VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO vliw
  CLASS BLOCK ;
  FOREIGN vliw ;
  ORIGIN 0.000 0.000 ;
  SIZE 2200.000 BY 850.000 ;
  PIN cache_PC[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.721000 ;
    PORT
      LAYER met2 ;
        RECT 26.770 846.000 27.050 850.000 ;
    END
  END cache_PC[0]
  PIN cache_PC[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 77.370 846.000 77.650 850.000 ;
    END
  END cache_PC[10]
  PIN cache_PC[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 82.430 846.000 82.710 850.000 ;
    END
  END cache_PC[11]
  PIN cache_PC[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 87.490 846.000 87.770 850.000 ;
    END
  END cache_PC[12]
  PIN cache_PC[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 92.550 846.000 92.830 850.000 ;
    END
  END cache_PC[13]
  PIN cache_PC[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 97.610 846.000 97.890 850.000 ;
    END
  END cache_PC[14]
  PIN cache_PC[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 102.670 846.000 102.950 850.000 ;
    END
  END cache_PC[15]
  PIN cache_PC[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 107.730 846.000 108.010 850.000 ;
    END
  END cache_PC[16]
  PIN cache_PC[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 112.790 846.000 113.070 850.000 ;
    END
  END cache_PC[17]
  PIN cache_PC[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 117.850 846.000 118.130 850.000 ;
    END
  END cache_PC[18]
  PIN cache_PC[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 122.910 846.000 123.190 850.000 ;
    END
  END cache_PC[19]
  PIN cache_PC[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 31.830 846.000 32.110 850.000 ;
    END
  END cache_PC[1]
  PIN cache_PC[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 127.970 846.000 128.250 850.000 ;
    END
  END cache_PC[20]
  PIN cache_PC[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 133.030 846.000 133.310 850.000 ;
    END
  END cache_PC[21]
  PIN cache_PC[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 138.090 846.000 138.370 850.000 ;
    END
  END cache_PC[22]
  PIN cache_PC[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 143.150 846.000 143.430 850.000 ;
    END
  END cache_PC[23]
  PIN cache_PC[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 148.210 846.000 148.490 850.000 ;
    END
  END cache_PC[24]
  PIN cache_PC[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 153.270 846.000 153.550 850.000 ;
    END
  END cache_PC[25]
  PIN cache_PC[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 158.330 846.000 158.610 850.000 ;
    END
  END cache_PC[26]
  PIN cache_PC[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 163.390 846.000 163.670 850.000 ;
    END
  END cache_PC[27]
  PIN cache_PC[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 36.890 846.000 37.170 850.000 ;
    END
  END cache_PC[2]
  PIN cache_PC[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.484000 ;
    PORT
      LAYER met2 ;
        RECT 41.950 846.000 42.230 850.000 ;
    END
  END cache_PC[3]
  PIN cache_PC[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 47.010 846.000 47.290 850.000 ;
    END
  END cache_PC[4]
  PIN cache_PC[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 52.070 846.000 52.350 850.000 ;
    END
  END cache_PC[5]
  PIN cache_PC[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 57.130 846.000 57.410 850.000 ;
    END
  END cache_PC[6]
  PIN cache_PC[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 62.190 846.000 62.470 850.000 ;
    END
  END cache_PC[7]
  PIN cache_PC[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 67.250 846.000 67.530 850.000 ;
    END
  END cache_PC[8]
  PIN cache_PC[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 72.310 846.000 72.590 850.000 ;
    END
  END cache_PC[9]
  PIN cache_entry[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 168.450 846.000 168.730 850.000 ;
    END
  END cache_entry[0]
  PIN cache_entry[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 674.450 846.000 674.730 850.000 ;
    END
  END cache_entry[100]
  PIN cache_entry[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 679.510 846.000 679.790 850.000 ;
    END
  END cache_entry[101]
  PIN cache_entry[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 684.570 846.000 684.850 850.000 ;
    END
  END cache_entry[102]
  PIN cache_entry[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 3.477600 ;
    PORT
      LAYER met2 ;
        RECT 689.630 846.000 689.910 850.000 ;
    END
  END cache_entry[103]
  PIN cache_entry[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 3.477600 ;
    PORT
      LAYER met2 ;
        RECT 694.690 846.000 694.970 850.000 ;
    END
  END cache_entry[104]
  PIN cache_entry[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 699.750 846.000 700.030 850.000 ;
    END
  END cache_entry[105]
  PIN cache_entry[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met2 ;
        RECT 704.810 846.000 705.090 850.000 ;
    END
  END cache_entry[106]
  PIN cache_entry[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 2.608200 ;
    PORT
      LAYER met2 ;
        RECT 709.870 846.000 710.150 850.000 ;
    END
  END cache_entry[107]
  PIN cache_entry[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 3.477600 ;
    PORT
      LAYER met2 ;
        RECT 714.930 846.000 715.210 850.000 ;
    END
  END cache_entry[108]
  PIN cache_entry[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 2.608200 ;
    PORT
      LAYER met2 ;
        RECT 719.990 846.000 720.270 850.000 ;
    END
  END cache_entry[109]
  PIN cache_entry[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 219.050 846.000 219.330 850.000 ;
    END
  END cache_entry[10]
  PIN cache_entry[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 12.171599 ;
    PORT
      LAYER met2 ;
        RECT 725.050 846.000 725.330 850.000 ;
    END
  END cache_entry[110]
  PIN cache_entry[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 730.110 846.000 730.390 850.000 ;
    END
  END cache_entry[111]
  PIN cache_entry[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 735.170 846.000 735.450 850.000 ;
    END
  END cache_entry[112]
  PIN cache_entry[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 740.230 846.000 740.510 850.000 ;
    END
  END cache_entry[113]
  PIN cache_entry[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 745.290 846.000 745.570 850.000 ;
    END
  END cache_entry[114]
  PIN cache_entry[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 750.350 846.000 750.630 850.000 ;
    END
  END cache_entry[115]
  PIN cache_entry[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 755.410 846.000 755.690 850.000 ;
    END
  END cache_entry[116]
  PIN cache_entry[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 760.470 846.000 760.750 850.000 ;
    END
  END cache_entry[117]
  PIN cache_entry[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 765.530 846.000 765.810 850.000 ;
    END
  END cache_entry[118]
  PIN cache_entry[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 770.590 846.000 770.870 850.000 ;
    END
  END cache_entry[119]
  PIN cache_entry[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 224.110 846.000 224.390 850.000 ;
    END
  END cache_entry[11]
  PIN cache_entry[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 775.650 846.000 775.930 850.000 ;
    END
  END cache_entry[120]
  PIN cache_entry[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 780.710 846.000 780.990 850.000 ;
    END
  END cache_entry[121]
  PIN cache_entry[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 785.770 846.000 786.050 850.000 ;
    END
  END cache_entry[122]
  PIN cache_entry[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 790.830 846.000 791.110 850.000 ;
    END
  END cache_entry[123]
  PIN cache_entry[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 795.890 846.000 796.170 850.000 ;
    END
  END cache_entry[124]
  PIN cache_entry[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 800.950 846.000 801.230 850.000 ;
    END
  END cache_entry[125]
  PIN cache_entry[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 806.010 846.000 806.290 850.000 ;
    END
  END cache_entry[126]
  PIN cache_entry[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 811.070 846.000 811.350 850.000 ;
    END
  END cache_entry[127]
  PIN cache_entry[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 229.170 846.000 229.450 850.000 ;
    END
  END cache_entry[12]
  PIN cache_entry[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 234.230 846.000 234.510 850.000 ;
    END
  END cache_entry[13]
  PIN cache_entry[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 239.290 846.000 239.570 850.000 ;
    END
  END cache_entry[14]
  PIN cache_entry[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 244.350 846.000 244.630 850.000 ;
    END
  END cache_entry[15]
  PIN cache_entry[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 249.410 846.000 249.690 850.000 ;
    END
  END cache_entry[16]
  PIN cache_entry[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 254.470 846.000 254.750 850.000 ;
    END
  END cache_entry[17]
  PIN cache_entry[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 259.530 846.000 259.810 850.000 ;
    END
  END cache_entry[18]
  PIN cache_entry[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 264.590 846.000 264.870 850.000 ;
    END
  END cache_entry[19]
  PIN cache_entry[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 173.510 846.000 173.790 850.000 ;
    END
  END cache_entry[1]
  PIN cache_entry[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 269.650 846.000 269.930 850.000 ;
    END
  END cache_entry[20]
  PIN cache_entry[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 274.710 846.000 274.990 850.000 ;
    END
  END cache_entry[21]
  PIN cache_entry[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 279.770 846.000 280.050 850.000 ;
    END
  END cache_entry[22]
  PIN cache_entry[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 284.830 846.000 285.110 850.000 ;
    END
  END cache_entry[23]
  PIN cache_entry[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 289.890 846.000 290.170 850.000 ;
    END
  END cache_entry[24]
  PIN cache_entry[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 294.950 846.000 295.230 850.000 ;
    END
  END cache_entry[25]
  PIN cache_entry[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 300.010 846.000 300.290 850.000 ;
    END
  END cache_entry[26]
  PIN cache_entry[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 305.070 846.000 305.350 850.000 ;
    END
  END cache_entry[27]
  PIN cache_entry[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 310.130 846.000 310.410 850.000 ;
    END
  END cache_entry[28]
  PIN cache_entry[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 315.190 846.000 315.470 850.000 ;
    END
  END cache_entry[29]
  PIN cache_entry[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 178.570 846.000 178.850 850.000 ;
    END
  END cache_entry[2]
  PIN cache_entry[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 320.250 846.000 320.530 850.000 ;
    END
  END cache_entry[30]
  PIN cache_entry[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 325.310 846.000 325.590 850.000 ;
    END
  END cache_entry[31]
  PIN cache_entry[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 330.370 846.000 330.650 850.000 ;
    END
  END cache_entry[32]
  PIN cache_entry[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 335.430 846.000 335.710 850.000 ;
    END
  END cache_entry[33]
  PIN cache_entry[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 340.490 846.000 340.770 850.000 ;
    END
  END cache_entry[34]
  PIN cache_entry[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 345.550 846.000 345.830 850.000 ;
    END
  END cache_entry[35]
  PIN cache_entry[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 350.610 846.000 350.890 850.000 ;
    END
  END cache_entry[36]
  PIN cache_entry[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 355.670 846.000 355.950 850.000 ;
    END
  END cache_entry[37]
  PIN cache_entry[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 360.730 846.000 361.010 850.000 ;
    END
  END cache_entry[38]
  PIN cache_entry[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 365.790 846.000 366.070 850.000 ;
    END
  END cache_entry[39]
  PIN cache_entry[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 183.630 846.000 183.910 850.000 ;
    END
  END cache_entry[3]
  PIN cache_entry[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 370.850 846.000 371.130 850.000 ;
    END
  END cache_entry[40]
  PIN cache_entry[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 375.910 846.000 376.190 850.000 ;
    END
  END cache_entry[41]
  PIN cache_entry[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 380.970 846.000 381.250 850.000 ;
    END
  END cache_entry[42]
  PIN cache_entry[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 386.030 846.000 386.310 850.000 ;
    END
  END cache_entry[43]
  PIN cache_entry[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 391.090 846.000 391.370 850.000 ;
    END
  END cache_entry[44]
  PIN cache_entry[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 396.150 846.000 396.430 850.000 ;
    END
  END cache_entry[45]
  PIN cache_entry[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 401.210 846.000 401.490 850.000 ;
    END
  END cache_entry[46]
  PIN cache_entry[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 406.270 846.000 406.550 850.000 ;
    END
  END cache_entry[47]
  PIN cache_entry[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 411.330 846.000 411.610 850.000 ;
    END
  END cache_entry[48]
  PIN cache_entry[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 416.390 846.000 416.670 850.000 ;
    END
  END cache_entry[49]
  PIN cache_entry[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 188.690 846.000 188.970 850.000 ;
    END
  END cache_entry[4]
  PIN cache_entry[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 421.450 846.000 421.730 850.000 ;
    END
  END cache_entry[50]
  PIN cache_entry[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 426.510 846.000 426.790 850.000 ;
    END
  END cache_entry[51]
  PIN cache_entry[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 431.570 846.000 431.850 850.000 ;
    END
  END cache_entry[52]
  PIN cache_entry[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 436.630 846.000 436.910 850.000 ;
    END
  END cache_entry[53]
  PIN cache_entry[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 441.690 846.000 441.970 850.000 ;
    END
  END cache_entry[54]
  PIN cache_entry[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 446.750 846.000 447.030 850.000 ;
    END
  END cache_entry[55]
  PIN cache_entry[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 451.810 846.000 452.090 850.000 ;
    END
  END cache_entry[56]
  PIN cache_entry[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 456.870 846.000 457.150 850.000 ;
    END
  END cache_entry[57]
  PIN cache_entry[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 461.930 846.000 462.210 850.000 ;
    END
  END cache_entry[58]
  PIN cache_entry[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 466.990 846.000 467.270 850.000 ;
    END
  END cache_entry[59]
  PIN cache_entry[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 193.750 846.000 194.030 850.000 ;
    END
  END cache_entry[5]
  PIN cache_entry[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 472.050 846.000 472.330 850.000 ;
    END
  END cache_entry[60]
  PIN cache_entry[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 477.110 846.000 477.390 850.000 ;
    END
  END cache_entry[61]
  PIN cache_entry[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 482.170 846.000 482.450 850.000 ;
    END
  END cache_entry[62]
  PIN cache_entry[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 487.230 846.000 487.510 850.000 ;
    END
  END cache_entry[63]
  PIN cache_entry[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 492.290 846.000 492.570 850.000 ;
    END
  END cache_entry[64]
  PIN cache_entry[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 497.350 846.000 497.630 850.000 ;
    END
  END cache_entry[65]
  PIN cache_entry[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 502.410 846.000 502.690 850.000 ;
    END
  END cache_entry[66]
  PIN cache_entry[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 507.470 846.000 507.750 850.000 ;
    END
  END cache_entry[67]
  PIN cache_entry[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 512.530 846.000 512.810 850.000 ;
    END
  END cache_entry[68]
  PIN cache_entry[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 517.590 846.000 517.870 850.000 ;
    END
  END cache_entry[69]
  PIN cache_entry[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 198.810 846.000 199.090 850.000 ;
    END
  END cache_entry[6]
  PIN cache_entry[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 522.650 846.000 522.930 850.000 ;
    END
  END cache_entry[70]
  PIN cache_entry[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 527.710 846.000 527.990 850.000 ;
    END
  END cache_entry[71]
  PIN cache_entry[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 532.770 846.000 533.050 850.000 ;
    END
  END cache_entry[72]
  PIN cache_entry[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 537.830 846.000 538.110 850.000 ;
    END
  END cache_entry[73]
  PIN cache_entry[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 542.890 846.000 543.170 850.000 ;
    END
  END cache_entry[74]
  PIN cache_entry[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 547.950 846.000 548.230 850.000 ;
    END
  END cache_entry[75]
  PIN cache_entry[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 553.010 846.000 553.290 850.000 ;
    END
  END cache_entry[76]
  PIN cache_entry[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 558.070 846.000 558.350 850.000 ;
    END
  END cache_entry[77]
  PIN cache_entry[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 563.130 846.000 563.410 850.000 ;
    END
  END cache_entry[78]
  PIN cache_entry[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 568.190 846.000 568.470 850.000 ;
    END
  END cache_entry[79]
  PIN cache_entry[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 203.870 846.000 204.150 850.000 ;
    END
  END cache_entry[7]
  PIN cache_entry[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 573.250 846.000 573.530 850.000 ;
    END
  END cache_entry[80]
  PIN cache_entry[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 578.310 846.000 578.590 850.000 ;
    END
  END cache_entry[81]
  PIN cache_entry[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 583.370 846.000 583.650 850.000 ;
    END
  END cache_entry[82]
  PIN cache_entry[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 588.430 846.000 588.710 850.000 ;
    END
  END cache_entry[83]
  PIN cache_entry[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 593.490 846.000 593.770 850.000 ;
    END
  END cache_entry[84]
  PIN cache_entry[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 598.550 846.000 598.830 850.000 ;
    END
  END cache_entry[85]
  PIN cache_entry[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 603.610 846.000 603.890 850.000 ;
    END
  END cache_entry[86]
  PIN cache_entry[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 608.670 846.000 608.950 850.000 ;
    END
  END cache_entry[87]
  PIN cache_entry[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 613.730 846.000 614.010 850.000 ;
    END
  END cache_entry[88]
  PIN cache_entry[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 618.790 846.000 619.070 850.000 ;
    END
  END cache_entry[89]
  PIN cache_entry[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 208.930 846.000 209.210 850.000 ;
    END
  END cache_entry[8]
  PIN cache_entry[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 623.850 846.000 624.130 850.000 ;
    END
  END cache_entry[90]
  PIN cache_entry[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 628.910 846.000 629.190 850.000 ;
    END
  END cache_entry[91]
  PIN cache_entry[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 633.970 846.000 634.250 850.000 ;
    END
  END cache_entry[92]
  PIN cache_entry[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 639.030 846.000 639.310 850.000 ;
    END
  END cache_entry[93]
  PIN cache_entry[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 644.090 846.000 644.370 850.000 ;
    END
  END cache_entry[94]
  PIN cache_entry[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 649.150 846.000 649.430 850.000 ;
    END
  END cache_entry[95]
  PIN cache_entry[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 2.608200 ;
    PORT
      LAYER met2 ;
        RECT 654.210 846.000 654.490 850.000 ;
    END
  END cache_entry[96]
  PIN cache_entry[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 3.477600 ;
    PORT
      LAYER met2 ;
        RECT 659.270 846.000 659.550 850.000 ;
    END
  END cache_entry[97]
  PIN cache_entry[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 2.608200 ;
    PORT
      LAYER met2 ;
        RECT 664.330 846.000 664.610 850.000 ;
    END
  END cache_entry[98]
  PIN cache_entry[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 669.390 846.000 669.670 850.000 ;
    END
  END cache_entry[99]
  PIN cache_entry[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 213.990 846.000 214.270 850.000 ;
    END
  END cache_entry[9]
  PIN cache_entry_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.484000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 102.040 2200.000 102.640 ;
    END
  END cache_entry_valid
  PIN cache_hit
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 93.880 2200.000 94.480 ;
    END
  END cache_hit
  PIN cache_invalidate
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 12.257999 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 96.600 2200.000 97.200 ;
    END
  END cache_invalidate
  PIN cache_new_entry[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END cache_new_entry[0]
  PIN cache_new_entry[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.737000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 915.950 0.000 916.230 4.000 ;
    END
  END cache_new_entry[100]
  PIN cache_new_entry[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.737000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 924.690 0.000 924.970 4.000 ;
    END
  END cache_new_entry[101]
  PIN cache_new_entry[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.737000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 933.430 0.000 933.710 4.000 ;
    END
  END cache_new_entry[102]
  PIN cache_new_entry[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.737000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 942.170 0.000 942.450 4.000 ;
    END
  END cache_new_entry[103]
  PIN cache_new_entry[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.737000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 950.910 0.000 951.190 4.000 ;
    END
  END cache_new_entry[104]
  PIN cache_new_entry[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.737000 ;
    ANTENNADIFFAREA 1.760400 ;
    PORT
      LAYER met2 ;
        RECT 959.650 0.000 959.930 4.000 ;
    END
  END cache_new_entry[105]
  PIN cache_new_entry[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.737000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 968.390 0.000 968.670 4.000 ;
    END
  END cache_new_entry[106]
  PIN cache_new_entry[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.737000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 977.130 0.000 977.410 4.000 ;
    END
  END cache_new_entry[107]
  PIN cache_new_entry[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.737000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 985.870 0.000 986.150 4.000 ;
    END
  END cache_new_entry[108]
  PIN cache_new_entry[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.737000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 994.610 0.000 994.890 4.000 ;
    END
  END cache_new_entry[109]
  PIN cache_new_entry[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 129.350 0.000 129.630 4.000 ;
    END
  END cache_new_entry[10]
  PIN cache_new_entry[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.747000 ;
    ANTENNADIFFAREA 2.195100 ;
    PORT
      LAYER met2 ;
        RECT 1003.350 0.000 1003.630 4.000 ;
    END
  END cache_new_entry[110]
  PIN cache_new_entry[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.994500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1012.090 0.000 1012.370 4.000 ;
    END
  END cache_new_entry[111]
  PIN cache_new_entry[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1020.830 0.000 1021.110 4.000 ;
    END
  END cache_new_entry[112]
  PIN cache_new_entry[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1029.570 0.000 1029.850 4.000 ;
    END
  END cache_new_entry[113]
  PIN cache_new_entry[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1038.310 0.000 1038.590 4.000 ;
    END
  END cache_new_entry[114]
  PIN cache_new_entry[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1047.050 0.000 1047.330 4.000 ;
    END
  END cache_new_entry[115]
  PIN cache_new_entry[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1055.790 0.000 1056.070 4.000 ;
    END
  END cache_new_entry[116]
  PIN cache_new_entry[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1064.530 0.000 1064.810 4.000 ;
    END
  END cache_new_entry[117]
  PIN cache_new_entry[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1073.270 0.000 1073.550 4.000 ;
    END
  END cache_new_entry[118]
  PIN cache_new_entry[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1082.010 0.000 1082.290 4.000 ;
    END
  END cache_new_entry[119]
  PIN cache_new_entry[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 138.090 0.000 138.370 4.000 ;
    END
  END cache_new_entry[11]
  PIN cache_new_entry[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1090.750 0.000 1091.030 4.000 ;
    END
  END cache_new_entry[120]
  PIN cache_new_entry[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1099.490 0.000 1099.770 4.000 ;
    END
  END cache_new_entry[121]
  PIN cache_new_entry[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1108.230 0.000 1108.510 4.000 ;
    END
  END cache_new_entry[122]
  PIN cache_new_entry[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1116.970 0.000 1117.250 4.000 ;
    END
  END cache_new_entry[123]
  PIN cache_new_entry[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1125.710 0.000 1125.990 4.000 ;
    END
  END cache_new_entry[124]
  PIN cache_new_entry[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1134.450 0.000 1134.730 4.000 ;
    END
  END cache_new_entry[125]
  PIN cache_new_entry[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1143.190 0.000 1143.470 4.000 ;
    END
  END cache_new_entry[126]
  PIN cache_new_entry[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1151.930 0.000 1152.210 4.000 ;
    END
  END cache_new_entry[127]
  PIN cache_new_entry[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 146.830 0.000 147.110 4.000 ;
    END
  END cache_new_entry[12]
  PIN cache_new_entry[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 155.570 0.000 155.850 4.000 ;
    END
  END cache_new_entry[13]
  PIN cache_new_entry[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 4.000 ;
    END
  END cache_new_entry[14]
  PIN cache_new_entry[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 173.050 0.000 173.330 4.000 ;
    END
  END cache_new_entry[15]
  PIN cache_new_entry[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 5.672700 ;
    PORT
      LAYER met2 ;
        RECT 181.790 0.000 182.070 4.000 ;
    END
  END cache_new_entry[16]
  PIN cache_new_entry[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 190.530 0.000 190.810 4.000 ;
    END
  END cache_new_entry[17]
  PIN cache_new_entry[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 199.270 0.000 199.550 4.000 ;
    END
  END cache_new_entry[18]
  PIN cache_new_entry[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 208.010 0.000 208.290 4.000 ;
    END
  END cache_new_entry[19]
  PIN cache_new_entry[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 50.690 0.000 50.970 4.000 ;
    END
  END cache_new_entry[1]
  PIN cache_new_entry[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 1.325700 ;
    PORT
      LAYER met2 ;
        RECT 216.750 0.000 217.030 4.000 ;
    END
  END cache_new_entry[20]
  PIN cache_new_entry[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 4.000 ;
    END
  END cache_new_entry[21]
  PIN cache_new_entry[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 234.230 0.000 234.510 4.000 ;
    END
  END cache_new_entry[22]
  PIN cache_new_entry[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 242.970 0.000 243.250 4.000 ;
    END
  END cache_new_entry[23]
  PIN cache_new_entry[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 251.710 0.000 251.990 4.000 ;
    END
  END cache_new_entry[24]
  PIN cache_new_entry[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 260.450 0.000 260.730 4.000 ;
    END
  END cache_new_entry[25]
  PIN cache_new_entry[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 269.190 0.000 269.470 4.000 ;
    END
  END cache_new_entry[26]
  PIN cache_new_entry[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 277.930 0.000 278.210 4.000 ;
    END
  END cache_new_entry[27]
  PIN cache_new_entry[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 286.670 0.000 286.950 4.000 ;
    END
  END cache_new_entry[28]
  PIN cache_new_entry[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 295.410 0.000 295.690 4.000 ;
    END
  END cache_new_entry[29]
  PIN cache_new_entry[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 59.430 0.000 59.710 4.000 ;
    END
  END cache_new_entry[2]
  PIN cache_new_entry[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 304.150 0.000 304.430 4.000 ;
    END
  END cache_new_entry[30]
  PIN cache_new_entry[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 312.890 0.000 313.170 4.000 ;
    END
  END cache_new_entry[31]
  PIN cache_new_entry[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 321.630 0.000 321.910 4.000 ;
    END
  END cache_new_entry[32]
  PIN cache_new_entry[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 1.325700 ;
    PORT
      LAYER met2 ;
        RECT 330.370 0.000 330.650 4.000 ;
    END
  END cache_new_entry[33]
  PIN cache_new_entry[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 1.325700 ;
    PORT
      LAYER met2 ;
        RECT 339.110 0.000 339.390 4.000 ;
    END
  END cache_new_entry[34]
  PIN cache_new_entry[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 347.850 0.000 348.130 4.000 ;
    END
  END cache_new_entry[35]
  PIN cache_new_entry[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 356.590 0.000 356.870 4.000 ;
    END
  END cache_new_entry[36]
  PIN cache_new_entry[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 365.330 0.000 365.610 4.000 ;
    END
  END cache_new_entry[37]
  PIN cache_new_entry[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 374.070 0.000 374.350 4.000 ;
    END
  END cache_new_entry[38]
  PIN cache_new_entry[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 382.810 0.000 383.090 4.000 ;
    END
  END cache_new_entry[39]
  PIN cache_new_entry[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 68.170 0.000 68.450 4.000 ;
    END
  END cache_new_entry[3]
  PIN cache_new_entry[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 391.550 0.000 391.830 4.000 ;
    END
  END cache_new_entry[40]
  PIN cache_new_entry[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 400.290 0.000 400.570 4.000 ;
    END
  END cache_new_entry[41]
  PIN cache_new_entry[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 409.030 0.000 409.310 4.000 ;
    END
  END cache_new_entry[42]
  PIN cache_new_entry[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 417.770 0.000 418.050 4.000 ;
    END
  END cache_new_entry[43]
  PIN cache_new_entry[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 426.510 0.000 426.790 4.000 ;
    END
  END cache_new_entry[44]
  PIN cache_new_entry[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 435.250 0.000 435.530 4.000 ;
    END
  END cache_new_entry[45]
  PIN cache_new_entry[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 1.325700 ;
    PORT
      LAYER met2 ;
        RECT 443.990 0.000 444.270 4.000 ;
    END
  END cache_new_entry[46]
  PIN cache_new_entry[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.489500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 452.730 0.000 453.010 4.000 ;
    END
  END cache_new_entry[47]
  PIN cache_new_entry[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 461.470 0.000 461.750 4.000 ;
    END
  END cache_new_entry[48]
  PIN cache_new_entry[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 470.210 0.000 470.490 4.000 ;
    END
  END cache_new_entry[49]
  PIN cache_new_entry[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 76.910 0.000 77.190 4.000 ;
    END
  END cache_new_entry[4]
  PIN cache_new_entry[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 478.950 0.000 479.230 4.000 ;
    END
  END cache_new_entry[50]
  PIN cache_new_entry[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 487.690 0.000 487.970 4.000 ;
    END
  END cache_new_entry[51]
  PIN cache_new_entry[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 496.430 0.000 496.710 4.000 ;
    END
  END cache_new_entry[52]
  PIN cache_new_entry[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 505.170 0.000 505.450 4.000 ;
    END
  END cache_new_entry[53]
  PIN cache_new_entry[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 513.910 0.000 514.190 4.000 ;
    END
  END cache_new_entry[54]
  PIN cache_new_entry[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 522.650 0.000 522.930 4.000 ;
    END
  END cache_new_entry[55]
  PIN cache_new_entry[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 531.390 0.000 531.670 4.000 ;
    END
  END cache_new_entry[56]
  PIN cache_new_entry[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 540.130 0.000 540.410 4.000 ;
    END
  END cache_new_entry[57]
  PIN cache_new_entry[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 548.870 0.000 549.150 4.000 ;
    END
  END cache_new_entry[58]
  PIN cache_new_entry[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 557.610 0.000 557.890 4.000 ;
    END
  END cache_new_entry[59]
  PIN cache_new_entry[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 85.650 0.000 85.930 4.000 ;
    END
  END cache_new_entry[5]
  PIN cache_new_entry[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 566.350 0.000 566.630 4.000 ;
    END
  END cache_new_entry[60]
  PIN cache_new_entry[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 1.325700 ;
    PORT
      LAYER met2 ;
        RECT 575.090 0.000 575.370 4.000 ;
    END
  END cache_new_entry[61]
  PIN cache_new_entry[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 1.760400 ;
    PORT
      LAYER met2 ;
        RECT 583.830 0.000 584.110 4.000 ;
    END
  END cache_new_entry[62]
  PIN cache_new_entry[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 592.570 0.000 592.850 4.000 ;
    END
  END cache_new_entry[63]
  PIN cache_new_entry[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 601.310 0.000 601.590 4.000 ;
    END
  END cache_new_entry[64]
  PIN cache_new_entry[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 610.050 0.000 610.330 4.000 ;
    END
  END cache_new_entry[65]
  PIN cache_new_entry[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 618.790 0.000 619.070 4.000 ;
    END
  END cache_new_entry[66]
  PIN cache_new_entry[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 1.325700 ;
    PORT
      LAYER met2 ;
        RECT 627.530 0.000 627.810 4.000 ;
    END
  END cache_new_entry[67]
  PIN cache_new_entry[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 636.270 0.000 636.550 4.000 ;
    END
  END cache_new_entry[68]
  PIN cache_new_entry[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 645.010 0.000 645.290 4.000 ;
    END
  END cache_new_entry[69]
  PIN cache_new_entry[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 94.390 0.000 94.670 4.000 ;
    END
  END cache_new_entry[6]
  PIN cache_new_entry[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 653.750 0.000 654.030 4.000 ;
    END
  END cache_new_entry[70]
  PIN cache_new_entry[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 12.236400 ;
    PORT
      LAYER met2 ;
        RECT 662.490 0.000 662.770 4.000 ;
    END
  END cache_new_entry[71]
  PIN cache_new_entry[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.499500 ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 671.230 0.000 671.510 4.000 ;
    END
  END cache_new_entry[72]
  PIN cache_new_entry[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 679.970 0.000 680.250 4.000 ;
    END
  END cache_new_entry[73]
  PIN cache_new_entry[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 4.368600 ;
    PORT
      LAYER met2 ;
        RECT 688.710 0.000 688.990 4.000 ;
    END
  END cache_new_entry[74]
  PIN cache_new_entry[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 697.450 0.000 697.730 4.000 ;
    END
  END cache_new_entry[75]
  PIN cache_new_entry[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 10.454400 ;
    PORT
      LAYER met2 ;
        RECT 706.190 0.000 706.470 4.000 ;
    END
  END cache_new_entry[76]
  PIN cache_new_entry[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 8.715600 ;
    PORT
      LAYER met2 ;
        RECT 714.930 0.000 715.210 4.000 ;
    END
  END cache_new_entry[77]
  PIN cache_new_entry[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 723.670 0.000 723.950 4.000 ;
    END
  END cache_new_entry[78]
  PIN cache_new_entry[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 732.410 0.000 732.690 4.000 ;
    END
  END cache_new_entry[79]
  PIN cache_new_entry[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END cache_new_entry[7]
  PIN cache_new_entry[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.499500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 741.150 0.000 741.430 4.000 ;
    END
  END cache_new_entry[80]
  PIN cache_new_entry[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 1.325700 ;
    PORT
      LAYER met2 ;
        RECT 749.890 0.000 750.170 4.000 ;
    END
  END cache_new_entry[81]
  PIN cache_new_entry[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 758.630 0.000 758.910 4.000 ;
    END
  END cache_new_entry[82]
  PIN cache_new_entry[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.499500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 767.370 0.000 767.650 4.000 ;
    END
  END cache_new_entry[83]
  PIN cache_new_entry[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.586500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 776.110 0.000 776.390 4.000 ;
    END
  END cache_new_entry[84]
  PIN cache_new_entry[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 784.850 0.000 785.130 4.000 ;
    END
  END cache_new_entry[85]
  PIN cache_new_entry[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 793.590 0.000 793.870 4.000 ;
    END
  END cache_new_entry[86]
  PIN cache_new_entry[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 802.330 0.000 802.610 4.000 ;
    END
  END cache_new_entry[87]
  PIN cache_new_entry[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 811.070 0.000 811.350 4.000 ;
    END
  END cache_new_entry[88]
  PIN cache_new_entry[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 819.810 0.000 820.090 4.000 ;
    END
  END cache_new_entry[89]
  PIN cache_new_entry[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 111.870 0.000 112.150 4.000 ;
    END
  END cache_new_entry[8]
  PIN cache_new_entry[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 828.550 0.000 828.830 4.000 ;
    END
  END cache_new_entry[90]
  PIN cache_new_entry[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 837.290 0.000 837.570 4.000 ;
    END
  END cache_new_entry[91]
  PIN cache_new_entry[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 846.030 0.000 846.310 4.000 ;
    END
  END cache_new_entry[92]
  PIN cache_new_entry[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 854.770 0.000 855.050 4.000 ;
    END
  END cache_new_entry[93]
  PIN cache_new_entry[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 863.510 0.000 863.790 4.000 ;
    END
  END cache_new_entry[94]
  PIN cache_new_entry[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 872.250 0.000 872.530 4.000 ;
    END
  END cache_new_entry[95]
  PIN cache_new_entry[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.737000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 880.990 0.000 881.270 4.000 ;
    END
  END cache_new_entry[96]
  PIN cache_new_entry[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.737000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 889.730 0.000 890.010 4.000 ;
    END
  END cache_new_entry[97]
  PIN cache_new_entry[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.737000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 898.470 0.000 898.750 4.000 ;
    END
  END cache_new_entry[98]
  PIN cache_new_entry[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.737000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 907.210 0.000 907.490 4.000 ;
    END
  END cache_new_entry[99]
  PIN cache_new_entry[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 120.610 0.000 120.890 4.000 ;
    END
  END cache_new_entry[9]
  PIN cache_rst
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 99.320 2200.000 99.920 ;
    END
  END cache_rst
  PIN curr_PC[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.275000 ;
    ANTENNADIFFAREA 1.760400 ;
    PORT
      LAYER met2 ;
        RECT 821.190 846.000 821.470 850.000 ;
    END
  END curr_PC[0]
  PIN curr_PC[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.967000 ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 871.790 846.000 872.070 850.000 ;
    END
  END curr_PC[10]
  PIN curr_PC[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.987000 ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 876.850 846.000 877.130 850.000 ;
    END
  END curr_PC[11]
  PIN curr_PC[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.588000 ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 881.910 846.000 882.190 850.000 ;
    END
  END curr_PC[12]
  PIN curr_PC[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.608000 ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 886.970 846.000 887.250 850.000 ;
    END
  END curr_PC[13]
  PIN curr_PC[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.845500 ;
    ANTENNADIFFAREA 4.411800 ;
    PORT
      LAYER met2 ;
        RECT 892.030 846.000 892.310 850.000 ;
    END
  END curr_PC[14]
  PIN curr_PC[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.865500 ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 897.090 846.000 897.370 850.000 ;
    END
  END curr_PC[15]
  PIN curr_PC[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.117500 ;
    ANTENNADIFFAREA 3.064500 ;
    PORT
      LAYER met2 ;
        RECT 902.150 846.000 902.430 850.000 ;
    END
  END curr_PC[16]
  PIN curr_PC[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.598000 ;
    ANTENNADIFFAREA 3.977100 ;
    PORT
      LAYER met2 ;
        RECT 907.210 846.000 907.490 850.000 ;
    END
  END curr_PC[17]
  PIN curr_PC[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.991500 ;
    ANTENNADIFFAREA 2.195100 ;
    PORT
      LAYER met2 ;
        RECT 912.270 846.000 912.550 850.000 ;
    END
  END curr_PC[18]
  PIN curr_PC[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.107500 ;
    ANTENNADIFFAREA 6.150600 ;
    PORT
      LAYER met2 ;
        RECT 917.330 846.000 917.610 850.000 ;
    END
  END curr_PC[19]
  PIN curr_PC[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.351500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 826.250 846.000 826.530 850.000 ;
    END
  END curr_PC[1]
  PIN curr_PC[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.093000 ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 922.390 846.000 922.670 850.000 ;
    END
  END curr_PC[20]
  PIN curr_PC[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.360500 ;
    ANTENNADIFFAREA 2.195100 ;
    PORT
      LAYER met2 ;
        RECT 927.450 846.000 927.730 850.000 ;
    END
  END curr_PC[21]
  PIN curr_PC[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.365000 ;
    ANTENNADIFFAREA 2.629800 ;
    PORT
      LAYER met2 ;
        RECT 932.510 846.000 932.790 850.000 ;
    END
  END curr_PC[22]
  PIN curr_PC[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.239000 ;
    ANTENNADIFFAREA 2.195100 ;
    PORT
      LAYER met2 ;
        RECT 937.570 846.000 937.850 850.000 ;
    END
  END curr_PC[23]
  PIN curr_PC[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.608000 ;
    ANTENNADIFFAREA 2.195100 ;
    PORT
      LAYER met2 ;
        RECT 942.630 846.000 942.910 850.000 ;
    END
  END curr_PC[24]
  PIN curr_PC[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.705000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 947.690 846.000 947.970 850.000 ;
    END
  END curr_PC[25]
  PIN curr_PC[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.363500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 952.750 846.000 953.030 850.000 ;
    END
  END curr_PC[26]
  PIN curr_PC[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.363500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 957.810 846.000 958.090 850.000 ;
    END
  END curr_PC[27]
  PIN curr_PC[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.654000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 831.310 846.000 831.590 850.000 ;
    END
  END curr_PC[2]
  PIN curr_PC[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 2.629800 ;
    PORT
      LAYER met2 ;
        RECT 836.370 846.000 836.650 850.000 ;
    END
  END curr_PC[3]
  PIN curr_PC[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.845500 ;
    ANTENNADIFFAREA 4.411800 ;
    PORT
      LAYER met2 ;
        RECT 841.430 846.000 841.710 850.000 ;
    END
  END curr_PC[4]
  PIN curr_PC[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.865500 ;
    ANTENNADIFFAREA 3.977100 ;
    PORT
      LAYER met2 ;
        RECT 846.490 846.000 846.770 850.000 ;
    END
  END curr_PC[5]
  PIN curr_PC[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.967000 ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 851.550 846.000 851.830 850.000 ;
    END
  END curr_PC[6]
  PIN curr_PC[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.987000 ;
    ANTENNADIFFAREA 3.977100 ;
    PORT
      LAYER met2 ;
        RECT 856.610 846.000 856.890 850.000 ;
    END
  END curr_PC[7]
  PIN curr_PC[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.845500 ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 861.670 846.000 861.950 850.000 ;
    END
  END curr_PC[8]
  PIN curr_PC[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.865500 ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 866.730 846.000 867.010 850.000 ;
    END
  END curr_PC[9]
  PIN custom_settings[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 2122.070 0.000 2122.350 4.000 ;
    END
  END custom_settings[0]
  PIN custom_settings[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 2130.810 0.000 2131.090 4.000 ;
    END
  END custom_settings[1]
  PIN custom_settings[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.719500 ;
    PORT
      LAYER met2 ;
        RECT 2139.550 0.000 2139.830 4.000 ;
    END
  END custom_settings[2]
  PIN custom_settings[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.719500 ;
    PORT
      LAYER met2 ;
        RECT 2148.290 0.000 2148.570 4.000 ;
    END
  END custom_settings[3]
  PIN custom_settings[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 2157.030 0.000 2157.310 4.000 ;
    END
  END custom_settings[4]
  PIN dest_idx0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 9.288000 ;
    PORT
      LAYER met2 ;
        RECT 1195.630 846.000 1195.910 850.000 ;
    END
  END dest_idx0[0]
  PIN dest_idx0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 6.318000 ;
    PORT
      LAYER met2 ;
        RECT 1200.690 846.000 1200.970 850.000 ;
    END
  END dest_idx0[1]
  PIN dest_idx0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 6.439500 ;
    PORT
      LAYER met2 ;
        RECT 1205.750 846.000 1206.030 850.000 ;
    END
  END dest_idx0[2]
  PIN dest_idx0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 9.531000 ;
    PORT
      LAYER met2 ;
        RECT 1210.810 846.000 1211.090 850.000 ;
    END
  END dest_idx0[3]
  PIN dest_idx0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 7.308000 ;
    PORT
      LAYER met2 ;
        RECT 1215.870 846.000 1216.150 850.000 ;
    END
  END dest_idx0[4]
  PIN dest_idx0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 6.934500 ;
    PORT
      LAYER met2 ;
        RECT 1220.930 846.000 1221.210 850.000 ;
    END
  END dest_idx0[5]
  PIN dest_idx1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 8.914500 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 229.880 2200.000 230.480 ;
    END
  END dest_idx1[0]
  PIN dest_idx1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.697000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 232.600 2200.000 233.200 ;
    END
  END dest_idx1[1]
  PIN dest_idx1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 6.070500 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 235.320 2200.000 235.920 ;
    END
  END dest_idx1[2]
  PIN dest_idx1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 8.419499 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 238.040 2200.000 238.640 ;
    END
  END dest_idx1[3]
  PIN dest_idx1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 7.186500 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 240.760 2200.000 241.360 ;
    END
  END dest_idx1[4]
  PIN dest_idx1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 6.813000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 243.480 2200.000 244.080 ;
    END
  END dest_idx1[5]
  PIN dest_idx2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.994500 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.440 4.000 225.040 ;
    END
  END dest_idx2[0]
  PIN dest_idx2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.744000 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.160 4.000 227.760 ;
    END
  END dest_idx2[1]
  PIN dest_idx2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.744000 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.880 4.000 230.480 ;
    END
  END dest_idx2[2]
  PIN dest_idx2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.994500 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 232.600 4.000 233.200 ;
    END
  END dest_idx2[3]
  PIN dest_idx2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.744000 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 0.000 235.320 4.000 235.920 ;
    END
  END dest_idx2[4]
  PIN dest_idx2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.744000 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.040 4.000 238.640 ;
    END
  END dest_idx2[5]
  PIN dest_mask0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.611000 ;
    PORT
      LAYER met2 ;
        RECT 1185.510 846.000 1185.790 850.000 ;
    END
  END dest_mask0[0]
  PIN dest_mask0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.363500 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met2 ;
        RECT 1190.570 846.000 1190.850 850.000 ;
    END
  END dest_mask0[1]
  PIN dest_mask1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.485000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 224.440 2200.000 225.040 ;
    END
  END dest_mask1[0]
  PIN dest_mask1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.980000 ;
    ANTENNADIFFAREA 3.477600 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 227.160 2200.000 227.760 ;
    END
  END dest_mask1[1]
  PIN dest_mask2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.000 4.000 219.600 ;
    END
  END dest_mask2[0]
  PIN dest_mask2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.737000 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.720 4.000 222.320 ;
    END
  END dest_mask2[1]
  PIN dest_pred0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.882000 ;
    ANTENNADIFFAREA 3.042900 ;
    PORT
      LAYER met2 ;
        RECT 1241.170 846.000 1241.450 850.000 ;
    END
  END dest_pred0[0]
  PIN dest_pred0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.882000 ;
    ANTENNADIFFAREA 3.042900 ;
    PORT
      LAYER met2 ;
        RECT 1246.230 846.000 1246.510 850.000 ;
    END
  END dest_pred0[1]
  PIN dest_pred0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.882000 ;
    ANTENNADIFFAREA 3.042900 ;
    PORT
      LAYER met2 ;
        RECT 1251.290 846.000 1251.570 850.000 ;
    END
  END dest_pred0[2]
  PIN dest_pred1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.625500 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 254.360 2200.000 254.960 ;
    END
  END dest_pred1[0]
  PIN dest_pred1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.877500 ;
    ANTENNADIFFAREA 2.608200 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 257.080 2200.000 257.680 ;
    END
  END dest_pred1[1]
  PIN dest_pred1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.877500 ;
    ANTENNADIFFAREA 2.608200 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 259.800 2200.000 260.400 ;
    END
  END dest_pred1[2]
  PIN dest_pred2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.630000 ;
    ANTENNADIFFAREA 2.173500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.920 4.000 249.520 ;
    END
  END dest_pred2[0]
  PIN dest_pred2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.368000 ;
    ANTENNADIFFAREA 2.608200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.640 4.000 252.240 ;
    END
  END dest_pred2[1]
  PIN dest_pred2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.494000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 254.360 4.000 254.960 ;
    END
  END dest_pred2[2]
  PIN dest_pred_val0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.882000 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met2 ;
        RECT 1256.350 846.000 1256.630 850.000 ;
    END
  END dest_pred_val0
  PIN dest_pred_val1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.999000 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 262.520 2200.000 263.120 ;
    END
  END dest_pred_val1
  PIN dest_pred_val2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.125000 ;
    ANTENNADIFFAREA 3.042900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 257.080 4.000 257.680 ;
    END
  END dest_pred_val2
  PIN dest_val0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1023.590 846.000 1023.870 850.000 ;
    END
  END dest_val0[0]
  PIN dest_val0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.475000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1074.190 846.000 1074.470 850.000 ;
    END
  END dest_val0[10]
  PIN dest_val0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.337000 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met2 ;
        RECT 1079.250 846.000 1079.530 850.000 ;
    END
  END dest_val0[11]
  PIN dest_val0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.485000 ;
    PORT
      LAYER met2 ;
        RECT 1084.310 846.000 1084.590 850.000 ;
    END
  END dest_val0[12]
  PIN dest_val0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.278000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1089.370 846.000 1089.650 850.000 ;
    END
  END dest_val0[13]
  PIN dest_val0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.416000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1094.430 846.000 1094.710 850.000 ;
    END
  END dest_val0[14]
  PIN dest_val0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.594500 ;
    PORT
      LAYER met2 ;
        RECT 1099.490 846.000 1099.770 850.000 ;
    END
  END dest_val0[15]
  PIN dest_val0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.230000 ;
    PORT
      LAYER met2 ;
        RECT 1104.550 846.000 1104.830 850.000 ;
    END
  END dest_val0[16]
  PIN dest_val0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.594500 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met2 ;
        RECT 1109.610 846.000 1109.890 850.000 ;
    END
  END dest_val0[17]
  PIN dest_val0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.224500 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met2 ;
        RECT 1114.670 846.000 1114.950 850.000 ;
    END
  END dest_val0[18]
  PIN dest_val0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.242000 ;
    PORT
      LAYER met2 ;
        RECT 1119.730 846.000 1120.010 850.000 ;
    END
  END dest_val0[19]
  PIN dest_val0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.134000 ;
    ANTENNADIFFAREA 2.608200 ;
    PORT
      LAYER met2 ;
        RECT 1028.650 846.000 1028.930 850.000 ;
    END
  END dest_val0[1]
  PIN dest_val0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.230000 ;
    PORT
      LAYER met2 ;
        RECT 1124.790 846.000 1125.070 850.000 ;
    END
  END dest_val0[20]
  PIN dest_val0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.846500 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met2 ;
        RECT 1129.850 846.000 1130.130 850.000 ;
    END
  END dest_val0[21]
  PIN dest_val0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.224500 ;
    PORT
      LAYER met2 ;
        RECT 1134.910 846.000 1135.190 850.000 ;
    END
  END dest_val0[22]
  PIN dest_val0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.416000 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met2 ;
        RECT 1139.970 846.000 1140.250 850.000 ;
    END
  END dest_val0[23]
  PIN dest_val0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.450500 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met2 ;
        RECT 1145.030 846.000 1145.310 850.000 ;
    END
  END dest_val0[24]
  PIN dest_val0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.450500 ;
    ANTENNADIFFAREA 3.912300 ;
    PORT
      LAYER met2 ;
        RECT 1150.090 846.000 1150.370 850.000 ;
    END
  END dest_val0[25]
  PIN dest_val0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807500 ;
    PORT
      LAYER met2 ;
        RECT 1155.150 846.000 1155.430 850.000 ;
    END
  END dest_val0[26]
  PIN dest_val0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.381500 ;
    ANTENNADIFFAREA 8.694000 ;
    PORT
      LAYER met2 ;
        RECT 1160.210 846.000 1160.490 850.000 ;
    END
  END dest_val0[27]
  PIN dest_val0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.644000 ;
    PORT
      LAYER met2 ;
        RECT 1165.270 846.000 1165.550 850.000 ;
    END
  END dest_val0[28]
  PIN dest_val0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 1170.330 846.000 1170.610 850.000 ;
    END
  END dest_val0[29]
  PIN dest_val0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.236500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1033.710 846.000 1033.990 850.000 ;
    END
  END dest_val0[2]
  PIN dest_val0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.124000 ;
    ANTENNADIFFAREA 2.173500 ;
    PORT
      LAYER met2 ;
        RECT 1175.390 846.000 1175.670 850.000 ;
    END
  END dest_val0[30]
  PIN dest_val0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.289000 ;
    PORT
      LAYER met2 ;
        RECT 1180.450 846.000 1180.730 850.000 ;
    END
  END dest_val0[31]
  PIN dest_val0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.794000 ;
    ANTENNADIFFAREA 5.651100 ;
    PORT
      LAYER met2 ;
        RECT 1038.770 846.000 1039.050 850.000 ;
    END
  END dest_val0[3]
  PIN dest_val0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1043.830 846.000 1044.110 850.000 ;
    END
  END dest_val0[4]
  PIN dest_val0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.007000 ;
    PORT
      LAYER met2 ;
        RECT 1048.890 846.000 1049.170 850.000 ;
    END
  END dest_val0[5]
  PIN dest_val0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.536500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1053.950 846.000 1054.230 850.000 ;
    END
  END dest_val0[6]
  PIN dest_val0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1059.010 846.000 1059.290 850.000 ;
    END
  END dest_val0[7]
  PIN dest_val0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.475000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1064.070 846.000 1064.350 850.000 ;
    END
  END dest_val0[8]
  PIN dest_val0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1069.130 846.000 1069.410 850.000 ;
    END
  END dest_val0[9]
  PIN dest_val1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 137.400 2200.000 138.000 ;
    END
  END dest_val1[0]
  PIN dest_val1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.980000 ;
    ANTENNADIFFAREA 2.173500 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 164.600 2200.000 165.200 ;
    END
  END dest_val1[10]
  PIN dest_val1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.406000 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 167.320 2200.000 167.920 ;
    END
  END dest_val1[11]
  PIN dest_val1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 170.040 2200.000 170.640 ;
    END
  END dest_val1[12]
  PIN dest_val1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.237500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 172.760 2200.000 173.360 ;
    END
  END dest_val1[13]
  PIN dest_val1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.168500 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 175.480 2200.000 176.080 ;
    END
  END dest_val1[14]
  PIN dest_val1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.485000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 178.200 2200.000 178.800 ;
    END
  END dest_val1[15]
  PIN dest_val1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.594500 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 180.920 2200.000 181.520 ;
    END
  END dest_val1[16]
  PIN dest_val1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.337000 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 183.640 2200.000 184.240 ;
    END
  END dest_val1[17]
  PIN dest_val1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.079500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 186.360 2200.000 186.960 ;
    END
  END dest_val1[18]
  PIN dest_val1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.485000 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 189.080 2200.000 189.680 ;
    END
  END dest_val1[19]
  PIN dest_val1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.203000 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 140.120 2200.000 140.720 ;
    END
  END dest_val1[1]
  PIN dest_val1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.732500 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 191.800 2200.000 192.400 ;
    END
  END dest_val1[20]
  PIN dest_val1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.227500 ;
    ANTENNADIFFAREA 3.042900 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 194.520 2200.000 195.120 ;
    END
  END dest_val1[21]
  PIN dest_val1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.079500 ;
    ANTENNADIFFAREA 2.608200 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 197.240 2200.000 197.840 ;
    END
  END dest_val1[22]
  PIN dest_val1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.842000 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 199.960 2200.000 200.560 ;
    END
  END dest_val1[23]
  PIN dest_val1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807500 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 202.680 2200.000 203.280 ;
    END
  END dest_val1[24]
  PIN dest_val1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.980000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 205.400 2200.000 206.000 ;
    END
  END dest_val1[25]
  PIN dest_val1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.842000 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 208.120 2200.000 208.720 ;
    END
  END dest_val1[26]
  PIN dest_val1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.450500 ;
    ANTENNADIFFAREA 6.085800 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 210.840 2200.000 211.440 ;
    END
  END dest_val1[27]
  PIN dest_val1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.203000 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 213.560 2200.000 214.160 ;
    END
  END dest_val1[28]
  PIN dest_val1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 216.280 2200.000 216.880 ;
    END
  END dest_val1[29]
  PIN dest_val1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.236500 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 142.840 2200.000 143.440 ;
    END
  END dest_val1[2]
  PIN dest_val1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.070000 ;
    ANTENNADIFFAREA 2.608200 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 219.000 2200.000 219.600 ;
    END
  END dest_val1[30]
  PIN dest_val1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 221.720 2200.000 222.320 ;
    END
  END dest_val1[31]
  PIN dest_val1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.863000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 145.560 2200.000 146.160 ;
    END
  END dest_val1[3]
  PIN dest_val1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 148.280 2200.000 148.880 ;
    END
  END dest_val1[4]
  PIN dest_val1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.828500 ;
    ANTENNADIFFAREA 3.042900 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 151.000 2200.000 151.600 ;
    END
  END dest_val1[5]
  PIN dest_val1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.915500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 153.720 2200.000 154.320 ;
    END
  END dest_val1[6]
  PIN dest_val1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 156.440 2200.000 157.040 ;
    END
  END dest_val1[7]
  PIN dest_val1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.311500 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 159.160 2200.000 159.760 ;
    END
  END dest_val1[8]
  PIN dest_val1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.167500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 161.880 2200.000 162.480 ;
    END
  END dest_val1[9]
  PIN dest_val2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.960 4.000 132.560 ;
    END
  END dest_val2[0]
  PIN dest_val2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.160 4.000 159.760 ;
    END
  END dest_val2[10]
  PIN dest_val2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.880 4.000 162.480 ;
    END
  END dest_val2[11]
  PIN dest_val2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 164.600 4.000 165.200 ;
    END
  END dest_val2[12]
  PIN dest_val2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 167.320 4.000 167.920 ;
    END
  END dest_val2[13]
  PIN dest_val2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END dest_val2[14]
  PIN dest_val2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.760 4.000 173.360 ;
    END
  END dest_val2[15]
  PIN dest_val2[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.347000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 175.480 4.000 176.080 ;
    END
  END dest_val2[16]
  PIN dest_val2[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.200 4.000 178.800 ;
    END
  END dest_val2[17]
  PIN dest_val2[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.621000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.920 4.000 181.520 ;
    END
  END dest_val2[18]
  PIN dest_val2[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.318000 ;
    ANTENNADIFFAREA 2.608200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END dest_val2[19]
  PIN dest_val2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    ANTENNADIFFAREA 3.042900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.680 4.000 135.280 ;
    END
  END dest_val2[1]
  PIN dest_val2[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 186.360 4.000 186.960 ;
    END
  END dest_val2[20]
  PIN dest_val2[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.080 4.000 189.680 ;
    END
  END dest_val2[21]
  PIN dest_val2[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.800 4.000 192.400 ;
    END
  END dest_val2[22]
  PIN dest_val2[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 194.520 4.000 195.120 ;
    END
  END dest_val2[23]
  PIN dest_val2[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.240 4.000 197.840 ;
    END
  END dest_val2[24]
  PIN dest_val2[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.485000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 199.960 4.000 200.560 ;
    END
  END dest_val2[25]
  PIN dest_val2[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.485000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 202.680 4.000 203.280 ;
    END
  END dest_val2[26]
  PIN dest_val2[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.485000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 205.400 4.000 206.000 ;
    END
  END dest_val2[27]
  PIN dest_val2[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 208.120 4.000 208.720 ;
    END
  END dest_val2[28]
  PIN dest_val2[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.840 4.000 211.440 ;
    END
  END dest_val2[29]
  PIN dest_val2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    ANTENNADIFFAREA 3.042900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.400 4.000 138.000 ;
    END
  END dest_val2[2]
  PIN dest_val2[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 213.560 4.000 214.160 ;
    END
  END dest_val2[30]
  PIN dest_val2[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.280 4.000 216.880 ;
    END
  END dest_val2[31]
  PIN dest_val2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.120 4.000 140.720 ;
    END
  END dest_val2[3]
  PIN dest_val2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    ANTENNADIFFAREA 2.608200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END dest_val2[4]
  PIN dest_val2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.560 4.000 146.160 ;
    END
  END dest_val2[5]
  PIN dest_val2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    ANTENNADIFFAREA 3.042900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.280 4.000 148.880 ;
    END
  END dest_val2[6]
  PIN dest_val2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    ANTENNADIFFAREA 3.042900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.000 4.000 151.600 ;
    END
  END dest_val2[7]
  PIN dest_val2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.720 4.000 154.320 ;
    END
  END dest_val2[8]
  PIN dest_val2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END dest_val2[9]
  PIN eu0_busy
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.485000 ;
    PORT
      LAYER met2 ;
        RECT 1625.730 846.000 1626.010 850.000 ;
    END
  END eu0_busy
  PIN eu0_instruction[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1630.790 846.000 1631.070 850.000 ;
    END
  END eu0_instruction[0]
  PIN eu0_instruction[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.499500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1681.390 846.000 1681.670 850.000 ;
    END
  END eu0_instruction[10]
  PIN eu0_instruction[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.499500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1686.450 846.000 1686.730 850.000 ;
    END
  END eu0_instruction[11]
  PIN eu0_instruction[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.499500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1691.510 846.000 1691.790 850.000 ;
    END
  END eu0_instruction[12]
  PIN eu0_instruction[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1696.570 846.000 1696.850 850.000 ;
    END
  END eu0_instruction[13]
  PIN eu0_instruction[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1701.630 846.000 1701.910 850.000 ;
    END
  END eu0_instruction[14]
  PIN eu0_instruction[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1706.690 846.000 1706.970 850.000 ;
    END
  END eu0_instruction[15]
  PIN eu0_instruction[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1711.750 846.000 1712.030 850.000 ;
    END
  END eu0_instruction[16]
  PIN eu0_instruction[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1716.810 846.000 1717.090 850.000 ;
    END
  END eu0_instruction[17]
  PIN eu0_instruction[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1721.870 846.000 1722.150 850.000 ;
    END
  END eu0_instruction[18]
  PIN eu0_instruction[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1726.930 846.000 1727.210 850.000 ;
    END
  END eu0_instruction[19]
  PIN eu0_instruction[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1635.850 846.000 1636.130 850.000 ;
    END
  END eu0_instruction[1]
  PIN eu0_instruction[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1731.990 846.000 1732.270 850.000 ;
    END
  END eu0_instruction[20]
  PIN eu0_instruction[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1737.050 846.000 1737.330 850.000 ;
    END
  END eu0_instruction[21]
  PIN eu0_instruction[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1742.110 846.000 1742.390 850.000 ;
    END
  END eu0_instruction[22]
  PIN eu0_instruction[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1747.170 846.000 1747.450 850.000 ;
    END
  END eu0_instruction[23]
  PIN eu0_instruction[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1752.230 846.000 1752.510 850.000 ;
    END
  END eu0_instruction[24]
  PIN eu0_instruction[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1757.290 846.000 1757.570 850.000 ;
    END
  END eu0_instruction[25]
  PIN eu0_instruction[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1762.350 846.000 1762.630 850.000 ;
    END
  END eu0_instruction[26]
  PIN eu0_instruction[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1767.410 846.000 1767.690 850.000 ;
    END
  END eu0_instruction[27]
  PIN eu0_instruction[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1772.470 846.000 1772.750 850.000 ;
    END
  END eu0_instruction[28]
  PIN eu0_instruction[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1777.530 846.000 1777.810 850.000 ;
    END
  END eu0_instruction[29]
  PIN eu0_instruction[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1640.910 846.000 1641.190 850.000 ;
    END
  END eu0_instruction[2]
  PIN eu0_instruction[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1782.590 846.000 1782.870 850.000 ;
    END
  END eu0_instruction[30]
  PIN eu0_instruction[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1787.650 846.000 1787.930 850.000 ;
    END
  END eu0_instruction[31]
  PIN eu0_instruction[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1792.710 846.000 1792.990 850.000 ;
    END
  END eu0_instruction[32]
  PIN eu0_instruction[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1797.770 846.000 1798.050 850.000 ;
    END
  END eu0_instruction[33]
  PIN eu0_instruction[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1802.830 846.000 1803.110 850.000 ;
    END
  END eu0_instruction[34]
  PIN eu0_instruction[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1807.890 846.000 1808.170 850.000 ;
    END
  END eu0_instruction[35]
  PIN eu0_instruction[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1812.950 846.000 1813.230 850.000 ;
    END
  END eu0_instruction[36]
  PIN eu0_instruction[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1818.010 846.000 1818.290 850.000 ;
    END
  END eu0_instruction[37]
  PIN eu0_instruction[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1823.070 846.000 1823.350 850.000 ;
    END
  END eu0_instruction[38]
  PIN eu0_instruction[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1828.130 846.000 1828.410 850.000 ;
    END
  END eu0_instruction[39]
  PIN eu0_instruction[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 12.236400 ;
    PORT
      LAYER met2 ;
        RECT 1645.970 846.000 1646.250 850.000 ;
    END
  END eu0_instruction[3]
  PIN eu0_instruction[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1833.190 846.000 1833.470 850.000 ;
    END
  END eu0_instruction[40]
  PIN eu0_instruction[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1838.250 846.000 1838.530 850.000 ;
    END
  END eu0_instruction[41]
  PIN eu0_instruction[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 12.236400 ;
    PORT
      LAYER met2 ;
        RECT 1651.030 846.000 1651.310 850.000 ;
    END
  END eu0_instruction[4]
  PIN eu0_instruction[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 12.236400 ;
    PORT
      LAYER met2 ;
        RECT 1656.090 846.000 1656.370 850.000 ;
    END
  END eu0_instruction[5]
  PIN eu0_instruction[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 7.020000 ;
    PORT
      LAYER met2 ;
        RECT 1661.150 846.000 1661.430 850.000 ;
    END
  END eu0_instruction[6]
  PIN eu0_instruction[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 10.454400 ;
    PORT
      LAYER met2 ;
        RECT 1666.210 846.000 1666.490 850.000 ;
    END
  END eu0_instruction[7]
  PIN eu0_instruction[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 10.454400 ;
    PORT
      LAYER met2 ;
        RECT 1671.270 846.000 1671.550 850.000 ;
    END
  END eu0_instruction[8]
  PIN eu0_instruction[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.499500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1676.330 846.000 1676.610 850.000 ;
    END
  END eu0_instruction[9]
  PIN eu1_busy
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.485000 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 461.080 2200.000 461.680 ;
    END
  END eu1_busy
  PIN eu1_instruction[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 463.800 2200.000 464.400 ;
    END
  END eu1_instruction[0]
  PIN eu1_instruction[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 491.000 2200.000 491.600 ;
    END
  END eu1_instruction[10]
  PIN eu1_instruction[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 493.720 2200.000 494.320 ;
    END
  END eu1_instruction[11]
  PIN eu1_instruction[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 496.440 2200.000 497.040 ;
    END
  END eu1_instruction[12]
  PIN eu1_instruction[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 499.160 2200.000 499.760 ;
    END
  END eu1_instruction[13]
  PIN eu1_instruction[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 501.880 2200.000 502.480 ;
    END
  END eu1_instruction[14]
  PIN eu1_instruction[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 504.600 2200.000 505.200 ;
    END
  END eu1_instruction[15]
  PIN eu1_instruction[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 507.320 2200.000 507.920 ;
    END
  END eu1_instruction[16]
  PIN eu1_instruction[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 510.040 2200.000 510.640 ;
    END
  END eu1_instruction[17]
  PIN eu1_instruction[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 512.760 2200.000 513.360 ;
    END
  END eu1_instruction[18]
  PIN eu1_instruction[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 515.480 2200.000 516.080 ;
    END
  END eu1_instruction[19]
  PIN eu1_instruction[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 466.520 2200.000 467.120 ;
    END
  END eu1_instruction[1]
  PIN eu1_instruction[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 518.200 2200.000 518.800 ;
    END
  END eu1_instruction[20]
  PIN eu1_instruction[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 520.920 2200.000 521.520 ;
    END
  END eu1_instruction[21]
  PIN eu1_instruction[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 523.640 2200.000 524.240 ;
    END
  END eu1_instruction[22]
  PIN eu1_instruction[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 526.360 2200.000 526.960 ;
    END
  END eu1_instruction[23]
  PIN eu1_instruction[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 529.080 2200.000 529.680 ;
    END
  END eu1_instruction[24]
  PIN eu1_instruction[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 531.800 2200.000 532.400 ;
    END
  END eu1_instruction[25]
  PIN eu1_instruction[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 534.520 2200.000 535.120 ;
    END
  END eu1_instruction[26]
  PIN eu1_instruction[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 537.240 2200.000 537.840 ;
    END
  END eu1_instruction[27]
  PIN eu1_instruction[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 539.960 2200.000 540.560 ;
    END
  END eu1_instruction[28]
  PIN eu1_instruction[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 542.680 2200.000 543.280 ;
    END
  END eu1_instruction[29]
  PIN eu1_instruction[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 469.240 2200.000 469.840 ;
    END
  END eu1_instruction[2]
  PIN eu1_instruction[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 545.400 2200.000 546.000 ;
    END
  END eu1_instruction[30]
  PIN eu1_instruction[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 548.120 2200.000 548.720 ;
    END
  END eu1_instruction[31]
  PIN eu1_instruction[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 550.840 2200.000 551.440 ;
    END
  END eu1_instruction[32]
  PIN eu1_instruction[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 553.560 2200.000 554.160 ;
    END
  END eu1_instruction[33]
  PIN eu1_instruction[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 556.280 2200.000 556.880 ;
    END
  END eu1_instruction[34]
  PIN eu1_instruction[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 559.000 2200.000 559.600 ;
    END
  END eu1_instruction[35]
  PIN eu1_instruction[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 561.720 2200.000 562.320 ;
    END
  END eu1_instruction[36]
  PIN eu1_instruction[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 564.440 2200.000 565.040 ;
    END
  END eu1_instruction[37]
  PIN eu1_instruction[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 567.160 2200.000 567.760 ;
    END
  END eu1_instruction[38]
  PIN eu1_instruction[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 569.880 2200.000 570.480 ;
    END
  END eu1_instruction[39]
  PIN eu1_instruction[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 471.960 2200.000 472.560 ;
    END
  END eu1_instruction[3]
  PIN eu1_instruction[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 572.600 2200.000 573.200 ;
    END
  END eu1_instruction[40]
  PIN eu1_instruction[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 575.320 2200.000 575.920 ;
    END
  END eu1_instruction[41]
  PIN eu1_instruction[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 474.680 2200.000 475.280 ;
    END
  END eu1_instruction[4]
  PIN eu1_instruction[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 477.400 2200.000 478.000 ;
    END
  END eu1_instruction[5]
  PIN eu1_instruction[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 480.120 2200.000 480.720 ;
    END
  END eu1_instruction[6]
  PIN eu1_instruction[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 482.840 2200.000 483.440 ;
    END
  END eu1_instruction[7]
  PIN eu1_instruction[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 485.560 2200.000 486.160 ;
    END
  END eu1_instruction[8]
  PIN eu1_instruction[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 488.280 2200.000 488.880 ;
    END
  END eu1_instruction[9]
  PIN eu2_busy
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.485000 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 0.000 455.640 4.000 456.240 ;
    END
  END eu2_busy
  PIN eu2_instruction[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 458.360 4.000 458.960 ;
    END
  END eu2_instruction[0]
  PIN eu2_instruction[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 485.560 4.000 486.160 ;
    END
  END eu2_instruction[10]
  PIN eu2_instruction[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 488.280 4.000 488.880 ;
    END
  END eu2_instruction[11]
  PIN eu2_instruction[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 491.000 4.000 491.600 ;
    END
  END eu2_instruction[12]
  PIN eu2_instruction[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 493.720 4.000 494.320 ;
    END
  END eu2_instruction[13]
  PIN eu2_instruction[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 496.440 4.000 497.040 ;
    END
  END eu2_instruction[14]
  PIN eu2_instruction[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 499.160 4.000 499.760 ;
    END
  END eu2_instruction[15]
  PIN eu2_instruction[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 501.880 4.000 502.480 ;
    END
  END eu2_instruction[16]
  PIN eu2_instruction[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 504.600 4.000 505.200 ;
    END
  END eu2_instruction[17]
  PIN eu2_instruction[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 507.320 4.000 507.920 ;
    END
  END eu2_instruction[18]
  PIN eu2_instruction[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 510.040 4.000 510.640 ;
    END
  END eu2_instruction[19]
  PIN eu2_instruction[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 461.080 4.000 461.680 ;
    END
  END eu2_instruction[1]
  PIN eu2_instruction[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 512.760 4.000 513.360 ;
    END
  END eu2_instruction[20]
  PIN eu2_instruction[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 515.480 4.000 516.080 ;
    END
  END eu2_instruction[21]
  PIN eu2_instruction[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 518.200 4.000 518.800 ;
    END
  END eu2_instruction[22]
  PIN eu2_instruction[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 520.920 4.000 521.520 ;
    END
  END eu2_instruction[23]
  PIN eu2_instruction[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 523.640 4.000 524.240 ;
    END
  END eu2_instruction[24]
  PIN eu2_instruction[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 526.360 4.000 526.960 ;
    END
  END eu2_instruction[25]
  PIN eu2_instruction[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 529.080 4.000 529.680 ;
    END
  END eu2_instruction[26]
  PIN eu2_instruction[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 531.800 4.000 532.400 ;
    END
  END eu2_instruction[27]
  PIN eu2_instruction[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 534.520 4.000 535.120 ;
    END
  END eu2_instruction[28]
  PIN eu2_instruction[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 537.240 4.000 537.840 ;
    END
  END eu2_instruction[29]
  PIN eu2_instruction[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 463.800 4.000 464.400 ;
    END
  END eu2_instruction[2]
  PIN eu2_instruction[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 539.960 4.000 540.560 ;
    END
  END eu2_instruction[30]
  PIN eu2_instruction[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 542.680 4.000 543.280 ;
    END
  END eu2_instruction[31]
  PIN eu2_instruction[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 545.400 4.000 546.000 ;
    END
  END eu2_instruction[32]
  PIN eu2_instruction[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 548.120 4.000 548.720 ;
    END
  END eu2_instruction[33]
  PIN eu2_instruction[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 550.840 4.000 551.440 ;
    END
  END eu2_instruction[34]
  PIN eu2_instruction[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 553.560 4.000 554.160 ;
    END
  END eu2_instruction[35]
  PIN eu2_instruction[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 556.280 4.000 556.880 ;
    END
  END eu2_instruction[36]
  PIN eu2_instruction[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 559.000 4.000 559.600 ;
    END
  END eu2_instruction[37]
  PIN eu2_instruction[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 561.720 4.000 562.320 ;
    END
  END eu2_instruction[38]
  PIN eu2_instruction[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 564.440 4.000 565.040 ;
    END
  END eu2_instruction[39]
  PIN eu2_instruction[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 466.520 4.000 467.120 ;
    END
  END eu2_instruction[3]
  PIN eu2_instruction[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 567.160 4.000 567.760 ;
    END
  END eu2_instruction[40]
  PIN eu2_instruction[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 569.880 4.000 570.480 ;
    END
  END eu2_instruction[41]
  PIN eu2_instruction[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 469.240 4.000 469.840 ;
    END
  END eu2_instruction[4]
  PIN eu2_instruction[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 471.960 4.000 472.560 ;
    END
  END eu2_instruction[5]
  PIN eu2_instruction[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 474.680 4.000 475.280 ;
    END
  END eu2_instruction[6]
  PIN eu2_instruction[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 477.400 4.000 478.000 ;
    END
  END eu2_instruction[7]
  PIN eu2_instruction[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 480.120 4.000 480.720 ;
    END
  END eu2_instruction[8]
  PIN eu2_instruction[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 482.840 4.000 483.440 ;
    END
  END eu2_instruction[9]
  PIN int_return0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met2 ;
        RECT 2172.210 846.000 2172.490 850.000 ;
    END
  END int_return0
  PIN int_return1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 9.998099 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 754.840 2200.000 755.440 ;
    END
  END int_return1
  PIN int_return2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 749.400 4.000 750.000 ;
    END
  END int_return2
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 1160.670 0.000 1160.950 4.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.232000 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met2 ;
        RECT 1248.070 0.000 1248.350 4.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.896000 ;
    PORT
      LAYER met2 ;
        RECT 1256.810 0.000 1257.090 4.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.863000 ;
    PORT
      LAYER met2 ;
        RECT 1265.550 0.000 1265.830 4.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.863000 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met2 ;
        RECT 1274.290 0.000 1274.570 4.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.863000 ;
    PORT
      LAYER met2 ;
        RECT 1283.030 0.000 1283.310 4.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.110500 ;
    ANTENNADIFFAREA 2.173500 ;
    PORT
      LAYER met2 ;
        RECT 1291.770 0.000 1292.050 4.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.110500 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met2 ;
        RECT 1300.510 0.000 1300.790 4.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.222000 ;
    PORT
      LAYER met2 ;
        RECT 1309.250 0.000 1309.530 4.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.459500 ;
    PORT
      LAYER met2 ;
        RECT 1317.990 0.000 1318.270 4.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1326.730 0.000 1327.010 4.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1169.410 0.000 1169.690 4.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1335.470 0.000 1335.750 4.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1344.210 0.000 1344.490 4.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1352.950 0.000 1353.230 4.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1361.690 0.000 1361.970 4.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1370.430 0.000 1370.710 4.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1379.170 0.000 1379.450 4.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.611000 ;
    PORT
      LAYER met2 ;
        RECT 1387.910 0.000 1388.190 4.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1396.650 0.000 1396.930 4.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1405.390 0.000 1405.670 4.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 1414.130 0.000 1414.410 4.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 1178.150 0.000 1178.430 4.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 2.173500 ;
    PORT
      LAYER met2 ;
        RECT 1422.870 0.000 1423.150 4.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.621000 ;
    PORT
      LAYER met2 ;
        RECT 1431.610 0.000 1431.890 4.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 1440.350 0.000 1440.630 4.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 1449.090 0.000 1449.370 4.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 2.608200 ;
    PORT
      LAYER met2 ;
        RECT 1457.830 0.000 1458.110 4.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met2 ;
        RECT 1466.570 0.000 1466.850 4.000 ;
    END
  END io_in[35]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.774500 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met2 ;
        RECT 1186.890 0.000 1187.170 4.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.727000 ;
    PORT
      LAYER met2 ;
        RECT 1195.630 0.000 1195.910 4.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.605500 ;
    PORT
      LAYER met2 ;
        RECT 1204.370 0.000 1204.650 4.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.863000 ;
    PORT
      LAYER met2 ;
        RECT 1213.110 0.000 1213.390 4.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.896000 ;
    PORT
      LAYER met2 ;
        RECT 1221.850 0.000 1222.130 4.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.232000 ;
    PORT
      LAYER met2 ;
        RECT 1230.590 0.000 1230.870 4.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.984500 ;
    PORT
      LAYER met2 ;
        RECT 1239.330 0.000 1239.610 4.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.484000 ;
    PORT
      LAYER met2 ;
        RECT 1475.310 0.000 1475.590 4.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1562.710 0.000 1562.990 4.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1571.450 0.000 1571.730 4.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1580.190 0.000 1580.470 4.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1588.930 0.000 1589.210 4.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1597.670 0.000 1597.950 4.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1606.410 0.000 1606.690 4.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1615.150 0.000 1615.430 4.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1623.890 0.000 1624.170 4.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 12.870000 ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1632.630 0.000 1632.910 4.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1641.370 0.000 1641.650 4.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1484.050 0.000 1484.330 4.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1650.110 0.000 1650.390 4.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1658.850 0.000 1659.130 4.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1667.590 0.000 1667.870 4.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1676.330 0.000 1676.610 4.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1685.070 0.000 1685.350 4.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1693.810 0.000 1694.090 4.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1702.550 0.000 1702.830 4.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1711.290 0.000 1711.570 4.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1720.030 0.000 1720.310 4.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1728.770 0.000 1729.050 4.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.484000 ;
    PORT
      LAYER met2 ;
        RECT 1492.790 0.000 1493.070 4.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 13.127399 ;
    PORT
      LAYER met2 ;
        RECT 1737.510 0.000 1737.790 4.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1746.250 0.000 1746.530 4.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1754.990 0.000 1755.270 4.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1763.730 0.000 1764.010 4.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1772.470 0.000 1772.750 4.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1781.210 0.000 1781.490 4.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1501.530 0.000 1501.810 4.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1510.270 0.000 1510.550 4.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1519.010 0.000 1519.290 4.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1527.750 0.000 1528.030 4.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1536.490 0.000 1536.770 4.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1545.230 0.000 1545.510 4.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1553.970 0.000 1554.250 4.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1789.950 0.000 1790.230 4.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1877.350 0.000 1877.630 4.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1886.090 0.000 1886.370 4.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1894.830 0.000 1895.110 4.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1903.570 0.000 1903.850 4.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1912.310 0.000 1912.590 4.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1921.050 0.000 1921.330 4.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1929.790 0.000 1930.070 4.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1938.530 0.000 1938.810 4.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1947.270 0.000 1947.550 4.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1956.010 0.000 1956.290 4.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1798.690 0.000 1798.970 4.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1964.750 0.000 1965.030 4.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1973.490 0.000 1973.770 4.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1982.230 0.000 1982.510 4.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1990.970 0.000 1991.250 4.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1999.710 0.000 1999.990 4.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 2008.450 0.000 2008.730 4.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2017.190 0.000 2017.470 4.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 9.585000 ;
    PORT
      LAYER met2 ;
        RECT 2025.930 0.000 2026.210 4.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 10.454400 ;
    PORT
      LAYER met2 ;
        RECT 2034.670 0.000 2034.950 4.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2043.410 0.000 2043.690 4.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1807.430 0.000 1807.710 4.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 2052.150 0.000 2052.430 4.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 2.195100 ;
    PORT
      LAYER met2 ;
        RECT 2060.890 0.000 2061.170 4.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 2069.630 0.000 2069.910 4.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 10.454400 ;
    PORT
      LAYER met2 ;
        RECT 2078.370 0.000 2078.650 4.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 3.499200 ;
    PORT
      LAYER met2 ;
        RECT 2087.110 0.000 2087.390 4.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 10.454400 ;
    PORT
      LAYER met2 ;
        RECT 2095.850 0.000 2096.130 4.000 ;
    END
  END io_out[35]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1816.170 0.000 1816.450 4.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1824.910 0.000 1825.190 4.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1833.650 0.000 1833.930 4.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1842.390 0.000 1842.670 4.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1851.130 0.000 1851.410 4.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1859.870 0.000 1860.150 4.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1868.610 0.000 1868.890 4.000 ;
    END
  END io_out[9]
  PIN is_load0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.237500 ;
    PORT
      LAYER met2 ;
        RECT 1423.330 846.000 1423.610 850.000 ;
    END
  END is_load0
  PIN is_load1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 352.280 2200.000 352.880 ;
    END
  END is_load1
  PIN is_load2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    ANTENNADIFFAREA 3.042900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.840 4.000 347.440 ;
    END
  END is_load2
  PIN is_store0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1428.390 846.000 1428.670 850.000 ;
    END
  END is_store0
  PIN is_store1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 355.000 2200.000 355.600 ;
    END
  END is_store1
  PIN is_store2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 3.477600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 349.560 4.000 350.160 ;
    END
  END is_store2
  PIN loadstore_address0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 3.912300 ;
    PORT
      LAYER met2 ;
        RECT 1261.410 846.000 1261.690 850.000 ;
    END
  END loadstore_address0[0]
  PIN loadstore_address0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 3.477600 ;
    PORT
      LAYER met2 ;
        RECT 1312.010 846.000 1312.290 850.000 ;
    END
  END loadstore_address0[10]
  PIN loadstore_address0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 1317.070 846.000 1317.350 850.000 ;
    END
  END loadstore_address0[11]
  PIN loadstore_address0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met2 ;
        RECT 1322.130 846.000 1322.410 850.000 ;
    END
  END loadstore_address0[12]
  PIN loadstore_address0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 3.912300 ;
    PORT
      LAYER met2 ;
        RECT 1327.190 846.000 1327.470 850.000 ;
    END
  END loadstore_address0[13]
  PIN loadstore_address0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 2.608200 ;
    PORT
      LAYER met2 ;
        RECT 1332.250 846.000 1332.530 850.000 ;
    END
  END loadstore_address0[14]
  PIN loadstore_address0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 3.477600 ;
    PORT
      LAYER met2 ;
        RECT 1337.310 846.000 1337.590 850.000 ;
    END
  END loadstore_address0[15]
  PIN loadstore_address0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 3.912300 ;
    PORT
      LAYER met2 ;
        RECT 1342.370 846.000 1342.650 850.000 ;
    END
  END loadstore_address0[16]
  PIN loadstore_address0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 3.042900 ;
    PORT
      LAYER met2 ;
        RECT 1347.430 846.000 1347.710 850.000 ;
    END
  END loadstore_address0[17]
  PIN loadstore_address0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 2.608200 ;
    PORT
      LAYER met2 ;
        RECT 1352.490 846.000 1352.770 850.000 ;
    END
  END loadstore_address0[18]
  PIN loadstore_address0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 2.173500 ;
    PORT
      LAYER met2 ;
        RECT 1357.550 846.000 1357.830 850.000 ;
    END
  END loadstore_address0[19]
  PIN loadstore_address0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.347000 ;
    PORT
      LAYER met2 ;
        RECT 1266.470 846.000 1266.750 850.000 ;
    END
  END loadstore_address0[1]
  PIN loadstore_address0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 3.042900 ;
    PORT
      LAYER met2 ;
        RECT 1362.610 846.000 1362.890 850.000 ;
    END
  END loadstore_address0[20]
  PIN loadstore_address0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 3.042900 ;
    PORT
      LAYER met2 ;
        RECT 1367.670 846.000 1367.950 850.000 ;
    END
  END loadstore_address0[21]
  PIN loadstore_address0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 3.042900 ;
    PORT
      LAYER met2 ;
        RECT 1372.730 846.000 1373.010 850.000 ;
    END
  END loadstore_address0[22]
  PIN loadstore_address0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met2 ;
        RECT 1377.790 846.000 1378.070 850.000 ;
    END
  END loadstore_address0[23]
  PIN loadstore_address0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met2 ;
        RECT 1382.850 846.000 1383.130 850.000 ;
    END
  END loadstore_address0[24]
  PIN loadstore_address0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met2 ;
        RECT 1387.910 846.000 1388.190 850.000 ;
    END
  END loadstore_address0[25]
  PIN loadstore_address0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1392.970 846.000 1393.250 850.000 ;
    END
  END loadstore_address0[26]
  PIN loadstore_address0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met2 ;
        RECT 1398.030 846.000 1398.310 850.000 ;
    END
  END loadstore_address0[27]
  PIN loadstore_address0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met2 ;
        RECT 1403.090 846.000 1403.370 850.000 ;
    END
  END loadstore_address0[28]
  PIN loadstore_address0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1408.150 846.000 1408.430 850.000 ;
    END
  END loadstore_address0[29]
  PIN loadstore_address0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1271.530 846.000 1271.810 850.000 ;
    END
  END loadstore_address0[2]
  PIN loadstore_address0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met2 ;
        RECT 1413.210 846.000 1413.490 850.000 ;
    END
  END loadstore_address0[30]
  PIN loadstore_address0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 2.173500 ;
    PORT
      LAYER met2 ;
        RECT 1418.270 846.000 1418.550 850.000 ;
    END
  END loadstore_address0[31]
  PIN loadstore_address0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 3.042900 ;
    PORT
      LAYER met2 ;
        RECT 1276.590 846.000 1276.870 850.000 ;
    END
  END loadstore_address0[3]
  PIN loadstore_address0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 5.651100 ;
    PORT
      LAYER met2 ;
        RECT 1281.650 846.000 1281.930 850.000 ;
    END
  END loadstore_address0[4]
  PIN loadstore_address0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 2.608200 ;
    PORT
      LAYER met2 ;
        RECT 1286.710 846.000 1286.990 850.000 ;
    END
  END loadstore_address0[5]
  PIN loadstore_address0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 3.042900 ;
    PORT
      LAYER met2 ;
        RECT 1291.770 846.000 1292.050 850.000 ;
    END
  END loadstore_address0[6]
  PIN loadstore_address0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 3.477600 ;
    PORT
      LAYER met2 ;
        RECT 1296.830 846.000 1297.110 850.000 ;
    END
  END loadstore_address0[7]
  PIN loadstore_address0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 3.912300 ;
    PORT
      LAYER met2 ;
        RECT 1301.890 846.000 1302.170 850.000 ;
    END
  END loadstore_address0[8]
  PIN loadstore_address0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 3.042900 ;
    PORT
      LAYER met2 ;
        RECT 1306.950 846.000 1307.230 850.000 ;
    END
  END loadstore_address0[9]
  PIN loadstore_address1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 265.240 2200.000 265.840 ;
    END
  END loadstore_address1[0]
  PIN loadstore_address1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 5.216400 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 292.440 2200.000 293.040 ;
    END
  END loadstore_address1[10]
  PIN loadstore_address1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 9.998099 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 295.160 2200.000 295.760 ;
    END
  END loadstore_address1[11]
  PIN loadstore_address1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 9.998099 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 297.880 2200.000 298.480 ;
    END
  END loadstore_address1[12]
  PIN loadstore_address1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 300.600 2200.000 301.200 ;
    END
  END loadstore_address1[13]
  PIN loadstore_address1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 303.320 2200.000 303.920 ;
    END
  END loadstore_address1[14]
  PIN loadstore_address1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 9.998099 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 306.040 2200.000 306.640 ;
    END
  END loadstore_address1[15]
  PIN loadstore_address1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 16.518600 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 308.760 2200.000 309.360 ;
    END
  END loadstore_address1[16]
  PIN loadstore_address1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 311.480 2200.000 312.080 ;
    END
  END loadstore_address1[17]
  PIN loadstore_address1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 9.998099 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 314.200 2200.000 314.800 ;
    END
  END loadstore_address1[18]
  PIN loadstore_address1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 316.920 2200.000 317.520 ;
    END
  END loadstore_address1[19]
  PIN loadstore_address1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 267.960 2200.000 268.560 ;
    END
  END loadstore_address1[1]
  PIN loadstore_address1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 319.640 2200.000 320.240 ;
    END
  END loadstore_address1[20]
  PIN loadstore_address1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 9.998099 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 322.360 2200.000 322.960 ;
    END
  END loadstore_address1[21]
  PIN loadstore_address1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 9.998099 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 325.080 2200.000 325.680 ;
    END
  END loadstore_address1[22]
  PIN loadstore_address1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 327.800 2200.000 328.400 ;
    END
  END loadstore_address1[23]
  PIN loadstore_address1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 12.606299 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 330.520 2200.000 331.120 ;
    END
  END loadstore_address1[24]
  PIN loadstore_address1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 9.998099 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 333.240 2200.000 333.840 ;
    END
  END loadstore_address1[25]
  PIN loadstore_address1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 335.960 2200.000 336.560 ;
    END
  END loadstore_address1[26]
  PIN loadstore_address1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 12.606299 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 338.680 2200.000 339.280 ;
    END
  END loadstore_address1[27]
  PIN loadstore_address1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 341.400 2200.000 342.000 ;
    END
  END loadstore_address1[28]
  PIN loadstore_address1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 9.998099 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 344.120 2200.000 344.720 ;
    END
  END loadstore_address1[29]
  PIN loadstore_address1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 270.680 2200.000 271.280 ;
    END
  END loadstore_address1[2]
  PIN loadstore_address1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 346.840 2200.000 347.440 ;
    END
  END loadstore_address1[30]
  PIN loadstore_address1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 9.998099 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 349.560 2200.000 350.160 ;
    END
  END loadstore_address1[31]
  PIN loadstore_address1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 273.400 2200.000 274.000 ;
    END
  END loadstore_address1[3]
  PIN loadstore_address1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 13.475699 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 276.120 2200.000 276.720 ;
    END
  END loadstore_address1[4]
  PIN loadstore_address1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 278.840 2200.000 279.440 ;
    END
  END loadstore_address1[5]
  PIN loadstore_address1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 281.560 2200.000 282.160 ;
    END
  END loadstore_address1[6]
  PIN loadstore_address1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 20.430899 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 284.280 2200.000 284.880 ;
    END
  END loadstore_address1[7]
  PIN loadstore_address1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 17.822701 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 287.000 2200.000 287.600 ;
    END
  END loadstore_address1[8]
  PIN loadstore_address1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 9.998099 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 289.720 2200.000 290.320 ;
    END
  END loadstore_address1[9]
  PIN loadstore_address2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 18.692099 ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.800 4.000 260.400 ;
    END
  END loadstore_address2[0]
  PIN loadstore_address2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 15.214499 ;
    PORT
      LAYER met3 ;
        RECT 0.000 287.000 4.000 287.600 ;
    END
  END loadstore_address2[10]
  PIN loadstore_address2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 15.214499 ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.720 4.000 290.320 ;
    END
  END loadstore_address2[11]
  PIN loadstore_address2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 9.563399 ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.440 4.000 293.040 ;
    END
  END loadstore_address2[12]
  PIN loadstore_address2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 9.998099 ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.160 4.000 295.760 ;
    END
  END loadstore_address2[13]
  PIN loadstore_address2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 12.606299 ;
    PORT
      LAYER met3 ;
        RECT 0.000 297.880 4.000 298.480 ;
    END
  END loadstore_address2[14]
  PIN loadstore_address2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 15.214499 ;
    PORT
      LAYER met3 ;
        RECT 0.000 300.600 4.000 301.200 ;
    END
  END loadstore_address2[15]
  PIN loadstore_address2[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 15.214499 ;
    PORT
      LAYER met3 ;
        RECT 0.000 303.320 4.000 303.920 ;
    END
  END loadstore_address2[16]
  PIN loadstore_address2[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 14.345099 ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.040 4.000 306.640 ;
    END
  END loadstore_address2[17]
  PIN loadstore_address2[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 32.167801 ;
    PORT
      LAYER met3 ;
        RECT 0.000 308.760 4.000 309.360 ;
    END
  END loadstore_address2[18]
  PIN loadstore_address2[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 13.475699 ;
    PORT
      LAYER met3 ;
        RECT 0.000 311.480 4.000 312.080 ;
    END
  END loadstore_address2[19]
  PIN loadstore_address2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 9.998099 ;
    PORT
      LAYER met3 ;
        RECT 0.000 262.520 4.000 263.120 ;
    END
  END loadstore_address2[1]
  PIN loadstore_address2[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 6.955200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 314.200 4.000 314.800 ;
    END
  END loadstore_address2[20]
  PIN loadstore_address2[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 26.081999 ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.920 4.000 317.520 ;
    END
  END loadstore_address2[21]
  PIN loadstore_address2[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 26.951399 ;
    PORT
      LAYER met3 ;
        RECT 0.000 319.640 4.000 320.240 ;
    END
  END loadstore_address2[22]
  PIN loadstore_address2[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 12.606299 ;
    PORT
      LAYER met3 ;
        RECT 0.000 322.360 4.000 322.960 ;
    END
  END loadstore_address2[23]
  PIN loadstore_address2[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 8.259300 ;
    PORT
      LAYER met3 ;
        RECT 0.000 325.080 4.000 325.680 ;
    END
  END loadstore_address2[24]
  PIN loadstore_address2[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 9.998099 ;
    PORT
      LAYER met3 ;
        RECT 0.000 327.800 4.000 328.400 ;
    END
  END loadstore_address2[25]
  PIN loadstore_address2[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 15.214499 ;
    PORT
      LAYER met3 ;
        RECT 0.000 330.520 4.000 331.120 ;
    END
  END loadstore_address2[26]
  PIN loadstore_address2[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 15.214499 ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.240 4.000 333.840 ;
    END
  END loadstore_address2[27]
  PIN loadstore_address2[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 335.960 4.000 336.560 ;
    END
  END loadstore_address2[28]
  PIN loadstore_address2[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 13.475699 ;
    PORT
      LAYER met3 ;
        RECT 0.000 338.680 4.000 339.280 ;
    END
  END loadstore_address2[29]
  PIN loadstore_address2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 15.214499 ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.240 4.000 265.840 ;
    END
  END loadstore_address2[2]
  PIN loadstore_address2[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 10.867499 ;
    PORT
      LAYER met3 ;
        RECT 0.000 341.400 4.000 342.000 ;
    END
  END loadstore_address2[30]
  PIN loadstore_address2[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 15.214499 ;
    PORT
      LAYER met3 ;
        RECT 0.000 344.120 4.000 344.720 ;
    END
  END loadstore_address2[31]
  PIN loadstore_address2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 15.214499 ;
    PORT
      LAYER met3 ;
        RECT 0.000 267.960 4.000 268.560 ;
    END
  END loadstore_address2[3]
  PIN loadstore_address2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 24.777899 ;
    PORT
      LAYER met3 ;
        RECT 0.000 270.680 4.000 271.280 ;
    END
  END loadstore_address2[4]
  PIN loadstore_address2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 10.867499 ;
    PORT
      LAYER met3 ;
        RECT 0.000 273.400 4.000 274.000 ;
    END
  END loadstore_address2[5]
  PIN loadstore_address2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 15.214499 ;
    PORT
      LAYER met3 ;
        RECT 0.000 276.120 4.000 276.720 ;
    END
  END loadstore_address2[6]
  PIN loadstore_address2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 18.257399 ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.840 4.000 279.440 ;
    END
  END loadstore_address2[7]
  PIN loadstore_address2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 16.953300 ;
    PORT
      LAYER met3 ;
        RECT 0.000 281.560 4.000 282.160 ;
    END
  END loadstore_address2[8]
  PIN loadstore_address2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 284.280 4.000 284.880 ;
    END
  END loadstore_address2[9]
  PIN loadstore_dest0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met2 ;
        RECT 1448.630 846.000 1448.910 850.000 ;
    END
  END loadstore_dest0[0]
  PIN loadstore_dest0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met2 ;
        RECT 1453.690 846.000 1453.970 850.000 ;
    END
  END loadstore_dest0[1]
  PIN loadstore_dest0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met2 ;
        RECT 1458.750 846.000 1459.030 850.000 ;
    END
  END loadstore_dest0[2]
  PIN loadstore_dest0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met2 ;
        RECT 1463.810 846.000 1464.090 850.000 ;
    END
  END loadstore_dest0[3]
  PIN loadstore_dest0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met2 ;
        RECT 1468.870 846.000 1469.150 850.000 ;
    END
  END loadstore_dest0[4]
  PIN loadstore_dest0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met2 ;
        RECT 1473.930 846.000 1474.210 850.000 ;
    END
  END loadstore_dest0[5]
  PIN loadstore_dest1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.237500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 365.880 2200.000 366.480 ;
    END
  END loadstore_dest1[0]
  PIN loadstore_dest1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.237500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 368.600 2200.000 369.200 ;
    END
  END loadstore_dest1[1]
  PIN loadstore_dest1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.485000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 371.320 2200.000 371.920 ;
    END
  END loadstore_dest1[2]
  PIN loadstore_dest1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.485000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 374.040 2200.000 374.640 ;
    END
  END loadstore_dest1[3]
  PIN loadstore_dest1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.485000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 376.760 2200.000 377.360 ;
    END
  END loadstore_dest1[4]
  PIN loadstore_dest1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.485000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 379.480 2200.000 380.080 ;
    END
  END loadstore_dest1[5]
  PIN loadstore_dest2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.237500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 360.440 4.000 361.040 ;
    END
  END loadstore_dest2[0]
  PIN loadstore_dest2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.237500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.160 4.000 363.760 ;
    END
  END loadstore_dest2[1]
  PIN loadstore_dest2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.485000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 365.880 4.000 366.480 ;
    END
  END loadstore_dest2[2]
  PIN loadstore_dest2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.485000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 368.600 4.000 369.200 ;
    END
  END loadstore_dest2[3]
  PIN loadstore_dest2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.485000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 371.320 4.000 371.920 ;
    END
  END loadstore_dest2[4]
  PIN loadstore_dest2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.485000 ;
    ANTENNADIFFAREA 2.173500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.040 4.000 374.640 ;
    END
  END loadstore_dest2[5]
  PIN loadstore_size0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met2 ;
        RECT 1438.510 846.000 1438.790 850.000 ;
    END
  END loadstore_size0[0]
  PIN loadstore_size0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 2.173500 ;
    PORT
      LAYER met2 ;
        RECT 1443.570 846.000 1443.850 850.000 ;
    END
  END loadstore_size0[1]
  PIN loadstore_size1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 360.440 2200.000 361.040 ;
    END
  END loadstore_size1[0]
  PIN loadstore_size1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 363.160 2200.000 363.760 ;
    END
  END loadstore_size1[1]
  PIN loadstore_size2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 15.214499 ;
    PORT
      LAYER met3 ;
        RECT 0.000 355.000 4.000 355.600 ;
    END
  END loadstore_size2[0]
  PIN loadstore_size2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 12.606299 ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.720 4.000 358.320 ;
    END
  END loadstore_size2[1]
  PIN new_PC0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1484.050 846.000 1484.330 850.000 ;
    END
  END new_PC0[0]
  PIN new_PC0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met2 ;
        RECT 1534.650 846.000 1534.930 850.000 ;
    END
  END new_PC0[10]
  PIN new_PC0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1539.710 846.000 1539.990 850.000 ;
    END
  END new_PC0[11]
  PIN new_PC0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1544.770 846.000 1545.050 850.000 ;
    END
  END new_PC0[12]
  PIN new_PC0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1549.830 846.000 1550.110 850.000 ;
    END
  END new_PC0[13]
  PIN new_PC0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1554.890 846.000 1555.170 850.000 ;
    END
  END new_PC0[14]
  PIN new_PC0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1559.950 846.000 1560.230 850.000 ;
    END
  END new_PC0[15]
  PIN new_PC0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 3.477600 ;
    PORT
      LAYER met2 ;
        RECT 1565.010 846.000 1565.290 850.000 ;
    END
  END new_PC0[16]
  PIN new_PC0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 5.216400 ;
    PORT
      LAYER met2 ;
        RECT 1570.070 846.000 1570.350 850.000 ;
    END
  END new_PC0[17]
  PIN new_PC0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1575.130 846.000 1575.410 850.000 ;
    END
  END new_PC0[18]
  PIN new_PC0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1580.190 846.000 1580.470 850.000 ;
    END
  END new_PC0[19]
  PIN new_PC0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 2.173500 ;
    PORT
      LAYER met2 ;
        RECT 1489.110 846.000 1489.390 850.000 ;
    END
  END new_PC0[1]
  PIN new_PC0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met2 ;
        RECT 1585.250 846.000 1585.530 850.000 ;
    END
  END new_PC0[20]
  PIN new_PC0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.347000 ;
    PORT
      LAYER met2 ;
        RECT 1590.310 846.000 1590.590 850.000 ;
    END
  END new_PC0[21]
  PIN new_PC0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1595.370 846.000 1595.650 850.000 ;
    END
  END new_PC0[22]
  PIN new_PC0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 2.173500 ;
    PORT
      LAYER met2 ;
        RECT 1600.430 846.000 1600.710 850.000 ;
    END
  END new_PC0[23]
  PIN new_PC0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1605.490 846.000 1605.770 850.000 ;
    END
  END new_PC0[24]
  PIN new_PC0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1610.550 846.000 1610.830 850.000 ;
    END
  END new_PC0[25]
  PIN new_PC0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1615.610 846.000 1615.890 850.000 ;
    END
  END new_PC0[26]
  PIN new_PC0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 3.912300 ;
    PORT
      LAYER met2 ;
        RECT 1620.670 846.000 1620.950 850.000 ;
    END
  END new_PC0[27]
  PIN new_PC0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 2.173500 ;
    PORT
      LAYER met2 ;
        RECT 1494.170 846.000 1494.450 850.000 ;
    END
  END new_PC0[2]
  PIN new_PC0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 7.389900 ;
    PORT
      LAYER met2 ;
        RECT 1499.230 846.000 1499.510 850.000 ;
    END
  END new_PC0[3]
  PIN new_PC0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 1504.290 846.000 1504.570 850.000 ;
    END
  END new_PC0[4]
  PIN new_PC0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1509.350 846.000 1509.630 850.000 ;
    END
  END new_PC0[5]
  PIN new_PC0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 5.216400 ;
    PORT
      LAYER met2 ;
        RECT 1514.410 846.000 1514.690 850.000 ;
    END
  END new_PC0[6]
  PIN new_PC0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1519.470 846.000 1519.750 850.000 ;
    END
  END new_PC0[7]
  PIN new_PC0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 1524.530 846.000 1524.810 850.000 ;
    END
  END new_PC0[8]
  PIN new_PC0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met2 ;
        RECT 1529.590 846.000 1529.870 850.000 ;
    END
  END new_PC0[9]
  PIN new_PC1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 384.920 2200.000 385.520 ;
    END
  END new_PC1[0]
  PIN new_PC1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 9.998099 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 412.120 2200.000 412.720 ;
    END
  END new_PC1[10]
  PIN new_PC1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 414.840 2200.000 415.440 ;
    END
  END new_PC1[11]
  PIN new_PC1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 417.560 2200.000 418.160 ;
    END
  END new_PC1[12]
  PIN new_PC1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 420.280 2200.000 420.880 ;
    END
  END new_PC1[13]
  PIN new_PC1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 423.000 2200.000 423.600 ;
    END
  END new_PC1[14]
  PIN new_PC1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 425.720 2200.000 426.320 ;
    END
  END new_PC1[15]
  PIN new_PC1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 428.440 2200.000 429.040 ;
    END
  END new_PC1[16]
  PIN new_PC1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 15.214499 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 431.160 2200.000 431.760 ;
    END
  END new_PC1[17]
  PIN new_PC1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 433.880 2200.000 434.480 ;
    END
  END new_PC1[18]
  PIN new_PC1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 436.600 2200.000 437.200 ;
    END
  END new_PC1[19]
  PIN new_PC1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 15.214499 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 387.640 2200.000 388.240 ;
    END
  END new_PC1[1]
  PIN new_PC1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 439.320 2200.000 439.920 ;
    END
  END new_PC1[20]
  PIN new_PC1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 442.040 2200.000 442.640 ;
    END
  END new_PC1[21]
  PIN new_PC1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 444.760 2200.000 445.360 ;
    END
  END new_PC1[22]
  PIN new_PC1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 447.480 2200.000 448.080 ;
    END
  END new_PC1[23]
  PIN new_PC1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 450.200 2200.000 450.800 ;
    END
  END new_PC1[24]
  PIN new_PC1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 452.920 2200.000 453.520 ;
    END
  END new_PC1[25]
  PIN new_PC1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 455.640 2200.000 456.240 ;
    END
  END new_PC1[26]
  PIN new_PC1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 458.360 2200.000 458.960 ;
    END
  END new_PC1[27]
  PIN new_PC1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 390.360 2200.000 390.960 ;
    END
  END new_PC1[2]
  PIN new_PC1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 15.214499 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 393.080 2200.000 393.680 ;
    END
  END new_PC1[3]
  PIN new_PC1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 9.998099 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 395.800 2200.000 396.400 ;
    END
  END new_PC1[4]
  PIN new_PC1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 398.520 2200.000 399.120 ;
    END
  END new_PC1[5]
  PIN new_PC1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 401.240 2200.000 401.840 ;
    END
  END new_PC1[6]
  PIN new_PC1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.304000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 403.960 2200.000 404.560 ;
    END
  END new_PC1[7]
  PIN new_PC1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 30.863699 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 406.680 2200.000 407.280 ;
    END
  END new_PC1[8]
  PIN new_PC1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 9.998099 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 409.400 2200.000 410.000 ;
    END
  END new_PC1[9]
  PIN new_PC2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 379.480 4.000 380.080 ;
    END
  END new_PC2[0]
  PIN new_PC2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 406.680 4.000 407.280 ;
    END
  END new_PC2[10]
  PIN new_PC2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 409.400 4.000 410.000 ;
    END
  END new_PC2[11]
  PIN new_PC2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 412.120 4.000 412.720 ;
    END
  END new_PC2[12]
  PIN new_PC2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 414.840 4.000 415.440 ;
    END
  END new_PC2[13]
  PIN new_PC2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 417.560 4.000 418.160 ;
    END
  END new_PC2[14]
  PIN new_PC2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 420.280 4.000 420.880 ;
    END
  END new_PC2[15]
  PIN new_PC2[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 423.000 4.000 423.600 ;
    END
  END new_PC2[16]
  PIN new_PC2[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 425.720 4.000 426.320 ;
    END
  END new_PC2[17]
  PIN new_PC2[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 428.440 4.000 429.040 ;
    END
  END new_PC2[18]
  PIN new_PC2[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 431.160 4.000 431.760 ;
    END
  END new_PC2[19]
  PIN new_PC2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 382.200 4.000 382.800 ;
    END
  END new_PC2[1]
  PIN new_PC2[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 433.880 4.000 434.480 ;
    END
  END new_PC2[20]
  PIN new_PC2[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 436.600 4.000 437.200 ;
    END
  END new_PC2[21]
  PIN new_PC2[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 439.320 4.000 439.920 ;
    END
  END new_PC2[22]
  PIN new_PC2[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 442.040 4.000 442.640 ;
    END
  END new_PC2[23]
  PIN new_PC2[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 444.760 4.000 445.360 ;
    END
  END new_PC2[24]
  PIN new_PC2[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 447.480 4.000 448.080 ;
    END
  END new_PC2[25]
  PIN new_PC2[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 450.200 4.000 450.800 ;
    END
  END new_PC2[26]
  PIN new_PC2[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 452.920 4.000 453.520 ;
    END
  END new_PC2[27]
  PIN new_PC2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.920 4.000 385.520 ;
    END
  END new_PC2[2]
  PIN new_PC2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 387.640 4.000 388.240 ;
    END
  END new_PC2[3]
  PIN new_PC2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 390.360 4.000 390.960 ;
    END
  END new_PC2[4]
  PIN new_PC2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 393.080 4.000 393.680 ;
    END
  END new_PC2[5]
  PIN new_PC2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 395.800 4.000 396.400 ;
    END
  END new_PC2[6]
  PIN new_PC2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 398.520 4.000 399.120 ;
    END
  END new_PC2[7]
  PIN new_PC2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 401.240 4.000 401.840 ;
    END
  END new_PC2[8]
  PIN new_PC2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 403.960 4.000 404.560 ;
    END
  END new_PC2[9]
  PIN pred_idx0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.630000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1225.990 846.000 1226.270 850.000 ;
    END
  END pred_idx0[0]
  PIN pred_idx0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.630000 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met2 ;
        RECT 1231.050 846.000 1231.330 850.000 ;
    END
  END pred_idx0[1]
  PIN pred_idx0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1236.110 846.000 1236.390 850.000 ;
    END
  END pred_idx0[2]
  PIN pred_idx1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.630000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 246.200 2200.000 246.800 ;
    END
  END pred_idx1[0]
  PIN pred_idx1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.630000 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 248.920 2200.000 249.520 ;
    END
  END pred_idx1[1]
  PIN pred_idx1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    ANTENNADIFFAREA 10.432799 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 251.640 2200.000 252.240 ;
    END
  END pred_idx1[2]
  PIN pred_idx2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.630000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.760 4.000 241.360 ;
    END
  END pred_idx2[0]
  PIN pred_idx2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.630000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 243.480 4.000 244.080 ;
    END
  END pred_idx2[1]
  PIN pred_idx2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 246.200 4.000 246.800 ;
    END
  END pred_idx2[2]
  PIN pred_val0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.962500 ;
    PORT
      LAYER met2 ;
        RECT 2167.150 846.000 2167.430 850.000 ;
    END
  END pred_val0
  PIN pred_val1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.962500 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 752.120 2200.000 752.720 ;
    END
  END pred_val1
  PIN pred_val2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.962500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 746.680 4.000 747.280 ;
    END
  END pred_val2
  PIN reg1_idx0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 962.870 846.000 963.150 850.000 ;
    END
  END reg1_idx0[0]
  PIN reg1_idx0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.980000 ;
    PORT
      LAYER met2 ;
        RECT 967.930 846.000 968.210 850.000 ;
    END
  END reg1_idx0[1]
  PIN reg1_idx0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.773500 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met2 ;
        RECT 972.990 846.000 973.270 850.000 ;
    END
  END reg1_idx0[2]
  PIN reg1_idx0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.980000 ;
    PORT
      LAYER met2 ;
        RECT 978.050 846.000 978.330 850.000 ;
    END
  END reg1_idx0[3]
  PIN reg1_idx0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.722500 ;
    PORT
      LAYER met2 ;
        RECT 983.110 846.000 983.390 850.000 ;
    END
  END reg1_idx0[4]
  PIN reg1_idx0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.475000 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met2 ;
        RECT 988.170 846.000 988.450 850.000 ;
    END
  END reg1_idx0[5]
  PIN reg1_idx1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 6.049500 ;
    ANTENNADIFFAREA 2.173500 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 104.760 2200.000 105.360 ;
    END
  END reg1_idx1[0]
  PIN reg1_idx1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.633500 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 107.480 2200.000 108.080 ;
    END
  END reg1_idx1[1]
  PIN reg1_idx1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 110.200 2200.000 110.800 ;
    END
  END reg1_idx1[2]
  PIN reg1_idx1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 112.920 2200.000 113.520 ;
    END
  END reg1_idx1[3]
  PIN reg1_idx1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.722500 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 115.640 2200.000 116.240 ;
    END
  END reg1_idx1[4]
  PIN reg1_idx1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.712500 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 118.360 2200.000 118.960 ;
    END
  END reg1_idx1[5]
  PIN reg1_idx2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.832000 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 0.000 99.320 4.000 99.920 ;
    END
  END reg1_idx2[0]
  PIN reg1_idx2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.970000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END reg1_idx2[1]
  PIN reg1_idx2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.398000 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.760 4.000 105.360 ;
    END
  END reg1_idx2[2]
  PIN reg1_idx2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.079500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 107.480 4.000 108.080 ;
    END
  END reg1_idx2[3]
  PIN reg1_idx2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.793000 ;
    ANTENNADIFFAREA 5.651100 ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.200 4.000 110.800 ;
    END
  END reg1_idx2[4]
  PIN reg1_idx2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.980000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.920 4.000 113.520 ;
    END
  END reg1_idx2[5]
  PIN reg1_val0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1843.310 846.000 1843.590 850.000 ;
    END
  END reg1_val0[0]
  PIN reg1_val0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1893.910 846.000 1894.190 850.000 ;
    END
  END reg1_val0[10]
  PIN reg1_val0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1898.970 846.000 1899.250 850.000 ;
    END
  END reg1_val0[11]
  PIN reg1_val0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1904.030 846.000 1904.310 850.000 ;
    END
  END reg1_val0[12]
  PIN reg1_val0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1909.090 846.000 1909.370 850.000 ;
    END
  END reg1_val0[13]
  PIN reg1_val0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1914.150 846.000 1914.430 850.000 ;
    END
  END reg1_val0[14]
  PIN reg1_val0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1919.210 846.000 1919.490 850.000 ;
    END
  END reg1_val0[15]
  PIN reg1_val0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1924.270 846.000 1924.550 850.000 ;
    END
  END reg1_val0[16]
  PIN reg1_val0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1929.330 846.000 1929.610 850.000 ;
    END
  END reg1_val0[17]
  PIN reg1_val0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1934.390 846.000 1934.670 850.000 ;
    END
  END reg1_val0[18]
  PIN reg1_val0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1939.450 846.000 1939.730 850.000 ;
    END
  END reg1_val0[19]
  PIN reg1_val0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1848.370 846.000 1848.650 850.000 ;
    END
  END reg1_val0[1]
  PIN reg1_val0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1944.510 846.000 1944.790 850.000 ;
    END
  END reg1_val0[20]
  PIN reg1_val0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1949.570 846.000 1949.850 850.000 ;
    END
  END reg1_val0[21]
  PIN reg1_val0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1954.630 846.000 1954.910 850.000 ;
    END
  END reg1_val0[22]
  PIN reg1_val0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1959.690 846.000 1959.970 850.000 ;
    END
  END reg1_val0[23]
  PIN reg1_val0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1964.750 846.000 1965.030 850.000 ;
    END
  END reg1_val0[24]
  PIN reg1_val0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1969.810 846.000 1970.090 850.000 ;
    END
  END reg1_val0[25]
  PIN reg1_val0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1974.870 846.000 1975.150 850.000 ;
    END
  END reg1_val0[26]
  PIN reg1_val0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1979.930 846.000 1980.210 850.000 ;
    END
  END reg1_val0[27]
  PIN reg1_val0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1984.990 846.000 1985.270 850.000 ;
    END
  END reg1_val0[28]
  PIN reg1_val0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1990.050 846.000 1990.330 850.000 ;
    END
  END reg1_val0[29]
  PIN reg1_val0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1853.430 846.000 1853.710 850.000 ;
    END
  END reg1_val0[2]
  PIN reg1_val0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1995.110 846.000 1995.390 850.000 ;
    END
  END reg1_val0[30]
  PIN reg1_val0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 2000.170 846.000 2000.450 850.000 ;
    END
  END reg1_val0[31]
  PIN reg1_val0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1858.490 846.000 1858.770 850.000 ;
    END
  END reg1_val0[3]
  PIN reg1_val0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1863.550 846.000 1863.830 850.000 ;
    END
  END reg1_val0[4]
  PIN reg1_val0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1868.610 846.000 1868.890 850.000 ;
    END
  END reg1_val0[5]
  PIN reg1_val0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1873.670 846.000 1873.950 850.000 ;
    END
  END reg1_val0[6]
  PIN reg1_val0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1878.730 846.000 1879.010 850.000 ;
    END
  END reg1_val0[7]
  PIN reg1_val0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1883.790 846.000 1884.070 850.000 ;
    END
  END reg1_val0[8]
  PIN reg1_val0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1888.850 846.000 1889.130 850.000 ;
    END
  END reg1_val0[9]
  PIN reg1_val1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 578.040 2200.000 578.640 ;
    END
  END reg1_val1[0]
  PIN reg1_val1[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 605.240 2200.000 605.840 ;
    END
  END reg1_val1[10]
  PIN reg1_val1[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 607.960 2200.000 608.560 ;
    END
  END reg1_val1[11]
  PIN reg1_val1[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 610.680 2200.000 611.280 ;
    END
  END reg1_val1[12]
  PIN reg1_val1[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 613.400 2200.000 614.000 ;
    END
  END reg1_val1[13]
  PIN reg1_val1[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 616.120 2200.000 616.720 ;
    END
  END reg1_val1[14]
  PIN reg1_val1[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 618.840 2200.000 619.440 ;
    END
  END reg1_val1[15]
  PIN reg1_val1[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 621.560 2200.000 622.160 ;
    END
  END reg1_val1[16]
  PIN reg1_val1[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 624.280 2200.000 624.880 ;
    END
  END reg1_val1[17]
  PIN reg1_val1[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 627.000 2200.000 627.600 ;
    END
  END reg1_val1[18]
  PIN reg1_val1[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 629.720 2200.000 630.320 ;
    END
  END reg1_val1[19]
  PIN reg1_val1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 580.760 2200.000 581.360 ;
    END
  END reg1_val1[1]
  PIN reg1_val1[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 632.440 2200.000 633.040 ;
    END
  END reg1_val1[20]
  PIN reg1_val1[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 635.160 2200.000 635.760 ;
    END
  END reg1_val1[21]
  PIN reg1_val1[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 637.880 2200.000 638.480 ;
    END
  END reg1_val1[22]
  PIN reg1_val1[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 640.600 2200.000 641.200 ;
    END
  END reg1_val1[23]
  PIN reg1_val1[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 643.320 2200.000 643.920 ;
    END
  END reg1_val1[24]
  PIN reg1_val1[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 646.040 2200.000 646.640 ;
    END
  END reg1_val1[25]
  PIN reg1_val1[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 648.760 2200.000 649.360 ;
    END
  END reg1_val1[26]
  PIN reg1_val1[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 651.480 2200.000 652.080 ;
    END
  END reg1_val1[27]
  PIN reg1_val1[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 654.200 2200.000 654.800 ;
    END
  END reg1_val1[28]
  PIN reg1_val1[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 656.920 2200.000 657.520 ;
    END
  END reg1_val1[29]
  PIN reg1_val1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 583.480 2200.000 584.080 ;
    END
  END reg1_val1[2]
  PIN reg1_val1[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 659.640 2200.000 660.240 ;
    END
  END reg1_val1[30]
  PIN reg1_val1[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 662.360 2200.000 662.960 ;
    END
  END reg1_val1[31]
  PIN reg1_val1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 586.200 2200.000 586.800 ;
    END
  END reg1_val1[3]
  PIN reg1_val1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 588.920 2200.000 589.520 ;
    END
  END reg1_val1[4]
  PIN reg1_val1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 591.640 2200.000 592.240 ;
    END
  END reg1_val1[5]
  PIN reg1_val1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 594.360 2200.000 594.960 ;
    END
  END reg1_val1[6]
  PIN reg1_val1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 597.080 2200.000 597.680 ;
    END
  END reg1_val1[7]
  PIN reg1_val1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 599.800 2200.000 600.400 ;
    END
  END reg1_val1[8]
  PIN reg1_val1[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 602.520 2200.000 603.120 ;
    END
  END reg1_val1[9]
  PIN reg1_val2[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 572.600 4.000 573.200 ;
    END
  END reg1_val2[0]
  PIN reg1_val2[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 599.800 4.000 600.400 ;
    END
  END reg1_val2[10]
  PIN reg1_val2[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 602.520 4.000 603.120 ;
    END
  END reg1_val2[11]
  PIN reg1_val2[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 605.240 4.000 605.840 ;
    END
  END reg1_val2[12]
  PIN reg1_val2[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 607.960 4.000 608.560 ;
    END
  END reg1_val2[13]
  PIN reg1_val2[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 610.680 4.000 611.280 ;
    END
  END reg1_val2[14]
  PIN reg1_val2[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 613.400 4.000 614.000 ;
    END
  END reg1_val2[15]
  PIN reg1_val2[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 616.120 4.000 616.720 ;
    END
  END reg1_val2[16]
  PIN reg1_val2[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 618.840 4.000 619.440 ;
    END
  END reg1_val2[17]
  PIN reg1_val2[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 621.560 4.000 622.160 ;
    END
  END reg1_val2[18]
  PIN reg1_val2[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 624.280 4.000 624.880 ;
    END
  END reg1_val2[19]
  PIN reg1_val2[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 575.320 4.000 575.920 ;
    END
  END reg1_val2[1]
  PIN reg1_val2[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 627.000 4.000 627.600 ;
    END
  END reg1_val2[20]
  PIN reg1_val2[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 629.720 4.000 630.320 ;
    END
  END reg1_val2[21]
  PIN reg1_val2[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 632.440 4.000 633.040 ;
    END
  END reg1_val2[22]
  PIN reg1_val2[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 635.160 4.000 635.760 ;
    END
  END reg1_val2[23]
  PIN reg1_val2[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 637.880 4.000 638.480 ;
    END
  END reg1_val2[24]
  PIN reg1_val2[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 640.600 4.000 641.200 ;
    END
  END reg1_val2[25]
  PIN reg1_val2[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 643.320 4.000 643.920 ;
    END
  END reg1_val2[26]
  PIN reg1_val2[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 646.040 4.000 646.640 ;
    END
  END reg1_val2[27]
  PIN reg1_val2[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 648.760 4.000 649.360 ;
    END
  END reg1_val2[28]
  PIN reg1_val2[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 651.480 4.000 652.080 ;
    END
  END reg1_val2[29]
  PIN reg1_val2[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 578.040 4.000 578.640 ;
    END
  END reg1_val2[2]
  PIN reg1_val2[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 654.200 4.000 654.800 ;
    END
  END reg1_val2[30]
  PIN reg1_val2[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 656.920 4.000 657.520 ;
    END
  END reg1_val2[31]
  PIN reg1_val2[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 580.760 4.000 581.360 ;
    END
  END reg1_val2[3]
  PIN reg1_val2[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 583.480 4.000 584.080 ;
    END
  END reg1_val2[4]
  PIN reg1_val2[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 586.200 4.000 586.800 ;
    END
  END reg1_val2[5]
  PIN reg1_val2[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 588.920 4.000 589.520 ;
    END
  END reg1_val2[6]
  PIN reg1_val2[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 591.640 4.000 592.240 ;
    END
  END reg1_val2[7]
  PIN reg1_val2[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 594.360 4.000 594.960 ;
    END
  END reg1_val2[8]
  PIN reg1_val2[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 597.080 4.000 597.680 ;
    END
  END reg1_val2[9]
  PIN reg2_idx0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.436500 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met2 ;
        RECT 993.230 846.000 993.510 850.000 ;
    END
  END reg2_idx0[0]
  PIN reg2_idx0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.970000 ;
    PORT
      LAYER met2 ;
        RECT 998.290 846.000 998.570 850.000 ;
    END
  END reg2_idx0[1]
  PIN reg2_idx0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 1003.350 846.000 1003.630 850.000 ;
    END
  END reg2_idx0[2]
  PIN reg2_idx0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.960000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1008.410 846.000 1008.690 850.000 ;
    END
  END reg2_idx0[3]
  PIN reg2_idx0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.722500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1013.470 846.000 1013.750 850.000 ;
    END
  END reg2_idx0[4]
  PIN reg2_idx0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 1018.530 846.000 1018.810 850.000 ;
    END
  END reg2_idx0[5]
  PIN reg2_idx1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 121.080 2200.000 121.680 ;
    END
  END reg2_idx1[0]
  PIN reg2_idx1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.722500 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 123.800 2200.000 124.400 ;
    END
  END reg2_idx1[1]
  PIN reg2_idx1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.574500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 126.520 2200.000 127.120 ;
    END
  END reg2_idx1[2]
  PIN reg2_idx1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.574500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 129.240 2200.000 129.840 ;
    END
  END reg2_idx1[3]
  PIN reg2_idx1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.722500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 131.960 2200.000 132.560 ;
    END
  END reg2_idx1[4]
  PIN reg2_idx1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.980000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 134.680 2200.000 135.280 ;
    END
  END reg2_idx1[5]
  PIN reg2_idx2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.426500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END reg2_idx2[0]
  PIN reg2_idx2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.360 4.000 118.960 ;
    END
  END reg2_idx2[1]
  PIN reg2_idx2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.080 4.000 121.680 ;
    END
  END reg2_idx2[2]
  PIN reg2_idx2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.059500 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.800 4.000 124.400 ;
    END
  END reg2_idx2[3]
  PIN reg2_idx2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.793000 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.520 4.000 127.120 ;
    END
  END reg2_idx2[4]
  PIN reg2_idx2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END reg2_idx2[5]
  PIN reg2_val0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 2005.230 846.000 2005.510 850.000 ;
    END
  END reg2_val0[0]
  PIN reg2_val0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 2055.830 846.000 2056.110 850.000 ;
    END
  END reg2_val0[10]
  PIN reg2_val0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 2060.890 846.000 2061.170 850.000 ;
    END
  END reg2_val0[11]
  PIN reg2_val0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 2065.950 846.000 2066.230 850.000 ;
    END
  END reg2_val0[12]
  PIN reg2_val0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 2071.010 846.000 2071.290 850.000 ;
    END
  END reg2_val0[13]
  PIN reg2_val0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 2076.070 846.000 2076.350 850.000 ;
    END
  END reg2_val0[14]
  PIN reg2_val0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 2081.130 846.000 2081.410 850.000 ;
    END
  END reg2_val0[15]
  PIN reg2_val0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 2086.190 846.000 2086.470 850.000 ;
    END
  END reg2_val0[16]
  PIN reg2_val0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 2091.250 846.000 2091.530 850.000 ;
    END
  END reg2_val0[17]
  PIN reg2_val0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 2096.310 846.000 2096.590 850.000 ;
    END
  END reg2_val0[18]
  PIN reg2_val0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 2101.370 846.000 2101.650 850.000 ;
    END
  END reg2_val0[19]
  PIN reg2_val0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 2010.290 846.000 2010.570 850.000 ;
    END
  END reg2_val0[1]
  PIN reg2_val0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 2106.430 846.000 2106.710 850.000 ;
    END
  END reg2_val0[20]
  PIN reg2_val0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 2111.490 846.000 2111.770 850.000 ;
    END
  END reg2_val0[21]
  PIN reg2_val0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 2116.550 846.000 2116.830 850.000 ;
    END
  END reg2_val0[22]
  PIN reg2_val0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 2121.610 846.000 2121.890 850.000 ;
    END
  END reg2_val0[23]
  PIN reg2_val0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 2126.670 846.000 2126.950 850.000 ;
    END
  END reg2_val0[24]
  PIN reg2_val0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 2131.730 846.000 2132.010 850.000 ;
    END
  END reg2_val0[25]
  PIN reg2_val0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 2136.790 846.000 2137.070 850.000 ;
    END
  END reg2_val0[26]
  PIN reg2_val0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 2141.850 846.000 2142.130 850.000 ;
    END
  END reg2_val0[27]
  PIN reg2_val0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 2146.910 846.000 2147.190 850.000 ;
    END
  END reg2_val0[28]
  PIN reg2_val0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 2151.970 846.000 2152.250 850.000 ;
    END
  END reg2_val0[29]
  PIN reg2_val0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 2015.350 846.000 2015.630 850.000 ;
    END
  END reg2_val0[2]
  PIN reg2_val0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 2157.030 846.000 2157.310 850.000 ;
    END
  END reg2_val0[30]
  PIN reg2_val0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 2162.090 846.000 2162.370 850.000 ;
    END
  END reg2_val0[31]
  PIN reg2_val0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 2020.410 846.000 2020.690 850.000 ;
    END
  END reg2_val0[3]
  PIN reg2_val0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 2025.470 846.000 2025.750 850.000 ;
    END
  END reg2_val0[4]
  PIN reg2_val0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 2030.530 846.000 2030.810 850.000 ;
    END
  END reg2_val0[5]
  PIN reg2_val0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 2035.590 846.000 2035.870 850.000 ;
    END
  END reg2_val0[6]
  PIN reg2_val0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 2040.650 846.000 2040.930 850.000 ;
    END
  END reg2_val0[7]
  PIN reg2_val0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 2045.710 846.000 2045.990 850.000 ;
    END
  END reg2_val0[8]
  PIN reg2_val0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 2050.770 846.000 2051.050 850.000 ;
    END
  END reg2_val0[9]
  PIN reg2_val1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 665.080 2200.000 665.680 ;
    END
  END reg2_val1[0]
  PIN reg2_val1[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 692.280 2200.000 692.880 ;
    END
  END reg2_val1[10]
  PIN reg2_val1[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 695.000 2200.000 695.600 ;
    END
  END reg2_val1[11]
  PIN reg2_val1[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 697.720 2200.000 698.320 ;
    END
  END reg2_val1[12]
  PIN reg2_val1[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 700.440 2200.000 701.040 ;
    END
  END reg2_val1[13]
  PIN reg2_val1[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 703.160 2200.000 703.760 ;
    END
  END reg2_val1[14]
  PIN reg2_val1[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 705.880 2200.000 706.480 ;
    END
  END reg2_val1[15]
  PIN reg2_val1[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 708.600 2200.000 709.200 ;
    END
  END reg2_val1[16]
  PIN reg2_val1[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 711.320 2200.000 711.920 ;
    END
  END reg2_val1[17]
  PIN reg2_val1[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 714.040 2200.000 714.640 ;
    END
  END reg2_val1[18]
  PIN reg2_val1[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 716.760 2200.000 717.360 ;
    END
  END reg2_val1[19]
  PIN reg2_val1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 667.800 2200.000 668.400 ;
    END
  END reg2_val1[1]
  PIN reg2_val1[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 719.480 2200.000 720.080 ;
    END
  END reg2_val1[20]
  PIN reg2_val1[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 722.200 2200.000 722.800 ;
    END
  END reg2_val1[21]
  PIN reg2_val1[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 724.920 2200.000 725.520 ;
    END
  END reg2_val1[22]
  PIN reg2_val1[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 727.640 2200.000 728.240 ;
    END
  END reg2_val1[23]
  PIN reg2_val1[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 730.360 2200.000 730.960 ;
    END
  END reg2_val1[24]
  PIN reg2_val1[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 733.080 2200.000 733.680 ;
    END
  END reg2_val1[25]
  PIN reg2_val1[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 735.800 2200.000 736.400 ;
    END
  END reg2_val1[26]
  PIN reg2_val1[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 738.520 2200.000 739.120 ;
    END
  END reg2_val1[27]
  PIN reg2_val1[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 741.240 2200.000 741.840 ;
    END
  END reg2_val1[28]
  PIN reg2_val1[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 743.960 2200.000 744.560 ;
    END
  END reg2_val1[29]
  PIN reg2_val1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 670.520 2200.000 671.120 ;
    END
  END reg2_val1[2]
  PIN reg2_val1[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 746.680 2200.000 747.280 ;
    END
  END reg2_val1[30]
  PIN reg2_val1[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 749.400 2200.000 750.000 ;
    END
  END reg2_val1[31]
  PIN reg2_val1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 673.240 2200.000 673.840 ;
    END
  END reg2_val1[3]
  PIN reg2_val1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 675.960 2200.000 676.560 ;
    END
  END reg2_val1[4]
  PIN reg2_val1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 678.680 2200.000 679.280 ;
    END
  END reg2_val1[5]
  PIN reg2_val1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 681.400 2200.000 682.000 ;
    END
  END reg2_val1[6]
  PIN reg2_val1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 684.120 2200.000 684.720 ;
    END
  END reg2_val1[7]
  PIN reg2_val1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 686.840 2200.000 687.440 ;
    END
  END reg2_val1[8]
  PIN reg2_val1[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 689.560 2200.000 690.160 ;
    END
  END reg2_val1[9]
  PIN reg2_val2[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 659.640 4.000 660.240 ;
    END
  END reg2_val2[0]
  PIN reg2_val2[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 686.840 4.000 687.440 ;
    END
  END reg2_val2[10]
  PIN reg2_val2[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 689.560 4.000 690.160 ;
    END
  END reg2_val2[11]
  PIN reg2_val2[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 692.280 4.000 692.880 ;
    END
  END reg2_val2[12]
  PIN reg2_val2[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 695.000 4.000 695.600 ;
    END
  END reg2_val2[13]
  PIN reg2_val2[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 697.720 4.000 698.320 ;
    END
  END reg2_val2[14]
  PIN reg2_val2[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 700.440 4.000 701.040 ;
    END
  END reg2_val2[15]
  PIN reg2_val2[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 703.160 4.000 703.760 ;
    END
  END reg2_val2[16]
  PIN reg2_val2[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 705.880 4.000 706.480 ;
    END
  END reg2_val2[17]
  PIN reg2_val2[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 708.600 4.000 709.200 ;
    END
  END reg2_val2[18]
  PIN reg2_val2[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 711.320 4.000 711.920 ;
    END
  END reg2_val2[19]
  PIN reg2_val2[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 662.360 4.000 662.960 ;
    END
  END reg2_val2[1]
  PIN reg2_val2[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 714.040 4.000 714.640 ;
    END
  END reg2_val2[20]
  PIN reg2_val2[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 716.760 4.000 717.360 ;
    END
  END reg2_val2[21]
  PIN reg2_val2[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 719.480 4.000 720.080 ;
    END
  END reg2_val2[22]
  PIN reg2_val2[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 722.200 4.000 722.800 ;
    END
  END reg2_val2[23]
  PIN reg2_val2[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 724.920 4.000 725.520 ;
    END
  END reg2_val2[24]
  PIN reg2_val2[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 727.640 4.000 728.240 ;
    END
  END reg2_val2[25]
  PIN reg2_val2[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 730.360 4.000 730.960 ;
    END
  END reg2_val2[26]
  PIN reg2_val2[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 733.080 4.000 733.680 ;
    END
  END reg2_val2[27]
  PIN reg2_val2[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 735.800 4.000 736.400 ;
    END
  END reg2_val2[28]
  PIN reg2_val2[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 738.520 4.000 739.120 ;
    END
  END reg2_val2[29]
  PIN reg2_val2[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 665.080 4.000 665.680 ;
    END
  END reg2_val2[2]
  PIN reg2_val2[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 741.240 4.000 741.840 ;
    END
  END reg2_val2[30]
  PIN reg2_val2[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 743.960 4.000 744.560 ;
    END
  END reg2_val2[31]
  PIN reg2_val2[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 667.800 4.000 668.400 ;
    END
  END reg2_val2[3]
  PIN reg2_val2[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 670.520 4.000 671.120 ;
    END
  END reg2_val2[4]
  PIN reg2_val2[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 673.240 4.000 673.840 ;
    END
  END reg2_val2[5]
  PIN reg2_val2[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 675.960 4.000 676.560 ;
    END
  END reg2_val2[6]
  PIN reg2_val2[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 678.680 4.000 679.280 ;
    END
  END reg2_val2[7]
  PIN reg2_val2[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 681.400 4.000 682.000 ;
    END
  END reg2_val2[8]
  PIN reg2_val2[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 684.120 4.000 684.720 ;
    END
  END reg2_val2[9]
  PIN rst_eu
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.862000 ;
    PORT
      LAYER met2 ;
        RECT 816.130 846.000 816.410 850.000 ;
    END
  END rst_eu
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.086000 ;
    PORT
      LAYER met2 ;
        RECT 2113.330 0.000 2113.610 4.000 ;
    END
  END rst_n
  PIN sign_extend0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 2.608200 ;
    PORT
      LAYER met2 ;
        RECT 1433.450 846.000 1433.730 850.000 ;
    END
  END sign_extend0
  PIN sign_extend1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 357.720 2200.000 358.320 ;
    END
  END sign_extend1
  PIN sign_extend2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 7.824600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 352.280 4.000 352.880 ;
    END
  END sign_extend2
  PIN take_branch0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.227500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1478.990 846.000 1479.270 850.000 ;
    END
  END take_branch0
  PIN take_branch1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 7.996500 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 382.200 2200.000 382.800 ;
    END
  END take_branch1
  PIN take_branch2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.475000 ;
    ANTENNADIFFAREA 2.173500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 376.760 4.000 377.360 ;
    END
  END take_branch2
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 838.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 838.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 838.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 838.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 838.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 838.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 838.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 838.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 838.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 838.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.040 10.640 1558.640 838.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1710.640 10.640 1712.240 838.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1864.240 10.640 1865.840 838.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2017.840 10.640 2019.440 838.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2171.440 10.640 2173.040 838.000 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 838.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 838.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 838.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 838.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 838.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 838.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 838.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 838.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 838.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 838.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1633.840 10.640 1635.440 838.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1787.440 10.640 1789.040 838.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1941.040 10.640 1942.640 838.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2094.640 10.640 2096.240 838.000 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 2104.590 0.000 2104.870 4.000 ;
    END
  END wb_clk_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2194.200 837.845 ;
      LAYER met1 ;
        RECT 5.520 0.380 2196.890 849.960 ;
      LAYER met2 ;
        RECT 6.070 845.720 26.490 849.990 ;
        RECT 27.330 845.720 31.550 849.990 ;
        RECT 32.390 845.720 36.610 849.990 ;
        RECT 37.450 845.720 41.670 849.990 ;
        RECT 42.510 845.720 46.730 849.990 ;
        RECT 47.570 845.720 51.790 849.990 ;
        RECT 52.630 845.720 56.850 849.990 ;
        RECT 57.690 845.720 61.910 849.990 ;
        RECT 62.750 845.720 66.970 849.990 ;
        RECT 67.810 845.720 72.030 849.990 ;
        RECT 72.870 845.720 77.090 849.990 ;
        RECT 77.930 845.720 82.150 849.990 ;
        RECT 82.990 845.720 87.210 849.990 ;
        RECT 88.050 845.720 92.270 849.990 ;
        RECT 93.110 845.720 97.330 849.990 ;
        RECT 98.170 845.720 102.390 849.990 ;
        RECT 103.230 845.720 107.450 849.990 ;
        RECT 108.290 845.720 112.510 849.990 ;
        RECT 113.350 845.720 117.570 849.990 ;
        RECT 118.410 845.720 122.630 849.990 ;
        RECT 123.470 845.720 127.690 849.990 ;
        RECT 128.530 845.720 132.750 849.990 ;
        RECT 133.590 845.720 137.810 849.990 ;
        RECT 138.650 845.720 142.870 849.990 ;
        RECT 143.710 845.720 147.930 849.990 ;
        RECT 148.770 845.720 152.990 849.990 ;
        RECT 153.830 845.720 158.050 849.990 ;
        RECT 158.890 845.720 163.110 849.990 ;
        RECT 163.950 845.720 168.170 849.990 ;
        RECT 169.010 845.720 173.230 849.990 ;
        RECT 174.070 845.720 178.290 849.990 ;
        RECT 179.130 845.720 183.350 849.990 ;
        RECT 184.190 845.720 188.410 849.990 ;
        RECT 189.250 845.720 193.470 849.990 ;
        RECT 194.310 845.720 198.530 849.990 ;
        RECT 199.370 845.720 203.590 849.990 ;
        RECT 204.430 845.720 208.650 849.990 ;
        RECT 209.490 845.720 213.710 849.990 ;
        RECT 214.550 845.720 218.770 849.990 ;
        RECT 219.610 845.720 223.830 849.990 ;
        RECT 224.670 845.720 228.890 849.990 ;
        RECT 229.730 845.720 233.950 849.990 ;
        RECT 234.790 845.720 239.010 849.990 ;
        RECT 239.850 845.720 244.070 849.990 ;
        RECT 244.910 845.720 249.130 849.990 ;
        RECT 249.970 845.720 254.190 849.990 ;
        RECT 255.030 845.720 259.250 849.990 ;
        RECT 260.090 845.720 264.310 849.990 ;
        RECT 265.150 845.720 269.370 849.990 ;
        RECT 270.210 845.720 274.430 849.990 ;
        RECT 275.270 845.720 279.490 849.990 ;
        RECT 280.330 845.720 284.550 849.990 ;
        RECT 285.390 845.720 289.610 849.990 ;
        RECT 290.450 845.720 294.670 849.990 ;
        RECT 295.510 845.720 299.730 849.990 ;
        RECT 300.570 845.720 304.790 849.990 ;
        RECT 305.630 845.720 309.850 849.990 ;
        RECT 310.690 845.720 314.910 849.990 ;
        RECT 315.750 845.720 319.970 849.990 ;
        RECT 320.810 845.720 325.030 849.990 ;
        RECT 325.870 845.720 330.090 849.990 ;
        RECT 330.930 845.720 335.150 849.990 ;
        RECT 335.990 845.720 340.210 849.990 ;
        RECT 341.050 845.720 345.270 849.990 ;
        RECT 346.110 845.720 350.330 849.990 ;
        RECT 351.170 845.720 355.390 849.990 ;
        RECT 356.230 845.720 360.450 849.990 ;
        RECT 361.290 845.720 365.510 849.990 ;
        RECT 366.350 845.720 370.570 849.990 ;
        RECT 371.410 845.720 375.630 849.990 ;
        RECT 376.470 845.720 380.690 849.990 ;
        RECT 381.530 845.720 385.750 849.990 ;
        RECT 386.590 845.720 390.810 849.990 ;
        RECT 391.650 845.720 395.870 849.990 ;
        RECT 396.710 845.720 400.930 849.990 ;
        RECT 401.770 845.720 405.990 849.990 ;
        RECT 406.830 845.720 411.050 849.990 ;
        RECT 411.890 845.720 416.110 849.990 ;
        RECT 416.950 845.720 421.170 849.990 ;
        RECT 422.010 845.720 426.230 849.990 ;
        RECT 427.070 845.720 431.290 849.990 ;
        RECT 432.130 845.720 436.350 849.990 ;
        RECT 437.190 845.720 441.410 849.990 ;
        RECT 442.250 845.720 446.470 849.990 ;
        RECT 447.310 845.720 451.530 849.990 ;
        RECT 452.370 845.720 456.590 849.990 ;
        RECT 457.430 845.720 461.650 849.990 ;
        RECT 462.490 845.720 466.710 849.990 ;
        RECT 467.550 845.720 471.770 849.990 ;
        RECT 472.610 845.720 476.830 849.990 ;
        RECT 477.670 845.720 481.890 849.990 ;
        RECT 482.730 845.720 486.950 849.990 ;
        RECT 487.790 845.720 492.010 849.990 ;
        RECT 492.850 845.720 497.070 849.990 ;
        RECT 497.910 845.720 502.130 849.990 ;
        RECT 502.970 845.720 507.190 849.990 ;
        RECT 508.030 845.720 512.250 849.990 ;
        RECT 513.090 845.720 517.310 849.990 ;
        RECT 518.150 845.720 522.370 849.990 ;
        RECT 523.210 845.720 527.430 849.990 ;
        RECT 528.270 845.720 532.490 849.990 ;
        RECT 533.330 845.720 537.550 849.990 ;
        RECT 538.390 845.720 542.610 849.990 ;
        RECT 543.450 845.720 547.670 849.990 ;
        RECT 548.510 845.720 552.730 849.990 ;
        RECT 553.570 845.720 557.790 849.990 ;
        RECT 558.630 845.720 562.850 849.990 ;
        RECT 563.690 845.720 567.910 849.990 ;
        RECT 568.750 845.720 572.970 849.990 ;
        RECT 573.810 845.720 578.030 849.990 ;
        RECT 578.870 845.720 583.090 849.990 ;
        RECT 583.930 845.720 588.150 849.990 ;
        RECT 588.990 845.720 593.210 849.990 ;
        RECT 594.050 845.720 598.270 849.990 ;
        RECT 599.110 845.720 603.330 849.990 ;
        RECT 604.170 845.720 608.390 849.990 ;
        RECT 609.230 845.720 613.450 849.990 ;
        RECT 614.290 845.720 618.510 849.990 ;
        RECT 619.350 845.720 623.570 849.990 ;
        RECT 624.410 845.720 628.630 849.990 ;
        RECT 629.470 845.720 633.690 849.990 ;
        RECT 634.530 845.720 638.750 849.990 ;
        RECT 639.590 845.720 643.810 849.990 ;
        RECT 644.650 845.720 648.870 849.990 ;
        RECT 649.710 845.720 653.930 849.990 ;
        RECT 654.770 845.720 658.990 849.990 ;
        RECT 659.830 845.720 664.050 849.990 ;
        RECT 664.890 845.720 669.110 849.990 ;
        RECT 669.950 845.720 674.170 849.990 ;
        RECT 675.010 845.720 679.230 849.990 ;
        RECT 680.070 845.720 684.290 849.990 ;
        RECT 685.130 845.720 689.350 849.990 ;
        RECT 690.190 845.720 694.410 849.990 ;
        RECT 695.250 845.720 699.470 849.990 ;
        RECT 700.310 845.720 704.530 849.990 ;
        RECT 705.370 845.720 709.590 849.990 ;
        RECT 710.430 845.720 714.650 849.990 ;
        RECT 715.490 845.720 719.710 849.990 ;
        RECT 720.550 845.720 724.770 849.990 ;
        RECT 725.610 845.720 729.830 849.990 ;
        RECT 730.670 845.720 734.890 849.990 ;
        RECT 735.730 845.720 739.950 849.990 ;
        RECT 740.790 845.720 745.010 849.990 ;
        RECT 745.850 845.720 750.070 849.990 ;
        RECT 750.910 845.720 755.130 849.990 ;
        RECT 755.970 845.720 760.190 849.990 ;
        RECT 761.030 845.720 765.250 849.990 ;
        RECT 766.090 845.720 770.310 849.990 ;
        RECT 771.150 845.720 775.370 849.990 ;
        RECT 776.210 845.720 780.430 849.990 ;
        RECT 781.270 845.720 785.490 849.990 ;
        RECT 786.330 845.720 790.550 849.990 ;
        RECT 791.390 845.720 795.610 849.990 ;
        RECT 796.450 845.720 800.670 849.990 ;
        RECT 801.510 845.720 805.730 849.990 ;
        RECT 806.570 845.720 810.790 849.990 ;
        RECT 811.630 845.720 815.850 849.990 ;
        RECT 816.690 845.720 820.910 849.990 ;
        RECT 821.750 845.720 825.970 849.990 ;
        RECT 826.810 845.720 831.030 849.990 ;
        RECT 831.870 845.720 836.090 849.990 ;
        RECT 836.930 845.720 841.150 849.990 ;
        RECT 841.990 845.720 846.210 849.990 ;
        RECT 847.050 845.720 851.270 849.990 ;
        RECT 852.110 845.720 856.330 849.990 ;
        RECT 857.170 845.720 861.390 849.990 ;
        RECT 862.230 845.720 866.450 849.990 ;
        RECT 867.290 845.720 871.510 849.990 ;
        RECT 872.350 845.720 876.570 849.990 ;
        RECT 877.410 845.720 881.630 849.990 ;
        RECT 882.470 845.720 886.690 849.990 ;
        RECT 887.530 845.720 891.750 849.990 ;
        RECT 892.590 845.720 896.810 849.990 ;
        RECT 897.650 845.720 901.870 849.990 ;
        RECT 902.710 845.720 906.930 849.990 ;
        RECT 907.770 845.720 911.990 849.990 ;
        RECT 912.830 845.720 917.050 849.990 ;
        RECT 917.890 845.720 922.110 849.990 ;
        RECT 922.950 845.720 927.170 849.990 ;
        RECT 928.010 845.720 932.230 849.990 ;
        RECT 933.070 845.720 937.290 849.990 ;
        RECT 938.130 845.720 942.350 849.990 ;
        RECT 943.190 845.720 947.410 849.990 ;
        RECT 948.250 845.720 952.470 849.990 ;
        RECT 953.310 845.720 957.530 849.990 ;
        RECT 958.370 845.720 962.590 849.990 ;
        RECT 963.430 845.720 967.650 849.990 ;
        RECT 968.490 845.720 972.710 849.990 ;
        RECT 973.550 845.720 977.770 849.990 ;
        RECT 978.610 845.720 982.830 849.990 ;
        RECT 983.670 845.720 987.890 849.990 ;
        RECT 988.730 845.720 992.950 849.990 ;
        RECT 993.790 845.720 998.010 849.990 ;
        RECT 998.850 845.720 1003.070 849.990 ;
        RECT 1003.910 845.720 1008.130 849.990 ;
        RECT 1008.970 845.720 1013.190 849.990 ;
        RECT 1014.030 845.720 1018.250 849.990 ;
        RECT 1019.090 845.720 1023.310 849.990 ;
        RECT 1024.150 845.720 1028.370 849.990 ;
        RECT 1029.210 845.720 1033.430 849.990 ;
        RECT 1034.270 845.720 1038.490 849.990 ;
        RECT 1039.330 845.720 1043.550 849.990 ;
        RECT 1044.390 845.720 1048.610 849.990 ;
        RECT 1049.450 845.720 1053.670 849.990 ;
        RECT 1054.510 845.720 1058.730 849.990 ;
        RECT 1059.570 845.720 1063.790 849.990 ;
        RECT 1064.630 845.720 1068.850 849.990 ;
        RECT 1069.690 845.720 1073.910 849.990 ;
        RECT 1074.750 845.720 1078.970 849.990 ;
        RECT 1079.810 845.720 1084.030 849.990 ;
        RECT 1084.870 845.720 1089.090 849.990 ;
        RECT 1089.930 845.720 1094.150 849.990 ;
        RECT 1094.990 845.720 1099.210 849.990 ;
        RECT 1100.050 845.720 1104.270 849.990 ;
        RECT 1105.110 845.720 1109.330 849.990 ;
        RECT 1110.170 845.720 1114.390 849.990 ;
        RECT 1115.230 845.720 1119.450 849.990 ;
        RECT 1120.290 845.720 1124.510 849.990 ;
        RECT 1125.350 845.720 1129.570 849.990 ;
        RECT 1130.410 845.720 1134.630 849.990 ;
        RECT 1135.470 845.720 1139.690 849.990 ;
        RECT 1140.530 845.720 1144.750 849.990 ;
        RECT 1145.590 845.720 1149.810 849.990 ;
        RECT 1150.650 845.720 1154.870 849.990 ;
        RECT 1155.710 845.720 1159.930 849.990 ;
        RECT 1160.770 845.720 1164.990 849.990 ;
        RECT 1165.830 845.720 1170.050 849.990 ;
        RECT 1170.890 845.720 1175.110 849.990 ;
        RECT 1175.950 845.720 1180.170 849.990 ;
        RECT 1181.010 845.720 1185.230 849.990 ;
        RECT 1186.070 845.720 1190.290 849.990 ;
        RECT 1191.130 845.720 1195.350 849.990 ;
        RECT 1196.190 845.720 1200.410 849.990 ;
        RECT 1201.250 845.720 1205.470 849.990 ;
        RECT 1206.310 845.720 1210.530 849.990 ;
        RECT 1211.370 845.720 1215.590 849.990 ;
        RECT 1216.430 845.720 1220.650 849.990 ;
        RECT 1221.490 845.720 1225.710 849.990 ;
        RECT 1226.550 845.720 1230.770 849.990 ;
        RECT 1231.610 845.720 1235.830 849.990 ;
        RECT 1236.670 845.720 1240.890 849.990 ;
        RECT 1241.730 845.720 1245.950 849.990 ;
        RECT 1246.790 845.720 1251.010 849.990 ;
        RECT 1251.850 845.720 1256.070 849.990 ;
        RECT 1256.910 845.720 1261.130 849.990 ;
        RECT 1261.970 845.720 1266.190 849.990 ;
        RECT 1267.030 845.720 1271.250 849.990 ;
        RECT 1272.090 845.720 1276.310 849.990 ;
        RECT 1277.150 845.720 1281.370 849.990 ;
        RECT 1282.210 845.720 1286.430 849.990 ;
        RECT 1287.270 845.720 1291.490 849.990 ;
        RECT 1292.330 845.720 1296.550 849.990 ;
        RECT 1297.390 845.720 1301.610 849.990 ;
        RECT 1302.450 845.720 1306.670 849.990 ;
        RECT 1307.510 845.720 1311.730 849.990 ;
        RECT 1312.570 845.720 1316.790 849.990 ;
        RECT 1317.630 845.720 1321.850 849.990 ;
        RECT 1322.690 845.720 1326.910 849.990 ;
        RECT 1327.750 845.720 1331.970 849.990 ;
        RECT 1332.810 845.720 1337.030 849.990 ;
        RECT 1337.870 845.720 1342.090 849.990 ;
        RECT 1342.930 845.720 1347.150 849.990 ;
        RECT 1347.990 845.720 1352.210 849.990 ;
        RECT 1353.050 845.720 1357.270 849.990 ;
        RECT 1358.110 845.720 1362.330 849.990 ;
        RECT 1363.170 845.720 1367.390 849.990 ;
        RECT 1368.230 845.720 1372.450 849.990 ;
        RECT 1373.290 845.720 1377.510 849.990 ;
        RECT 1378.350 845.720 1382.570 849.990 ;
        RECT 1383.410 845.720 1387.630 849.990 ;
        RECT 1388.470 845.720 1392.690 849.990 ;
        RECT 1393.530 845.720 1397.750 849.990 ;
        RECT 1398.590 845.720 1402.810 849.990 ;
        RECT 1403.650 845.720 1407.870 849.990 ;
        RECT 1408.710 845.720 1412.930 849.990 ;
        RECT 1413.770 845.720 1417.990 849.990 ;
        RECT 1418.830 845.720 1423.050 849.990 ;
        RECT 1423.890 845.720 1428.110 849.990 ;
        RECT 1428.950 845.720 1433.170 849.990 ;
        RECT 1434.010 845.720 1438.230 849.990 ;
        RECT 1439.070 845.720 1443.290 849.990 ;
        RECT 1444.130 845.720 1448.350 849.990 ;
        RECT 1449.190 845.720 1453.410 849.990 ;
        RECT 1454.250 845.720 1458.470 849.990 ;
        RECT 1459.310 845.720 1463.530 849.990 ;
        RECT 1464.370 845.720 1468.590 849.990 ;
        RECT 1469.430 845.720 1473.650 849.990 ;
        RECT 1474.490 845.720 1478.710 849.990 ;
        RECT 1479.550 845.720 1483.770 849.990 ;
        RECT 1484.610 845.720 1488.830 849.990 ;
        RECT 1489.670 845.720 1493.890 849.990 ;
        RECT 1494.730 845.720 1498.950 849.990 ;
        RECT 1499.790 845.720 1504.010 849.990 ;
        RECT 1504.850 845.720 1509.070 849.990 ;
        RECT 1509.910 845.720 1514.130 849.990 ;
        RECT 1514.970 845.720 1519.190 849.990 ;
        RECT 1520.030 845.720 1524.250 849.990 ;
        RECT 1525.090 845.720 1529.310 849.990 ;
        RECT 1530.150 845.720 1534.370 849.990 ;
        RECT 1535.210 845.720 1539.430 849.990 ;
        RECT 1540.270 845.720 1544.490 849.990 ;
        RECT 1545.330 845.720 1549.550 849.990 ;
        RECT 1550.390 845.720 1554.610 849.990 ;
        RECT 1555.450 845.720 1559.670 849.990 ;
        RECT 1560.510 845.720 1564.730 849.990 ;
        RECT 1565.570 845.720 1569.790 849.990 ;
        RECT 1570.630 845.720 1574.850 849.990 ;
        RECT 1575.690 845.720 1579.910 849.990 ;
        RECT 1580.750 845.720 1584.970 849.990 ;
        RECT 1585.810 845.720 1590.030 849.990 ;
        RECT 1590.870 845.720 1595.090 849.990 ;
        RECT 1595.930 845.720 1600.150 849.990 ;
        RECT 1600.990 845.720 1605.210 849.990 ;
        RECT 1606.050 845.720 1610.270 849.990 ;
        RECT 1611.110 845.720 1615.330 849.990 ;
        RECT 1616.170 845.720 1620.390 849.990 ;
        RECT 1621.230 845.720 1625.450 849.990 ;
        RECT 1626.290 845.720 1630.510 849.990 ;
        RECT 1631.350 845.720 1635.570 849.990 ;
        RECT 1636.410 845.720 1640.630 849.990 ;
        RECT 1641.470 845.720 1645.690 849.990 ;
        RECT 1646.530 845.720 1650.750 849.990 ;
        RECT 1651.590 845.720 1655.810 849.990 ;
        RECT 1656.650 845.720 1660.870 849.990 ;
        RECT 1661.710 845.720 1665.930 849.990 ;
        RECT 1666.770 845.720 1670.990 849.990 ;
        RECT 1671.830 845.720 1676.050 849.990 ;
        RECT 1676.890 845.720 1681.110 849.990 ;
        RECT 1681.950 845.720 1686.170 849.990 ;
        RECT 1687.010 845.720 1691.230 849.990 ;
        RECT 1692.070 845.720 1696.290 849.990 ;
        RECT 1697.130 845.720 1701.350 849.990 ;
        RECT 1702.190 845.720 1706.410 849.990 ;
        RECT 1707.250 845.720 1711.470 849.990 ;
        RECT 1712.310 845.720 1716.530 849.990 ;
        RECT 1717.370 845.720 1721.590 849.990 ;
        RECT 1722.430 845.720 1726.650 849.990 ;
        RECT 1727.490 845.720 1731.710 849.990 ;
        RECT 1732.550 845.720 1736.770 849.990 ;
        RECT 1737.610 845.720 1741.830 849.990 ;
        RECT 1742.670 845.720 1746.890 849.990 ;
        RECT 1747.730 845.720 1751.950 849.990 ;
        RECT 1752.790 845.720 1757.010 849.990 ;
        RECT 1757.850 845.720 1762.070 849.990 ;
        RECT 1762.910 845.720 1767.130 849.990 ;
        RECT 1767.970 845.720 1772.190 849.990 ;
        RECT 1773.030 845.720 1777.250 849.990 ;
        RECT 1778.090 845.720 1782.310 849.990 ;
        RECT 1783.150 845.720 1787.370 849.990 ;
        RECT 1788.210 845.720 1792.430 849.990 ;
        RECT 1793.270 845.720 1797.490 849.990 ;
        RECT 1798.330 845.720 1802.550 849.990 ;
        RECT 1803.390 845.720 1807.610 849.990 ;
        RECT 1808.450 845.720 1812.670 849.990 ;
        RECT 1813.510 845.720 1817.730 849.990 ;
        RECT 1818.570 845.720 1822.790 849.990 ;
        RECT 1823.630 845.720 1827.850 849.990 ;
        RECT 1828.690 845.720 1832.910 849.990 ;
        RECT 1833.750 845.720 1837.970 849.990 ;
        RECT 1838.810 845.720 1843.030 849.990 ;
        RECT 1843.870 845.720 1848.090 849.990 ;
        RECT 1848.930 845.720 1853.150 849.990 ;
        RECT 1853.990 845.720 1858.210 849.990 ;
        RECT 1859.050 845.720 1863.270 849.990 ;
        RECT 1864.110 845.720 1868.330 849.990 ;
        RECT 1869.170 845.720 1873.390 849.990 ;
        RECT 1874.230 845.720 1878.450 849.990 ;
        RECT 1879.290 845.720 1883.510 849.990 ;
        RECT 1884.350 845.720 1888.570 849.990 ;
        RECT 1889.410 845.720 1893.630 849.990 ;
        RECT 1894.470 845.720 1898.690 849.990 ;
        RECT 1899.530 845.720 1903.750 849.990 ;
        RECT 1904.590 845.720 1908.810 849.990 ;
        RECT 1909.650 845.720 1913.870 849.990 ;
        RECT 1914.710 845.720 1918.930 849.990 ;
        RECT 1919.770 845.720 1923.990 849.990 ;
        RECT 1924.830 845.720 1929.050 849.990 ;
        RECT 1929.890 845.720 1934.110 849.990 ;
        RECT 1934.950 845.720 1939.170 849.990 ;
        RECT 1940.010 845.720 1944.230 849.990 ;
        RECT 1945.070 845.720 1949.290 849.990 ;
        RECT 1950.130 845.720 1954.350 849.990 ;
        RECT 1955.190 845.720 1959.410 849.990 ;
        RECT 1960.250 845.720 1964.470 849.990 ;
        RECT 1965.310 845.720 1969.530 849.990 ;
        RECT 1970.370 845.720 1974.590 849.990 ;
        RECT 1975.430 845.720 1979.650 849.990 ;
        RECT 1980.490 845.720 1984.710 849.990 ;
        RECT 1985.550 845.720 1989.770 849.990 ;
        RECT 1990.610 845.720 1994.830 849.990 ;
        RECT 1995.670 845.720 1999.890 849.990 ;
        RECT 2000.730 845.720 2004.950 849.990 ;
        RECT 2005.790 845.720 2010.010 849.990 ;
        RECT 2010.850 845.720 2015.070 849.990 ;
        RECT 2015.910 845.720 2020.130 849.990 ;
        RECT 2020.970 845.720 2025.190 849.990 ;
        RECT 2026.030 845.720 2030.250 849.990 ;
        RECT 2031.090 845.720 2035.310 849.990 ;
        RECT 2036.150 845.720 2040.370 849.990 ;
        RECT 2041.210 845.720 2045.430 849.990 ;
        RECT 2046.270 845.720 2050.490 849.990 ;
        RECT 2051.330 845.720 2055.550 849.990 ;
        RECT 2056.390 845.720 2060.610 849.990 ;
        RECT 2061.450 845.720 2065.670 849.990 ;
        RECT 2066.510 845.720 2070.730 849.990 ;
        RECT 2071.570 845.720 2075.790 849.990 ;
        RECT 2076.630 845.720 2080.850 849.990 ;
        RECT 2081.690 845.720 2085.910 849.990 ;
        RECT 2086.750 845.720 2090.970 849.990 ;
        RECT 2091.810 845.720 2096.030 849.990 ;
        RECT 2096.870 845.720 2101.090 849.990 ;
        RECT 2101.930 845.720 2106.150 849.990 ;
        RECT 2106.990 845.720 2111.210 849.990 ;
        RECT 2112.050 845.720 2116.270 849.990 ;
        RECT 2117.110 845.720 2121.330 849.990 ;
        RECT 2122.170 845.720 2126.390 849.990 ;
        RECT 2127.230 845.720 2131.450 849.990 ;
        RECT 2132.290 845.720 2136.510 849.990 ;
        RECT 2137.350 845.720 2141.570 849.990 ;
        RECT 2142.410 845.720 2146.630 849.990 ;
        RECT 2147.470 845.720 2151.690 849.990 ;
        RECT 2152.530 845.720 2156.750 849.990 ;
        RECT 2157.590 845.720 2161.810 849.990 ;
        RECT 2162.650 845.720 2166.870 849.990 ;
        RECT 2167.710 845.720 2171.930 849.990 ;
        RECT 2172.770 845.720 2196.860 849.990 ;
        RECT 6.070 4.280 2196.860 845.720 ;
        RECT 6.070 0.155 41.670 4.280 ;
        RECT 42.510 0.155 50.410 4.280 ;
        RECT 51.250 0.155 59.150 4.280 ;
        RECT 59.990 0.155 67.890 4.280 ;
        RECT 68.730 0.155 76.630 4.280 ;
        RECT 77.470 0.155 85.370 4.280 ;
        RECT 86.210 0.155 94.110 4.280 ;
        RECT 94.950 0.155 102.850 4.280 ;
        RECT 103.690 0.155 111.590 4.280 ;
        RECT 112.430 0.155 120.330 4.280 ;
        RECT 121.170 0.155 129.070 4.280 ;
        RECT 129.910 0.155 137.810 4.280 ;
        RECT 138.650 0.155 146.550 4.280 ;
        RECT 147.390 0.155 155.290 4.280 ;
        RECT 156.130 0.155 164.030 4.280 ;
        RECT 164.870 0.155 172.770 4.280 ;
        RECT 173.610 0.155 181.510 4.280 ;
        RECT 182.350 0.155 190.250 4.280 ;
        RECT 191.090 0.155 198.990 4.280 ;
        RECT 199.830 0.155 207.730 4.280 ;
        RECT 208.570 0.155 216.470 4.280 ;
        RECT 217.310 0.155 225.210 4.280 ;
        RECT 226.050 0.155 233.950 4.280 ;
        RECT 234.790 0.155 242.690 4.280 ;
        RECT 243.530 0.155 251.430 4.280 ;
        RECT 252.270 0.155 260.170 4.280 ;
        RECT 261.010 0.155 268.910 4.280 ;
        RECT 269.750 0.155 277.650 4.280 ;
        RECT 278.490 0.155 286.390 4.280 ;
        RECT 287.230 0.155 295.130 4.280 ;
        RECT 295.970 0.155 303.870 4.280 ;
        RECT 304.710 0.155 312.610 4.280 ;
        RECT 313.450 0.155 321.350 4.280 ;
        RECT 322.190 0.155 330.090 4.280 ;
        RECT 330.930 0.155 338.830 4.280 ;
        RECT 339.670 0.155 347.570 4.280 ;
        RECT 348.410 0.155 356.310 4.280 ;
        RECT 357.150 0.155 365.050 4.280 ;
        RECT 365.890 0.155 373.790 4.280 ;
        RECT 374.630 0.155 382.530 4.280 ;
        RECT 383.370 0.155 391.270 4.280 ;
        RECT 392.110 0.155 400.010 4.280 ;
        RECT 400.850 0.155 408.750 4.280 ;
        RECT 409.590 0.155 417.490 4.280 ;
        RECT 418.330 0.155 426.230 4.280 ;
        RECT 427.070 0.155 434.970 4.280 ;
        RECT 435.810 0.155 443.710 4.280 ;
        RECT 444.550 0.155 452.450 4.280 ;
        RECT 453.290 0.155 461.190 4.280 ;
        RECT 462.030 0.155 469.930 4.280 ;
        RECT 470.770 0.155 478.670 4.280 ;
        RECT 479.510 0.155 487.410 4.280 ;
        RECT 488.250 0.155 496.150 4.280 ;
        RECT 496.990 0.155 504.890 4.280 ;
        RECT 505.730 0.155 513.630 4.280 ;
        RECT 514.470 0.155 522.370 4.280 ;
        RECT 523.210 0.155 531.110 4.280 ;
        RECT 531.950 0.155 539.850 4.280 ;
        RECT 540.690 0.155 548.590 4.280 ;
        RECT 549.430 0.155 557.330 4.280 ;
        RECT 558.170 0.155 566.070 4.280 ;
        RECT 566.910 0.155 574.810 4.280 ;
        RECT 575.650 0.155 583.550 4.280 ;
        RECT 584.390 0.155 592.290 4.280 ;
        RECT 593.130 0.155 601.030 4.280 ;
        RECT 601.870 0.155 609.770 4.280 ;
        RECT 610.610 0.155 618.510 4.280 ;
        RECT 619.350 0.155 627.250 4.280 ;
        RECT 628.090 0.155 635.990 4.280 ;
        RECT 636.830 0.155 644.730 4.280 ;
        RECT 645.570 0.155 653.470 4.280 ;
        RECT 654.310 0.155 662.210 4.280 ;
        RECT 663.050 0.155 670.950 4.280 ;
        RECT 671.790 0.155 679.690 4.280 ;
        RECT 680.530 0.155 688.430 4.280 ;
        RECT 689.270 0.155 697.170 4.280 ;
        RECT 698.010 0.155 705.910 4.280 ;
        RECT 706.750 0.155 714.650 4.280 ;
        RECT 715.490 0.155 723.390 4.280 ;
        RECT 724.230 0.155 732.130 4.280 ;
        RECT 732.970 0.155 740.870 4.280 ;
        RECT 741.710 0.155 749.610 4.280 ;
        RECT 750.450 0.155 758.350 4.280 ;
        RECT 759.190 0.155 767.090 4.280 ;
        RECT 767.930 0.155 775.830 4.280 ;
        RECT 776.670 0.155 784.570 4.280 ;
        RECT 785.410 0.155 793.310 4.280 ;
        RECT 794.150 0.155 802.050 4.280 ;
        RECT 802.890 0.155 810.790 4.280 ;
        RECT 811.630 0.155 819.530 4.280 ;
        RECT 820.370 0.155 828.270 4.280 ;
        RECT 829.110 0.155 837.010 4.280 ;
        RECT 837.850 0.155 845.750 4.280 ;
        RECT 846.590 0.155 854.490 4.280 ;
        RECT 855.330 0.155 863.230 4.280 ;
        RECT 864.070 0.155 871.970 4.280 ;
        RECT 872.810 0.155 880.710 4.280 ;
        RECT 881.550 0.155 889.450 4.280 ;
        RECT 890.290 0.155 898.190 4.280 ;
        RECT 899.030 0.155 906.930 4.280 ;
        RECT 907.770 0.155 915.670 4.280 ;
        RECT 916.510 0.155 924.410 4.280 ;
        RECT 925.250 0.155 933.150 4.280 ;
        RECT 933.990 0.155 941.890 4.280 ;
        RECT 942.730 0.155 950.630 4.280 ;
        RECT 951.470 0.155 959.370 4.280 ;
        RECT 960.210 0.155 968.110 4.280 ;
        RECT 968.950 0.155 976.850 4.280 ;
        RECT 977.690 0.155 985.590 4.280 ;
        RECT 986.430 0.155 994.330 4.280 ;
        RECT 995.170 0.155 1003.070 4.280 ;
        RECT 1003.910 0.155 1011.810 4.280 ;
        RECT 1012.650 0.155 1020.550 4.280 ;
        RECT 1021.390 0.155 1029.290 4.280 ;
        RECT 1030.130 0.155 1038.030 4.280 ;
        RECT 1038.870 0.155 1046.770 4.280 ;
        RECT 1047.610 0.155 1055.510 4.280 ;
        RECT 1056.350 0.155 1064.250 4.280 ;
        RECT 1065.090 0.155 1072.990 4.280 ;
        RECT 1073.830 0.155 1081.730 4.280 ;
        RECT 1082.570 0.155 1090.470 4.280 ;
        RECT 1091.310 0.155 1099.210 4.280 ;
        RECT 1100.050 0.155 1107.950 4.280 ;
        RECT 1108.790 0.155 1116.690 4.280 ;
        RECT 1117.530 0.155 1125.430 4.280 ;
        RECT 1126.270 0.155 1134.170 4.280 ;
        RECT 1135.010 0.155 1142.910 4.280 ;
        RECT 1143.750 0.155 1151.650 4.280 ;
        RECT 1152.490 0.155 1160.390 4.280 ;
        RECT 1161.230 0.155 1169.130 4.280 ;
        RECT 1169.970 0.155 1177.870 4.280 ;
        RECT 1178.710 0.155 1186.610 4.280 ;
        RECT 1187.450 0.155 1195.350 4.280 ;
        RECT 1196.190 0.155 1204.090 4.280 ;
        RECT 1204.930 0.155 1212.830 4.280 ;
        RECT 1213.670 0.155 1221.570 4.280 ;
        RECT 1222.410 0.155 1230.310 4.280 ;
        RECT 1231.150 0.155 1239.050 4.280 ;
        RECT 1239.890 0.155 1247.790 4.280 ;
        RECT 1248.630 0.155 1256.530 4.280 ;
        RECT 1257.370 0.155 1265.270 4.280 ;
        RECT 1266.110 0.155 1274.010 4.280 ;
        RECT 1274.850 0.155 1282.750 4.280 ;
        RECT 1283.590 0.155 1291.490 4.280 ;
        RECT 1292.330 0.155 1300.230 4.280 ;
        RECT 1301.070 0.155 1308.970 4.280 ;
        RECT 1309.810 0.155 1317.710 4.280 ;
        RECT 1318.550 0.155 1326.450 4.280 ;
        RECT 1327.290 0.155 1335.190 4.280 ;
        RECT 1336.030 0.155 1343.930 4.280 ;
        RECT 1344.770 0.155 1352.670 4.280 ;
        RECT 1353.510 0.155 1361.410 4.280 ;
        RECT 1362.250 0.155 1370.150 4.280 ;
        RECT 1370.990 0.155 1378.890 4.280 ;
        RECT 1379.730 0.155 1387.630 4.280 ;
        RECT 1388.470 0.155 1396.370 4.280 ;
        RECT 1397.210 0.155 1405.110 4.280 ;
        RECT 1405.950 0.155 1413.850 4.280 ;
        RECT 1414.690 0.155 1422.590 4.280 ;
        RECT 1423.430 0.155 1431.330 4.280 ;
        RECT 1432.170 0.155 1440.070 4.280 ;
        RECT 1440.910 0.155 1448.810 4.280 ;
        RECT 1449.650 0.155 1457.550 4.280 ;
        RECT 1458.390 0.155 1466.290 4.280 ;
        RECT 1467.130 0.155 1475.030 4.280 ;
        RECT 1475.870 0.155 1483.770 4.280 ;
        RECT 1484.610 0.155 1492.510 4.280 ;
        RECT 1493.350 0.155 1501.250 4.280 ;
        RECT 1502.090 0.155 1509.990 4.280 ;
        RECT 1510.830 0.155 1518.730 4.280 ;
        RECT 1519.570 0.155 1527.470 4.280 ;
        RECT 1528.310 0.155 1536.210 4.280 ;
        RECT 1537.050 0.155 1544.950 4.280 ;
        RECT 1545.790 0.155 1553.690 4.280 ;
        RECT 1554.530 0.155 1562.430 4.280 ;
        RECT 1563.270 0.155 1571.170 4.280 ;
        RECT 1572.010 0.155 1579.910 4.280 ;
        RECT 1580.750 0.155 1588.650 4.280 ;
        RECT 1589.490 0.155 1597.390 4.280 ;
        RECT 1598.230 0.155 1606.130 4.280 ;
        RECT 1606.970 0.155 1614.870 4.280 ;
        RECT 1615.710 0.155 1623.610 4.280 ;
        RECT 1624.450 0.155 1632.350 4.280 ;
        RECT 1633.190 0.155 1641.090 4.280 ;
        RECT 1641.930 0.155 1649.830 4.280 ;
        RECT 1650.670 0.155 1658.570 4.280 ;
        RECT 1659.410 0.155 1667.310 4.280 ;
        RECT 1668.150 0.155 1676.050 4.280 ;
        RECT 1676.890 0.155 1684.790 4.280 ;
        RECT 1685.630 0.155 1693.530 4.280 ;
        RECT 1694.370 0.155 1702.270 4.280 ;
        RECT 1703.110 0.155 1711.010 4.280 ;
        RECT 1711.850 0.155 1719.750 4.280 ;
        RECT 1720.590 0.155 1728.490 4.280 ;
        RECT 1729.330 0.155 1737.230 4.280 ;
        RECT 1738.070 0.155 1745.970 4.280 ;
        RECT 1746.810 0.155 1754.710 4.280 ;
        RECT 1755.550 0.155 1763.450 4.280 ;
        RECT 1764.290 0.155 1772.190 4.280 ;
        RECT 1773.030 0.155 1780.930 4.280 ;
        RECT 1781.770 0.155 1789.670 4.280 ;
        RECT 1790.510 0.155 1798.410 4.280 ;
        RECT 1799.250 0.155 1807.150 4.280 ;
        RECT 1807.990 0.155 1815.890 4.280 ;
        RECT 1816.730 0.155 1824.630 4.280 ;
        RECT 1825.470 0.155 1833.370 4.280 ;
        RECT 1834.210 0.155 1842.110 4.280 ;
        RECT 1842.950 0.155 1850.850 4.280 ;
        RECT 1851.690 0.155 1859.590 4.280 ;
        RECT 1860.430 0.155 1868.330 4.280 ;
        RECT 1869.170 0.155 1877.070 4.280 ;
        RECT 1877.910 0.155 1885.810 4.280 ;
        RECT 1886.650 0.155 1894.550 4.280 ;
        RECT 1895.390 0.155 1903.290 4.280 ;
        RECT 1904.130 0.155 1912.030 4.280 ;
        RECT 1912.870 0.155 1920.770 4.280 ;
        RECT 1921.610 0.155 1929.510 4.280 ;
        RECT 1930.350 0.155 1938.250 4.280 ;
        RECT 1939.090 0.155 1946.990 4.280 ;
        RECT 1947.830 0.155 1955.730 4.280 ;
        RECT 1956.570 0.155 1964.470 4.280 ;
        RECT 1965.310 0.155 1973.210 4.280 ;
        RECT 1974.050 0.155 1981.950 4.280 ;
        RECT 1982.790 0.155 1990.690 4.280 ;
        RECT 1991.530 0.155 1999.430 4.280 ;
        RECT 2000.270 0.155 2008.170 4.280 ;
        RECT 2009.010 0.155 2016.910 4.280 ;
        RECT 2017.750 0.155 2025.650 4.280 ;
        RECT 2026.490 0.155 2034.390 4.280 ;
        RECT 2035.230 0.155 2043.130 4.280 ;
        RECT 2043.970 0.155 2051.870 4.280 ;
        RECT 2052.710 0.155 2060.610 4.280 ;
        RECT 2061.450 0.155 2069.350 4.280 ;
        RECT 2070.190 0.155 2078.090 4.280 ;
        RECT 2078.930 0.155 2086.830 4.280 ;
        RECT 2087.670 0.155 2095.570 4.280 ;
        RECT 2096.410 0.155 2104.310 4.280 ;
        RECT 2105.150 0.155 2113.050 4.280 ;
        RECT 2113.890 0.155 2121.790 4.280 ;
        RECT 2122.630 0.155 2130.530 4.280 ;
        RECT 2131.370 0.155 2139.270 4.280 ;
        RECT 2140.110 0.155 2148.010 4.280 ;
        RECT 2148.850 0.155 2156.750 4.280 ;
        RECT 2157.590 0.155 2196.860 4.280 ;
      LAYER met3 ;
        RECT 4.000 755.840 2196.000 846.425 ;
        RECT 4.000 754.440 2195.600 755.840 ;
        RECT 4.000 753.120 2196.000 754.440 ;
        RECT 4.000 751.720 2195.600 753.120 ;
        RECT 4.000 750.400 2196.000 751.720 ;
        RECT 4.400 749.000 2195.600 750.400 ;
        RECT 4.000 747.680 2196.000 749.000 ;
        RECT 4.400 746.280 2195.600 747.680 ;
        RECT 4.000 744.960 2196.000 746.280 ;
        RECT 4.400 743.560 2195.600 744.960 ;
        RECT 4.000 742.240 2196.000 743.560 ;
        RECT 4.400 740.840 2195.600 742.240 ;
        RECT 4.000 739.520 2196.000 740.840 ;
        RECT 4.400 738.120 2195.600 739.520 ;
        RECT 4.000 736.800 2196.000 738.120 ;
        RECT 4.400 735.400 2195.600 736.800 ;
        RECT 4.000 734.080 2196.000 735.400 ;
        RECT 4.400 732.680 2195.600 734.080 ;
        RECT 4.000 731.360 2196.000 732.680 ;
        RECT 4.400 729.960 2195.600 731.360 ;
        RECT 4.000 728.640 2196.000 729.960 ;
        RECT 4.400 727.240 2195.600 728.640 ;
        RECT 4.000 725.920 2196.000 727.240 ;
        RECT 4.400 724.520 2195.600 725.920 ;
        RECT 4.000 723.200 2196.000 724.520 ;
        RECT 4.400 721.800 2195.600 723.200 ;
        RECT 4.000 720.480 2196.000 721.800 ;
        RECT 4.400 719.080 2195.600 720.480 ;
        RECT 4.000 717.760 2196.000 719.080 ;
        RECT 4.400 716.360 2195.600 717.760 ;
        RECT 4.000 715.040 2196.000 716.360 ;
        RECT 4.400 713.640 2195.600 715.040 ;
        RECT 4.000 712.320 2196.000 713.640 ;
        RECT 4.400 710.920 2195.600 712.320 ;
        RECT 4.000 709.600 2196.000 710.920 ;
        RECT 4.400 708.200 2195.600 709.600 ;
        RECT 4.000 706.880 2196.000 708.200 ;
        RECT 4.400 705.480 2195.600 706.880 ;
        RECT 4.000 704.160 2196.000 705.480 ;
        RECT 4.400 702.760 2195.600 704.160 ;
        RECT 4.000 701.440 2196.000 702.760 ;
        RECT 4.400 700.040 2195.600 701.440 ;
        RECT 4.000 698.720 2196.000 700.040 ;
        RECT 4.400 697.320 2195.600 698.720 ;
        RECT 4.000 696.000 2196.000 697.320 ;
        RECT 4.400 694.600 2195.600 696.000 ;
        RECT 4.000 693.280 2196.000 694.600 ;
        RECT 4.400 691.880 2195.600 693.280 ;
        RECT 4.000 690.560 2196.000 691.880 ;
        RECT 4.400 689.160 2195.600 690.560 ;
        RECT 4.000 687.840 2196.000 689.160 ;
        RECT 4.400 686.440 2195.600 687.840 ;
        RECT 4.000 685.120 2196.000 686.440 ;
        RECT 4.400 683.720 2195.600 685.120 ;
        RECT 4.000 682.400 2196.000 683.720 ;
        RECT 4.400 681.000 2195.600 682.400 ;
        RECT 4.000 679.680 2196.000 681.000 ;
        RECT 4.400 678.280 2195.600 679.680 ;
        RECT 4.000 676.960 2196.000 678.280 ;
        RECT 4.400 675.560 2195.600 676.960 ;
        RECT 4.000 674.240 2196.000 675.560 ;
        RECT 4.400 672.840 2195.600 674.240 ;
        RECT 4.000 671.520 2196.000 672.840 ;
        RECT 4.400 670.120 2195.600 671.520 ;
        RECT 4.000 668.800 2196.000 670.120 ;
        RECT 4.400 667.400 2195.600 668.800 ;
        RECT 4.000 666.080 2196.000 667.400 ;
        RECT 4.400 664.680 2195.600 666.080 ;
        RECT 4.000 663.360 2196.000 664.680 ;
        RECT 4.400 661.960 2195.600 663.360 ;
        RECT 4.000 660.640 2196.000 661.960 ;
        RECT 4.400 659.240 2195.600 660.640 ;
        RECT 4.000 657.920 2196.000 659.240 ;
        RECT 4.400 656.520 2195.600 657.920 ;
        RECT 4.000 655.200 2196.000 656.520 ;
        RECT 4.400 653.800 2195.600 655.200 ;
        RECT 4.000 652.480 2196.000 653.800 ;
        RECT 4.400 651.080 2195.600 652.480 ;
        RECT 4.000 649.760 2196.000 651.080 ;
        RECT 4.400 648.360 2195.600 649.760 ;
        RECT 4.000 647.040 2196.000 648.360 ;
        RECT 4.400 645.640 2195.600 647.040 ;
        RECT 4.000 644.320 2196.000 645.640 ;
        RECT 4.400 642.920 2195.600 644.320 ;
        RECT 4.000 641.600 2196.000 642.920 ;
        RECT 4.400 640.200 2195.600 641.600 ;
        RECT 4.000 638.880 2196.000 640.200 ;
        RECT 4.400 637.480 2195.600 638.880 ;
        RECT 4.000 636.160 2196.000 637.480 ;
        RECT 4.400 634.760 2195.600 636.160 ;
        RECT 4.000 633.440 2196.000 634.760 ;
        RECT 4.400 632.040 2195.600 633.440 ;
        RECT 4.000 630.720 2196.000 632.040 ;
        RECT 4.400 629.320 2195.600 630.720 ;
        RECT 4.000 628.000 2196.000 629.320 ;
        RECT 4.400 626.600 2195.600 628.000 ;
        RECT 4.000 625.280 2196.000 626.600 ;
        RECT 4.400 623.880 2195.600 625.280 ;
        RECT 4.000 622.560 2196.000 623.880 ;
        RECT 4.400 621.160 2195.600 622.560 ;
        RECT 4.000 619.840 2196.000 621.160 ;
        RECT 4.400 618.440 2195.600 619.840 ;
        RECT 4.000 617.120 2196.000 618.440 ;
        RECT 4.400 615.720 2195.600 617.120 ;
        RECT 4.000 614.400 2196.000 615.720 ;
        RECT 4.400 613.000 2195.600 614.400 ;
        RECT 4.000 611.680 2196.000 613.000 ;
        RECT 4.400 610.280 2195.600 611.680 ;
        RECT 4.000 608.960 2196.000 610.280 ;
        RECT 4.400 607.560 2195.600 608.960 ;
        RECT 4.000 606.240 2196.000 607.560 ;
        RECT 4.400 604.840 2195.600 606.240 ;
        RECT 4.000 603.520 2196.000 604.840 ;
        RECT 4.400 602.120 2195.600 603.520 ;
        RECT 4.000 600.800 2196.000 602.120 ;
        RECT 4.400 599.400 2195.600 600.800 ;
        RECT 4.000 598.080 2196.000 599.400 ;
        RECT 4.400 596.680 2195.600 598.080 ;
        RECT 4.000 595.360 2196.000 596.680 ;
        RECT 4.400 593.960 2195.600 595.360 ;
        RECT 4.000 592.640 2196.000 593.960 ;
        RECT 4.400 591.240 2195.600 592.640 ;
        RECT 4.000 589.920 2196.000 591.240 ;
        RECT 4.400 588.520 2195.600 589.920 ;
        RECT 4.000 587.200 2196.000 588.520 ;
        RECT 4.400 585.800 2195.600 587.200 ;
        RECT 4.000 584.480 2196.000 585.800 ;
        RECT 4.400 583.080 2195.600 584.480 ;
        RECT 4.000 581.760 2196.000 583.080 ;
        RECT 4.400 580.360 2195.600 581.760 ;
        RECT 4.000 579.040 2196.000 580.360 ;
        RECT 4.400 577.640 2195.600 579.040 ;
        RECT 4.000 576.320 2196.000 577.640 ;
        RECT 4.400 574.920 2195.600 576.320 ;
        RECT 4.000 573.600 2196.000 574.920 ;
        RECT 4.400 572.200 2195.600 573.600 ;
        RECT 4.000 570.880 2196.000 572.200 ;
        RECT 4.400 569.480 2195.600 570.880 ;
        RECT 4.000 568.160 2196.000 569.480 ;
        RECT 4.400 566.760 2195.600 568.160 ;
        RECT 4.000 565.440 2196.000 566.760 ;
        RECT 4.400 564.040 2195.600 565.440 ;
        RECT 4.000 562.720 2196.000 564.040 ;
        RECT 4.400 561.320 2195.600 562.720 ;
        RECT 4.000 560.000 2196.000 561.320 ;
        RECT 4.400 558.600 2195.600 560.000 ;
        RECT 4.000 557.280 2196.000 558.600 ;
        RECT 4.400 555.880 2195.600 557.280 ;
        RECT 4.000 554.560 2196.000 555.880 ;
        RECT 4.400 553.160 2195.600 554.560 ;
        RECT 4.000 551.840 2196.000 553.160 ;
        RECT 4.400 550.440 2195.600 551.840 ;
        RECT 4.000 549.120 2196.000 550.440 ;
        RECT 4.400 547.720 2195.600 549.120 ;
        RECT 4.000 546.400 2196.000 547.720 ;
        RECT 4.400 545.000 2195.600 546.400 ;
        RECT 4.000 543.680 2196.000 545.000 ;
        RECT 4.400 542.280 2195.600 543.680 ;
        RECT 4.000 540.960 2196.000 542.280 ;
        RECT 4.400 539.560 2195.600 540.960 ;
        RECT 4.000 538.240 2196.000 539.560 ;
        RECT 4.400 536.840 2195.600 538.240 ;
        RECT 4.000 535.520 2196.000 536.840 ;
        RECT 4.400 534.120 2195.600 535.520 ;
        RECT 4.000 532.800 2196.000 534.120 ;
        RECT 4.400 531.400 2195.600 532.800 ;
        RECT 4.000 530.080 2196.000 531.400 ;
        RECT 4.400 528.680 2195.600 530.080 ;
        RECT 4.000 527.360 2196.000 528.680 ;
        RECT 4.400 525.960 2195.600 527.360 ;
        RECT 4.000 524.640 2196.000 525.960 ;
        RECT 4.400 523.240 2195.600 524.640 ;
        RECT 4.000 521.920 2196.000 523.240 ;
        RECT 4.400 520.520 2195.600 521.920 ;
        RECT 4.000 519.200 2196.000 520.520 ;
        RECT 4.400 517.800 2195.600 519.200 ;
        RECT 4.000 516.480 2196.000 517.800 ;
        RECT 4.400 515.080 2195.600 516.480 ;
        RECT 4.000 513.760 2196.000 515.080 ;
        RECT 4.400 512.360 2195.600 513.760 ;
        RECT 4.000 511.040 2196.000 512.360 ;
        RECT 4.400 509.640 2195.600 511.040 ;
        RECT 4.000 508.320 2196.000 509.640 ;
        RECT 4.400 506.920 2195.600 508.320 ;
        RECT 4.000 505.600 2196.000 506.920 ;
        RECT 4.400 504.200 2195.600 505.600 ;
        RECT 4.000 502.880 2196.000 504.200 ;
        RECT 4.400 501.480 2195.600 502.880 ;
        RECT 4.000 500.160 2196.000 501.480 ;
        RECT 4.400 498.760 2195.600 500.160 ;
        RECT 4.000 497.440 2196.000 498.760 ;
        RECT 4.400 496.040 2195.600 497.440 ;
        RECT 4.000 494.720 2196.000 496.040 ;
        RECT 4.400 493.320 2195.600 494.720 ;
        RECT 4.000 492.000 2196.000 493.320 ;
        RECT 4.400 490.600 2195.600 492.000 ;
        RECT 4.000 489.280 2196.000 490.600 ;
        RECT 4.400 487.880 2195.600 489.280 ;
        RECT 4.000 486.560 2196.000 487.880 ;
        RECT 4.400 485.160 2195.600 486.560 ;
        RECT 4.000 483.840 2196.000 485.160 ;
        RECT 4.400 482.440 2195.600 483.840 ;
        RECT 4.000 481.120 2196.000 482.440 ;
        RECT 4.400 479.720 2195.600 481.120 ;
        RECT 4.000 478.400 2196.000 479.720 ;
        RECT 4.400 477.000 2195.600 478.400 ;
        RECT 4.000 475.680 2196.000 477.000 ;
        RECT 4.400 474.280 2195.600 475.680 ;
        RECT 4.000 472.960 2196.000 474.280 ;
        RECT 4.400 471.560 2195.600 472.960 ;
        RECT 4.000 470.240 2196.000 471.560 ;
        RECT 4.400 468.840 2195.600 470.240 ;
        RECT 4.000 467.520 2196.000 468.840 ;
        RECT 4.400 466.120 2195.600 467.520 ;
        RECT 4.000 464.800 2196.000 466.120 ;
        RECT 4.400 463.400 2195.600 464.800 ;
        RECT 4.000 462.080 2196.000 463.400 ;
        RECT 4.400 460.680 2195.600 462.080 ;
        RECT 4.000 459.360 2196.000 460.680 ;
        RECT 4.400 457.960 2195.600 459.360 ;
        RECT 4.000 456.640 2196.000 457.960 ;
        RECT 4.400 455.240 2195.600 456.640 ;
        RECT 4.000 453.920 2196.000 455.240 ;
        RECT 4.400 452.520 2195.600 453.920 ;
        RECT 4.000 451.200 2196.000 452.520 ;
        RECT 4.400 449.800 2195.600 451.200 ;
        RECT 4.000 448.480 2196.000 449.800 ;
        RECT 4.400 447.080 2195.600 448.480 ;
        RECT 4.000 445.760 2196.000 447.080 ;
        RECT 4.400 444.360 2195.600 445.760 ;
        RECT 4.000 443.040 2196.000 444.360 ;
        RECT 4.400 441.640 2195.600 443.040 ;
        RECT 4.000 440.320 2196.000 441.640 ;
        RECT 4.400 438.920 2195.600 440.320 ;
        RECT 4.000 437.600 2196.000 438.920 ;
        RECT 4.400 436.200 2195.600 437.600 ;
        RECT 4.000 434.880 2196.000 436.200 ;
        RECT 4.400 433.480 2195.600 434.880 ;
        RECT 4.000 432.160 2196.000 433.480 ;
        RECT 4.400 430.760 2195.600 432.160 ;
        RECT 4.000 429.440 2196.000 430.760 ;
        RECT 4.400 428.040 2195.600 429.440 ;
        RECT 4.000 426.720 2196.000 428.040 ;
        RECT 4.400 425.320 2195.600 426.720 ;
        RECT 4.000 424.000 2196.000 425.320 ;
        RECT 4.400 422.600 2195.600 424.000 ;
        RECT 4.000 421.280 2196.000 422.600 ;
        RECT 4.400 419.880 2195.600 421.280 ;
        RECT 4.000 418.560 2196.000 419.880 ;
        RECT 4.400 417.160 2195.600 418.560 ;
        RECT 4.000 415.840 2196.000 417.160 ;
        RECT 4.400 414.440 2195.600 415.840 ;
        RECT 4.000 413.120 2196.000 414.440 ;
        RECT 4.400 411.720 2195.600 413.120 ;
        RECT 4.000 410.400 2196.000 411.720 ;
        RECT 4.400 409.000 2195.600 410.400 ;
        RECT 4.000 407.680 2196.000 409.000 ;
        RECT 4.400 406.280 2195.600 407.680 ;
        RECT 4.000 404.960 2196.000 406.280 ;
        RECT 4.400 403.560 2195.600 404.960 ;
        RECT 4.000 402.240 2196.000 403.560 ;
        RECT 4.400 400.840 2195.600 402.240 ;
        RECT 4.000 399.520 2196.000 400.840 ;
        RECT 4.400 398.120 2195.600 399.520 ;
        RECT 4.000 396.800 2196.000 398.120 ;
        RECT 4.400 395.400 2195.600 396.800 ;
        RECT 4.000 394.080 2196.000 395.400 ;
        RECT 4.400 392.680 2195.600 394.080 ;
        RECT 4.000 391.360 2196.000 392.680 ;
        RECT 4.400 389.960 2195.600 391.360 ;
        RECT 4.000 388.640 2196.000 389.960 ;
        RECT 4.400 387.240 2195.600 388.640 ;
        RECT 4.000 385.920 2196.000 387.240 ;
        RECT 4.400 384.520 2195.600 385.920 ;
        RECT 4.000 383.200 2196.000 384.520 ;
        RECT 4.400 381.800 2195.600 383.200 ;
        RECT 4.000 380.480 2196.000 381.800 ;
        RECT 4.400 379.080 2195.600 380.480 ;
        RECT 4.000 377.760 2196.000 379.080 ;
        RECT 4.400 376.360 2195.600 377.760 ;
        RECT 4.000 375.040 2196.000 376.360 ;
        RECT 4.400 373.640 2195.600 375.040 ;
        RECT 4.000 372.320 2196.000 373.640 ;
        RECT 4.400 370.920 2195.600 372.320 ;
        RECT 4.000 369.600 2196.000 370.920 ;
        RECT 4.400 368.200 2195.600 369.600 ;
        RECT 4.000 366.880 2196.000 368.200 ;
        RECT 4.400 365.480 2195.600 366.880 ;
        RECT 4.000 364.160 2196.000 365.480 ;
        RECT 4.400 362.760 2195.600 364.160 ;
        RECT 4.000 361.440 2196.000 362.760 ;
        RECT 4.400 360.040 2195.600 361.440 ;
        RECT 4.000 358.720 2196.000 360.040 ;
        RECT 4.400 357.320 2195.600 358.720 ;
        RECT 4.000 356.000 2196.000 357.320 ;
        RECT 4.400 354.600 2195.600 356.000 ;
        RECT 4.000 353.280 2196.000 354.600 ;
        RECT 4.400 351.880 2195.600 353.280 ;
        RECT 4.000 350.560 2196.000 351.880 ;
        RECT 4.400 349.160 2195.600 350.560 ;
        RECT 4.000 347.840 2196.000 349.160 ;
        RECT 4.400 346.440 2195.600 347.840 ;
        RECT 4.000 345.120 2196.000 346.440 ;
        RECT 4.400 343.720 2195.600 345.120 ;
        RECT 4.000 342.400 2196.000 343.720 ;
        RECT 4.400 341.000 2195.600 342.400 ;
        RECT 4.000 339.680 2196.000 341.000 ;
        RECT 4.400 338.280 2195.600 339.680 ;
        RECT 4.000 336.960 2196.000 338.280 ;
        RECT 4.400 335.560 2195.600 336.960 ;
        RECT 4.000 334.240 2196.000 335.560 ;
        RECT 4.400 332.840 2195.600 334.240 ;
        RECT 4.000 331.520 2196.000 332.840 ;
        RECT 4.400 330.120 2195.600 331.520 ;
        RECT 4.000 328.800 2196.000 330.120 ;
        RECT 4.400 327.400 2195.600 328.800 ;
        RECT 4.000 326.080 2196.000 327.400 ;
        RECT 4.400 324.680 2195.600 326.080 ;
        RECT 4.000 323.360 2196.000 324.680 ;
        RECT 4.400 321.960 2195.600 323.360 ;
        RECT 4.000 320.640 2196.000 321.960 ;
        RECT 4.400 319.240 2195.600 320.640 ;
        RECT 4.000 317.920 2196.000 319.240 ;
        RECT 4.400 316.520 2195.600 317.920 ;
        RECT 4.000 315.200 2196.000 316.520 ;
        RECT 4.400 313.800 2195.600 315.200 ;
        RECT 4.000 312.480 2196.000 313.800 ;
        RECT 4.400 311.080 2195.600 312.480 ;
        RECT 4.000 309.760 2196.000 311.080 ;
        RECT 4.400 308.360 2195.600 309.760 ;
        RECT 4.000 307.040 2196.000 308.360 ;
        RECT 4.400 305.640 2195.600 307.040 ;
        RECT 4.000 304.320 2196.000 305.640 ;
        RECT 4.400 302.920 2195.600 304.320 ;
        RECT 4.000 301.600 2196.000 302.920 ;
        RECT 4.400 300.200 2195.600 301.600 ;
        RECT 4.000 298.880 2196.000 300.200 ;
        RECT 4.400 297.480 2195.600 298.880 ;
        RECT 4.000 296.160 2196.000 297.480 ;
        RECT 4.400 294.760 2195.600 296.160 ;
        RECT 4.000 293.440 2196.000 294.760 ;
        RECT 4.400 292.040 2195.600 293.440 ;
        RECT 4.000 290.720 2196.000 292.040 ;
        RECT 4.400 289.320 2195.600 290.720 ;
        RECT 4.000 288.000 2196.000 289.320 ;
        RECT 4.400 286.600 2195.600 288.000 ;
        RECT 4.000 285.280 2196.000 286.600 ;
        RECT 4.400 283.880 2195.600 285.280 ;
        RECT 4.000 282.560 2196.000 283.880 ;
        RECT 4.400 281.160 2195.600 282.560 ;
        RECT 4.000 279.840 2196.000 281.160 ;
        RECT 4.400 278.440 2195.600 279.840 ;
        RECT 4.000 277.120 2196.000 278.440 ;
        RECT 4.400 275.720 2195.600 277.120 ;
        RECT 4.000 274.400 2196.000 275.720 ;
        RECT 4.400 273.000 2195.600 274.400 ;
        RECT 4.000 271.680 2196.000 273.000 ;
        RECT 4.400 270.280 2195.600 271.680 ;
        RECT 4.000 268.960 2196.000 270.280 ;
        RECT 4.400 267.560 2195.600 268.960 ;
        RECT 4.000 266.240 2196.000 267.560 ;
        RECT 4.400 264.840 2195.600 266.240 ;
        RECT 4.000 263.520 2196.000 264.840 ;
        RECT 4.400 262.120 2195.600 263.520 ;
        RECT 4.000 260.800 2196.000 262.120 ;
        RECT 4.400 259.400 2195.600 260.800 ;
        RECT 4.000 258.080 2196.000 259.400 ;
        RECT 4.400 256.680 2195.600 258.080 ;
        RECT 4.000 255.360 2196.000 256.680 ;
        RECT 4.400 253.960 2195.600 255.360 ;
        RECT 4.000 252.640 2196.000 253.960 ;
        RECT 4.400 251.240 2195.600 252.640 ;
        RECT 4.000 249.920 2196.000 251.240 ;
        RECT 4.400 248.520 2195.600 249.920 ;
        RECT 4.000 247.200 2196.000 248.520 ;
        RECT 4.400 245.800 2195.600 247.200 ;
        RECT 4.000 244.480 2196.000 245.800 ;
        RECT 4.400 243.080 2195.600 244.480 ;
        RECT 4.000 241.760 2196.000 243.080 ;
        RECT 4.400 240.360 2195.600 241.760 ;
        RECT 4.000 239.040 2196.000 240.360 ;
        RECT 4.400 237.640 2195.600 239.040 ;
        RECT 4.000 236.320 2196.000 237.640 ;
        RECT 4.400 234.920 2195.600 236.320 ;
        RECT 4.000 233.600 2196.000 234.920 ;
        RECT 4.400 232.200 2195.600 233.600 ;
        RECT 4.000 230.880 2196.000 232.200 ;
        RECT 4.400 229.480 2195.600 230.880 ;
        RECT 4.000 228.160 2196.000 229.480 ;
        RECT 4.400 226.760 2195.600 228.160 ;
        RECT 4.000 225.440 2196.000 226.760 ;
        RECT 4.400 224.040 2195.600 225.440 ;
        RECT 4.000 222.720 2196.000 224.040 ;
        RECT 4.400 221.320 2195.600 222.720 ;
        RECT 4.000 220.000 2196.000 221.320 ;
        RECT 4.400 218.600 2195.600 220.000 ;
        RECT 4.000 217.280 2196.000 218.600 ;
        RECT 4.400 215.880 2195.600 217.280 ;
        RECT 4.000 214.560 2196.000 215.880 ;
        RECT 4.400 213.160 2195.600 214.560 ;
        RECT 4.000 211.840 2196.000 213.160 ;
        RECT 4.400 210.440 2195.600 211.840 ;
        RECT 4.000 209.120 2196.000 210.440 ;
        RECT 4.400 207.720 2195.600 209.120 ;
        RECT 4.000 206.400 2196.000 207.720 ;
        RECT 4.400 205.000 2195.600 206.400 ;
        RECT 4.000 203.680 2196.000 205.000 ;
        RECT 4.400 202.280 2195.600 203.680 ;
        RECT 4.000 200.960 2196.000 202.280 ;
        RECT 4.400 199.560 2195.600 200.960 ;
        RECT 4.000 198.240 2196.000 199.560 ;
        RECT 4.400 196.840 2195.600 198.240 ;
        RECT 4.000 195.520 2196.000 196.840 ;
        RECT 4.400 194.120 2195.600 195.520 ;
        RECT 4.000 192.800 2196.000 194.120 ;
        RECT 4.400 191.400 2195.600 192.800 ;
        RECT 4.000 190.080 2196.000 191.400 ;
        RECT 4.400 188.680 2195.600 190.080 ;
        RECT 4.000 187.360 2196.000 188.680 ;
        RECT 4.400 185.960 2195.600 187.360 ;
        RECT 4.000 184.640 2196.000 185.960 ;
        RECT 4.400 183.240 2195.600 184.640 ;
        RECT 4.000 181.920 2196.000 183.240 ;
        RECT 4.400 180.520 2195.600 181.920 ;
        RECT 4.000 179.200 2196.000 180.520 ;
        RECT 4.400 177.800 2195.600 179.200 ;
        RECT 4.000 176.480 2196.000 177.800 ;
        RECT 4.400 175.080 2195.600 176.480 ;
        RECT 4.000 173.760 2196.000 175.080 ;
        RECT 4.400 172.360 2195.600 173.760 ;
        RECT 4.000 171.040 2196.000 172.360 ;
        RECT 4.400 169.640 2195.600 171.040 ;
        RECT 4.000 168.320 2196.000 169.640 ;
        RECT 4.400 166.920 2195.600 168.320 ;
        RECT 4.000 165.600 2196.000 166.920 ;
        RECT 4.400 164.200 2195.600 165.600 ;
        RECT 4.000 162.880 2196.000 164.200 ;
        RECT 4.400 161.480 2195.600 162.880 ;
        RECT 4.000 160.160 2196.000 161.480 ;
        RECT 4.400 158.760 2195.600 160.160 ;
        RECT 4.000 157.440 2196.000 158.760 ;
        RECT 4.400 156.040 2195.600 157.440 ;
        RECT 4.000 154.720 2196.000 156.040 ;
        RECT 4.400 153.320 2195.600 154.720 ;
        RECT 4.000 152.000 2196.000 153.320 ;
        RECT 4.400 150.600 2195.600 152.000 ;
        RECT 4.000 149.280 2196.000 150.600 ;
        RECT 4.400 147.880 2195.600 149.280 ;
        RECT 4.000 146.560 2196.000 147.880 ;
        RECT 4.400 145.160 2195.600 146.560 ;
        RECT 4.000 143.840 2196.000 145.160 ;
        RECT 4.400 142.440 2195.600 143.840 ;
        RECT 4.000 141.120 2196.000 142.440 ;
        RECT 4.400 139.720 2195.600 141.120 ;
        RECT 4.000 138.400 2196.000 139.720 ;
        RECT 4.400 137.000 2195.600 138.400 ;
        RECT 4.000 135.680 2196.000 137.000 ;
        RECT 4.400 134.280 2195.600 135.680 ;
        RECT 4.000 132.960 2196.000 134.280 ;
        RECT 4.400 131.560 2195.600 132.960 ;
        RECT 4.000 130.240 2196.000 131.560 ;
        RECT 4.400 128.840 2195.600 130.240 ;
        RECT 4.000 127.520 2196.000 128.840 ;
        RECT 4.400 126.120 2195.600 127.520 ;
        RECT 4.000 124.800 2196.000 126.120 ;
        RECT 4.400 123.400 2195.600 124.800 ;
        RECT 4.000 122.080 2196.000 123.400 ;
        RECT 4.400 120.680 2195.600 122.080 ;
        RECT 4.000 119.360 2196.000 120.680 ;
        RECT 4.400 117.960 2195.600 119.360 ;
        RECT 4.000 116.640 2196.000 117.960 ;
        RECT 4.400 115.240 2195.600 116.640 ;
        RECT 4.000 113.920 2196.000 115.240 ;
        RECT 4.400 112.520 2195.600 113.920 ;
        RECT 4.000 111.200 2196.000 112.520 ;
        RECT 4.400 109.800 2195.600 111.200 ;
        RECT 4.000 108.480 2196.000 109.800 ;
        RECT 4.400 107.080 2195.600 108.480 ;
        RECT 4.000 105.760 2196.000 107.080 ;
        RECT 4.400 104.360 2195.600 105.760 ;
        RECT 4.000 103.040 2196.000 104.360 ;
        RECT 4.400 101.640 2195.600 103.040 ;
        RECT 4.000 100.320 2196.000 101.640 ;
        RECT 4.400 98.920 2195.600 100.320 ;
        RECT 4.000 97.600 2196.000 98.920 ;
        RECT 4.000 96.200 2195.600 97.600 ;
        RECT 4.000 94.880 2196.000 96.200 ;
        RECT 4.000 93.480 2195.600 94.880 ;
        RECT 4.000 0.175 2196.000 93.480 ;
      LAYER met4 ;
        RECT 16.855 838.400 2184.705 845.745 ;
        RECT 16.855 10.240 20.640 838.400 ;
        RECT 23.040 10.240 97.440 838.400 ;
        RECT 99.840 10.240 174.240 838.400 ;
        RECT 176.640 10.240 251.040 838.400 ;
        RECT 253.440 10.240 327.840 838.400 ;
        RECT 330.240 10.240 404.640 838.400 ;
        RECT 407.040 10.240 481.440 838.400 ;
        RECT 483.840 10.240 558.240 838.400 ;
        RECT 560.640 10.240 635.040 838.400 ;
        RECT 637.440 10.240 711.840 838.400 ;
        RECT 714.240 10.240 788.640 838.400 ;
        RECT 791.040 10.240 865.440 838.400 ;
        RECT 867.840 10.240 942.240 838.400 ;
        RECT 944.640 10.240 1019.040 838.400 ;
        RECT 1021.440 10.240 1095.840 838.400 ;
        RECT 1098.240 10.240 1172.640 838.400 ;
        RECT 1175.040 10.240 1249.440 838.400 ;
        RECT 1251.840 10.240 1326.240 838.400 ;
        RECT 1328.640 10.240 1403.040 838.400 ;
        RECT 1405.440 10.240 1479.840 838.400 ;
        RECT 1482.240 10.240 1556.640 838.400 ;
        RECT 1559.040 10.240 1633.440 838.400 ;
        RECT 1635.840 10.240 1710.240 838.400 ;
        RECT 1712.640 10.240 1787.040 838.400 ;
        RECT 1789.440 10.240 1863.840 838.400 ;
        RECT 1866.240 10.240 1940.640 838.400 ;
        RECT 1943.040 10.240 2017.440 838.400 ;
        RECT 2019.840 10.240 2094.240 838.400 ;
        RECT 2096.640 10.240 2171.040 838.400 ;
        RECT 2173.440 10.240 2184.705 838.400 ;
        RECT 16.855 0.175 2184.705 10.240 ;
  END
END vliw
END LIBRARY

