* NGSPICE file created from scrapcpu.ext - technology: sky130B

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_4 abstract view
.subckt sky130_fd_sc_hd__o2111a_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_4 abstract view
.subckt sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

.subckt scrapcpu io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15]
+ io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22] io_in[23]
+ io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30] io_in[31]
+ io_in[32] io_in[33] io_in[34] io_in[35] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14]
+ io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21]
+ io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29]
+ io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[3]
+ io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9] io_out[0] io_out[10]
+ io_out[11] io_out[12] io_out[13] io_out[14] io_out[15] io_out[16] io_out[17] io_out[18]
+ io_out[19] io_out[1] io_out[20] io_out[21] io_out[22] io_out[23] io_out[24] io_out[25]
+ io_out[26] io_out[27] io_out[28] io_out[29] io_out[2] io_out[30] io_out[31] io_out[32]
+ io_out[33] io_out[34] io_out[35] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ io_out[8] io_out[9] rst_n vccd1 vssd1 wb_clk_i
XTAP_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3155_ _2948_/A _2886_/A _3137_/C vssd1 vssd1 vccd1 vccd1 _3155_/X sky130_fd_sc_hd__a21o_1
X_3086_ _3086_/A _3086_/B vssd1 vssd1 vccd1 vccd1 _3691_/D sky130_fd_sc_hd__and2_1
X_2106_ _3193_/A0 hold401/X _2111_/S vssd1 vssd1 vccd1 vccd1 _2106_/X sky130_fd_sc_hd__mux2_1
X_2037_ _2854_/B _2035_/X _2036_/Y _1760_/A vssd1 vssd1 vccd1 vccd1 _2037_/X sky130_fd_sc_hd__o22a_1
XANTENNA__2651__A0 _2651_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2939_ _3103_/A _2939_/B vssd1 vssd1 vccd1 vccd1 _3623_/D sky130_fd_sc_hd__and2_1
XFILLER_0_17_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2403__A0 _2475_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold362 _2580_/X vssd1 vssd1 vccd1 vccd1 _3518_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold351 _3299_/Q vssd1 vssd1 vccd1 vccd1 hold351/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold340 _2235_/X vssd1 vssd1 vccd1 vccd1 _3266_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold395 _3535_/Q vssd1 vssd1 vccd1 vccd1 hold395/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold373 _3374_/Q vssd1 vssd1 vccd1 vccd1 hold373/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold384 _2652_/X vssd1 vssd1 vccd1 vccd1 _3580_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout75_A _2659_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1051 _2874_/X vssd1 vssd1 vccd1 vccd1 _2875_/B1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1040 _3313_/Q vssd1 vssd1 vccd1 vccd1 hold1040/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1073 _3600_/Q vssd1 vssd1 vccd1 vccd1 _2982_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1084 _3618_/Q vssd1 vssd1 vccd1 vccd1 _2966_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1062 _3346_/Q vssd1 vssd1 vccd1 vccd1 hold1062/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2084__B _2084_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2974__S _2987_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1684__A1 _2797_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2330__C1 _3108_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_48_wb_clk_i_A clkbuf_3_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_46_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3189__A1 _3203_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_84 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3773_ _3773_/A vssd1 vssd1 vccd1 vccd1 _3773_/X sky130_fd_sc_hd__buf_1
XFILLER_0_54_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2724_ _3626_/Q _2714_/B _2721_/Y _2710_/A vssd1 vssd1 vccd1 vccd1 _2724_/X sky130_fd_sc_hd__o211a_1
X_2655_ _2655_/A0 hold433/X _2660_/S vssd1 vssd1 vccd1 vccd1 _2655_/X sky130_fd_sc_hd__mux2_1
X_1606_ _3599_/Q vssd1 vssd1 vccd1 vccd1 _1606_/Y sky130_fd_sc_hd__inv_2
X_2586_ _2656_/A0 hold371/X _2590_/S vssd1 vssd1 vccd1 vccd1 _2586_/X sky130_fd_sc_hd__mux2_1
Xfanout127 _1849_/S1 vssd1 vssd1 vccd1 vccd1 _2219_/C sky130_fd_sc_hd__clkbuf_8
Xfanout116 hold1021/X vssd1 vssd1 vccd1 vccd1 _2195_/B sky130_fd_sc_hd__buf_8
Xfanout138 _1954_/S vssd1 vssd1 vccd1 vccd1 _2005_/S sky130_fd_sc_hd__clkbuf_8
Xfanout105 _1716_/X vssd1 vssd1 vccd1 vccd1 _2022_/A sky130_fd_sc_hd__clkbuf_8
Xfanout149 _2859_/A vssd1 vssd1 vccd1 vccd1 _1979_/A sky130_fd_sc_hd__buf_4
XFILLER_0_38_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3207_ _3636_/CLK _3207_/D vssd1 vssd1 vccd1 vccd1 _3207_/Q sky130_fd_sc_hd__dfxtp_1
X_3138_ hold957/X _3131_/X _3137_/X _3166_/C1 vssd1 vssd1 vccd1 vccd1 _3138_/X sky130_fd_sc_hd__o211a_1
X_3069_ _3019_/Y _3068_/Y _3062_/X vssd1 vssd1 vccd1 vccd1 _3069_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_49_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2624__A0 _2097_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold170 _2415_/X vssd1 vssd1 vccd1 vccd1 _3382_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold192 _2594_/X vssd1 vssd1 vccd1 vccd1 _3530_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold181 _3470_/Q vssd1 vssd1 vccd1 vccd1 hold181/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_28_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2091__A1 hold918/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2918__A1 _1712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2918__B2 _2940_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2440_ hold980/X _2650_/A0 _2443_/S vssd1 vssd1 vccd1 vccd1 _3402_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_51_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2371_ _3198_/A0 hold675/X _2371_/S vssd1 vssd1 vccd1 vccd1 _2371_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_75_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1902__A _2085_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_4_wb_clk_i_A clkbuf_leaf_5_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__2606__A0 _2655_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout125_A _1849_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2707_ _2762_/A _2707_/B _2707_/C vssd1 vssd1 vccd1 vccd1 _2779_/A sky130_fd_sc_hd__and3_1
Xscrapcpu_172 vssd1 vssd1 vccd1 vccd1 scrapcpu_172/HI io_out[29] sky130_fd_sc_hd__conb_1
X_3687_ _3692_/CLK _3687_/D vssd1 vssd1 vccd1 vccd1 _3687_/Q sky130_fd_sc_hd__dfxtp_1
Xscrapcpu_161 vssd1 vssd1 vccd1 vccd1 scrapcpu_161/HI io_oeb[7] sky130_fd_sc_hd__conb_1
X_2638_ _2097_/X hold599/X _2639_/S vssd1 vssd1 vccd1 vccd1 _2638_/X sky130_fd_sc_hd__mux2_1
X_2569_ _2660_/A0 hold701/X _2569_/S vssd1 vssd1 vccd1 vccd1 _2569_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_4_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1820__A1 _2076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1887__A1 _1889_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1982__S1 _1760_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output19_A _3769_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1940_ _1889_/A _1936_/Y _1938_/Y _1939_/Y vssd1 vssd1 vccd1 vccd1 _1940_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_28_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1871_ _2720_/B _2720_/C vssd1 vssd1 vccd1 vccd1 _2701_/B sky130_fd_sc_hd__and2_2
XFILLER_0_43_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3610_ _3646_/CLK _3610_/D vssd1 vssd1 vccd1 vccd1 _3610_/Q sky130_fd_sc_hd__dfxtp_1
X_3541_ _3543_/CLK _3541_/D vssd1 vssd1 vccd1 vccd1 _3541_/Q sky130_fd_sc_hd__dfxtp_1
Xhold917 _1682_/X vssd1 vssd1 vccd1 vccd1 _3243_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold906 _3620_/Q vssd1 vssd1 vccd1 vccd1 _2924_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_24_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold928 _3168_/X vssd1 vssd1 vccd1 vccd1 _3719_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3472_ _3744_/CLK _3472_/D vssd1 vssd1 vccd1 vccd1 _3472_/Q sky130_fd_sc_hd__dfxtp_1
Xhold939 _3002_/Y vssd1 vssd1 vccd1 vccd1 hold939/X sky130_fd_sc_hd__dlygate4sd3_1
X_2423_ hold317/X _2656_/A0 _2427_/S vssd1 vssd1 vccd1 vccd1 _2423_/X sky130_fd_sc_hd__mux2_1
X_2354_ hold985/X _2351_/Y _2353_/X _3058_/A vssd1 vssd1 vccd1 vccd1 _3328_/D sky130_fd_sc_hd__o211a_1
X_2285_ _2650_/A0 hold503/X _2288_/S vssd1 vssd1 vccd1 vccd1 _2285_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_79_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1807__A _2085_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3739_ _3739_/CLK _3739_/D vssd1 vssd1 vccd1 vccd1 _3739_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1869__A1 _1626_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2294__A1 _2651_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2070_ _2195_/B _2036_/Y _2069_/X _2854_/B vssd1 vssd1 vccd1 vccd1 _2070_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_72_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2982__S _2987_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2972_ hold447/X _3624_/Q _2999_/S vssd1 vssd1 vccd1 vccd1 _2972_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2037__A1 _2854_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2037__B2 _1760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1923_ _2682_/B _2682_/C vssd1 vssd1 vccd1 vccd1 _2687_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_73 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1854_ _2244_/A _1849_/X _2087_/A vssd1 vssd1 vccd1 vccd1 _1854_/Y sky130_fd_sc_hd__o21ai_1
Xhold703 _3553_/Q vssd1 vssd1 vccd1 vccd1 hold703/X sky130_fd_sc_hd__dlygate4sd3_1
X_1785_ _2185_/A _1785_/B vssd1 vssd1 vccd1 vccd1 _1785_/Y sky130_fd_sc_hd__nor2_1
Xhold736 _2382_/X vssd1 vssd1 vccd1 vccd1 _3354_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3524_ _3539_/CLK _3524_/D vssd1 vssd1 vccd1 vccd1 _3524_/Q sky130_fd_sc_hd__dfxtp_1
Xhold714 _2564_/X vssd1 vssd1 vccd1 vccd1 _3504_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold725 _3214_/Q vssd1 vssd1 vccd1 vccd1 hold725/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold758 _2590_/X vssd1 vssd1 vccd1 vccd1 _3527_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold769 _3524_/Q vssd1 vssd1 vccd1 vccd1 hold769/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold747 _3352_/Q vssd1 vssd1 vccd1 vccd1 hold747/X sky130_fd_sc_hd__dlygate4sd3_1
X_3455_ _3739_/CLK _3455_/D vssd1 vssd1 vccd1 vccd1 _3455_/Q sky130_fd_sc_hd__dfxtp_1
X_2406_ _3198_/A0 hold721/X _2406_/S vssd1 vssd1 vccd1 vccd1 _2406_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3170__C1 _3172_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3386_ _3654_/CLK _3386_/D vssd1 vssd1 vccd1 vccd1 _3386_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2458__A _2570_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2337_ _3198_/A0 hold743/X _2337_/S vssd1 vssd1 vccd1 vccd1 _2337_/X sky130_fd_sc_hd__mux2_1
X_2268_ _2268_/A _2278_/B vssd1 vssd1 vccd1 vccd1 _2268_/X sky130_fd_sc_hd__or2_1
X_2199_ _2643_/A1 hold461/X _2202_/S vssd1 vssd1 vccd1 vccd1 _2199_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2193__A _2195_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold30 hold30/A vssd1 vssd1 vccd1 vccd1 hold30/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 hold41/A vssd1 vssd1 vccd1 vccd1 hold41/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold63 hold63/A vssd1 vssd1 vccd1 vccd1 hold63/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold52 hold52/A vssd1 vssd1 vccd1 vccd1 hold52/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 hold74/A vssd1 vssd1 vccd1 vccd1 hold74/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 hold85/A vssd1 vssd1 vccd1 vccd1 hold85/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2267__A1 _3058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold96 hold96/A vssd1 vssd1 vccd1 vccd1 hold96/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_85_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_3_7__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_3_7__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__3199__A _3199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2019__A1 _2479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_14_wb_clk_i clkbuf_3_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3543_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_26_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2977__S _2987_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3240_ _3575_/CLK _3240_/D vssd1 vssd1 vccd1 vccd1 _3240_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3152__C1 _3103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3171_ _3171_/A _3181_/B vssd1 vssd1 vccd1 vccd1 _3171_/X sky130_fd_sc_hd__or2_1
XANTENNA__1702__B1 _2876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2122_ _3720_/Q _3719_/Q _2146_/A vssd1 vssd1 vccd1 vccd1 _2154_/B sky130_fd_sc_hd__and3_1
XANTENNA__2428__D _2480_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2258__A1 _2659_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2053_ _3183_/B _3096_/A vssd1 vssd1 vccd1 vccd1 _2169_/B sky130_fd_sc_hd__nand2_2
XANTENNA__1910__A _2014_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1769__B1 _2854_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2955_ _2955_/A _2955_/B vssd1 vssd1 vccd1 vccd1 _2959_/S sky130_fd_sc_hd__or2_2
XFILLER_0_29_297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2886_ _2886_/A vssd1 vssd1 vccd1 vccd1 _3137_/B sky130_fd_sc_hd__inv_2
X_1906_ _2244_/A _1902_/Y _1904_/X _1905_/Y vssd1 vssd1 vccd1 vccd1 _1906_/X sky130_fd_sc_hd__a31o_1
X_1837_ hold31/A hold17/A hold9/A _3424_/Q _2244_/B _2185_/C vssd1 vssd1 vccd1 vccd1
+ _1838_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_32_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold511 _3569_/Q vssd1 vssd1 vccd1 vccd1 hold511/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold500 _2233_/X vssd1 vssd1 vccd1 vccd1 _3264_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold522 _2532_/X vssd1 vssd1 vccd1 vccd1 _3477_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold533 _3537_/Q vssd1 vssd1 vccd1 vccd1 hold533/X sky130_fd_sc_hd__dlygate4sd3_1
X_3507_ _3543_/CLK _3507_/D vssd1 vssd1 vccd1 vccd1 _3507_/Q sky130_fd_sc_hd__dfxtp_1
Xhold544 _2240_/X vssd1 vssd1 vccd1 vccd1 _3270_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1768_ _1713_/X _2868_/C _2731_/A2 hold767/X vssd1 vssd1 vccd1 vccd1 _1768_/X sky130_fd_sc_hd__o22a_1
Xhold588 _2469_/X vssd1 vssd1 vccd1 vccd1 _3427_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold555 _3254_/Q vssd1 vssd1 vccd1 vccd1 hold555/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold577 _3302_/Q vssd1 vssd1 vccd1 vccd1 hold577/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1699_ hold836/X _1698_/X _2961_/A vssd1 vssd1 vccd1 vccd1 _1699_/Y sky130_fd_sc_hd__a21oi_1
Xhold566 _2980_/X vssd1 vssd1 vccd1 vccd1 _3655_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold599 _3568_/Q vssd1 vssd1 vccd1 vccd1 hold599/X sky130_fd_sc_hd__dlygate4sd3_1
X_3438_ _3743_/CLK hold70/X vssd1 vssd1 vccd1 vccd1 hold69/A sky130_fd_sc_hd__dfxtp_1
X_3369_ _3543_/CLK _3369_/D vssd1 vssd1 vccd1 vccd1 _3369_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2249__A1 _2650_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput20 _3770_/X vssd1 vssd1 vccd1 vccd1 io_oeb[11] sky130_fd_sc_hd__buf_12
Xoutput31 _3622_/Q vssd1 vssd1 vccd1 vccd1 io_oeb[32] sky130_fd_sc_hd__buf_12
Xoutput42 _3402_/Q vssd1 vssd1 vccd1 vccd1 io_out[11] sky130_fd_sc_hd__buf_12
Xoutput64 _3313_/Q vssd1 vssd1 vccd1 vccd1 io_out[4] sky130_fd_sc_hd__buf_12
Xoutput53 _3310_/Q vssd1 vssd1 vccd1 vccd1 io_out[21] sky130_fd_sc_hd__buf_12
XANTENNA__1714__B _2195_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1730__A _1889_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_38_wb_clk_i_A clkbuf_3_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_85_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2740_ _2714_/B _2740_/B vssd1 vssd1 vccd1 vccd1 _2740_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_26_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2671_ _3599_/Q _2868_/D vssd1 vssd1 vccd1 vccd1 _2851_/A sky130_fd_sc_hd__and2_1
X_1622_ _2480_/A vssd1 vssd1 vccd1 vccd1 _2479_/A sky130_fd_sc_hd__inv_4
XFILLER_0_1_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3223_ _3308_/CLK _3223_/D vssd1 vssd1 vccd1 vccd1 _3223_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1687__C1 _1979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3154_ hold838/X _3131_/X hold889/X _3103_/A vssd1 vssd1 vccd1 vccd1 _3154_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_27_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1640__A _3045_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3085_ _3085_/A0 _3084_/Y _3085_/S vssd1 vssd1 vccd1 vccd1 _3085_/X sky130_fd_sc_hd__mux2_1
X_2105_ _2570_/A _2365_/A vssd1 vssd1 vccd1 vccd1 _2111_/S sky130_fd_sc_hd__nand2_4
X_2036_ _2731_/A2 _2034_/X _2083_/B vssd1 vssd1 vccd1 vccd1 _2036_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_0_9_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout155_A _3172_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1837__S0 _2244_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2938_ _2941_/A _2931_/Y _2937_/Y _2944_/B vssd1 vssd1 vccd1 vccd1 _2938_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_17_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2869_ _2701_/B _2867_/X _2868_/X _2866_/Y vssd1 vssd1 vccd1 vccd1 _2869_/X sky130_fd_sc_hd__o31a_1
XFILLER_0_32_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold341 _3520_/Q vssd1 vssd1 vccd1 vccd1 hold341/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold352 _2284_/X vssd1 vssd1 vccd1 vccd1 _3299_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold330 _2493_/X vssd1 vssd1 vccd1 vccd1 _3446_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold396 _2600_/X vssd1 vssd1 vccd1 vccd1 _3535_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold385 _3671_/Q vssd1 vssd1 vccd1 vccd1 hold385/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold374 _2405_/X vssd1 vssd1 vccd1 vccd1 _3374_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold363 _3360_/Q vssd1 vssd1 vccd1 vccd1 hold363/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1030 _3687_/Q vssd1 vssd1 vccd1 vccd1 _3053_/A sky130_fd_sc_hd__buf_1
Xhold1041 _2318_/Y vssd1 vssd1 vccd1 vccd1 _2320_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1052 _2875_/X vssd1 vssd1 vccd1 vccd1 _3613_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1085 _3622_/Q vssd1 vssd1 vccd1 vccd1 _2941_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1693__A2 _2960_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1063 _3610_/Q vssd1 vssd1 vccd1 vccd1 _2998_/A1 sky130_fd_sc_hd__buf_1
Xhold1074 _3616_/Q vssd1 vssd1 vccd1 vccd1 _2964_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2365__B _2598_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2642__A1 _2091_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1828__S0 _1760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1905__B1 _2087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2556__A _3192_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2881__A1 _3613_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3772_ _3772_/A vssd1 vssd1 vccd1 vccd1 _3772_/X sky130_fd_sc_hd__buf_1
XFILLER_0_54_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2397__A0 _2658_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2723_ _2723_/A vssd1 vssd1 vccd1 vccd1 _2723_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_89_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2654_ _2654_/A _2654_/B vssd1 vssd1 vccd1 vccd1 _2660_/S sky130_fd_sc_hd__nand2_4
X_2585_ _2655_/A0 hold227/X _2590_/S vssd1 vssd1 vccd1 vccd1 _2585_/X sky130_fd_sc_hd__mux2_1
X_1605_ _2929_/A vssd1 vssd1 vccd1 vccd1 _1605_/Y sky130_fd_sc_hd__inv_2
Xfanout128 _1849_/S1 vssd1 vssd1 vccd1 vccd1 _2289_/C sky130_fd_sc_hd__buf_4
Xfanout106 _1630_/X vssd1 vssd1 vccd1 vccd1 _3045_/B sky130_fd_sc_hd__clkbuf_8
Xfanout117 _2480_/A vssd1 vssd1 vccd1 vccd1 _2228_/A sky130_fd_sc_hd__clkbuf_8
Xfanout139 _3346_/Q vssd1 vssd1 vccd1 vccd1 _1954_/S sky130_fd_sc_hd__buf_4
X_3206_ _3666_/CLK _3206_/D vssd1 vssd1 vccd1 vccd1 _3206_/Q sky130_fd_sc_hd__dfxtp_1
X_3137_ _3137_/A _3137_/B _3137_/C vssd1 vssd1 vccd1 vccd1 _3137_/X sky130_fd_sc_hd__or3_1
XANTENNA__2185__B _2244_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3068_ _3007_/A _3066_/X _3067_/X vssd1 vssd1 vccd1 vccd1 _3068_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_54_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2019_ _2479_/A _1991_/X _1998_/X _2018_/Y vssd1 vssd1 vccd1 vccd1 _2022_/B sky130_fd_sc_hd__a31o_1
XFILLER_0_92_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold171 _3432_/Q vssd1 vssd1 vccd1 vccd1 hold171/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold160 _2536_/X vssd1 vssd1 vccd1 vccd1 _3480_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold182 _2524_/X vssd1 vssd1 vccd1 vccd1 _3470_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold193 _3456_/Q vssd1 vssd1 vccd1 vccd1 hold193/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2091__A2 _2084_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2674__A_N _2868_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2370_ _3197_/A0 hold493/X _2371_/S vssd1 vssd1 vccd1 vccd1 _2370_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2985__S _2987_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3686_ _3692_/CLK _3686_/D vssd1 vssd1 vccd1 vccd1 _3686_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2706_ _2755_/B _2705_/B _2705_/C vssd1 vssd1 vccd1 vccd1 _2707_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2637_ _2658_/A0 hold661/X _2639_/S vssd1 vssd1 vccd1 vccd1 _2637_/X sky130_fd_sc_hd__mux2_1
Xscrapcpu_173 vssd1 vssd1 vccd1 vccd1 scrapcpu_173/HI io_out[31] sky130_fd_sc_hd__conb_1
Xscrapcpu_162 vssd1 vssd1 vccd1 vccd1 scrapcpu_162/HI io_oeb[8] sky130_fd_sc_hd__conb_1
XFILLER_0_64_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2568_ _2659_/A0 hold453/X _2569_/S vssd1 vssd1 vccd1 vccd1 _2568_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_10_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2499_ _2076_/A hold833/X _2499_/S vssd1 vssd1 vccd1 vccd1 _2499_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2196__A _2619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3022__A1 _3045_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_39_wb_clk_i clkbuf_3_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3723_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_clkbuf_3_5__f_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1870_ _1870_/A _1922_/B vssd1 vssd1 vccd1 vccd1 _2720_/C sky130_fd_sc_hd__or2_1
XANTENNA__1884__S _1937_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3540_ _3739_/CLK _3540_/D vssd1 vssd1 vccd1 vccd1 _3540_/Q sky130_fd_sc_hd__dfxtp_1
Xhold918 _3595_/Q vssd1 vssd1 vccd1 vccd1 hold918/X sky130_fd_sc_hd__clkbuf_2
Xhold907 _2922_/X vssd1 vssd1 vccd1 vccd1 _3620_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_51_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3471_ _3744_/CLK hold78/X vssd1 vssd1 vccd1 vccd1 hold77/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold929 _3680_/Q vssd1 vssd1 vccd1 vccd1 _3033_/A sky130_fd_sc_hd__dlygate4sd3_1
X_2422_ hold143/X _2655_/A0 _2427_/S vssd1 vssd1 vccd1 vccd1 _2422_/X sky130_fd_sc_hd__mux2_1
X_2353_ _2353_/A _2363_/B vssd1 vssd1 vccd1 vccd1 _2353_/X sky130_fd_sc_hd__or2_1
XFILLER_0_19_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2284_ _2355_/A hold351/X _2288_/S vssd1 vssd1 vccd1 vccd1 _2284_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1999_ _3391_/Q _3585_/Q _3567_/Q _3555_/Q _2000_/S0 _2289_/C vssd1 vssd1 vccd1 vccd1
+ _1999_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_70_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3738_ _3738_/CLK _3738_/D vssd1 vssd1 vccd1 vccd1 _3738_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3669_ _3670_/CLK _3669_/D vssd1 vssd1 vccd1 vccd1 _3669_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2279__C1 _3058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_3_6__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_3_6__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_38_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2506__A0 _3198_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2971_ hold409/X _3623_/Q _2999_/S vssd1 vssd1 vccd1 vccd1 _2971_/X sky130_fd_sc_hd__mux2_1
X_1922_ _1922_/A _1922_/B vssd1 vssd1 vccd1 vccd1 _2682_/C sky130_fd_sc_hd__or2_1
X_1853_ _3769_/A _2005_/S _2085_/C _1852_/Y vssd1 vssd1 vccd1 vccd1 _1853_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_71_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1908__A _2085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1784_ hold59/A _3479_/Q _3417_/Q _3429_/Q _2244_/B _2185_/C vssd1 vssd1 vccd1 vccd1
+ _1785_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_21_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold715 _3517_/Q vssd1 vssd1 vccd1 vccd1 hold715/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold704 _2621_/X vssd1 vssd1 vccd1 vccd1 _3553_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3523_ _3561_/CLK _3523_/D vssd1 vssd1 vccd1 vccd1 _3523_/Q sky130_fd_sc_hd__dfxtp_1
Xhold726 _2108_/X vssd1 vssd1 vccd1 vccd1 _3214_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold737 _3421_/Q vssd1 vssd1 vccd1 vccd1 hold737/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold748 _2380_/X vssd1 vssd1 vccd1 vccd1 _3352_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold759 _3656_/Q vssd1 vssd1 vccd1 vccd1 hold759/X sky130_fd_sc_hd__dlygate4sd3_1
X_3454_ _3737_/CLK _3454_/D vssd1 vssd1 vccd1 vccd1 _3454_/Q sky130_fd_sc_hd__dfxtp_1
X_2405_ _3197_/A0 hold373/X _2406_/S vssd1 vssd1 vccd1 vccd1 _2405_/X sky130_fd_sc_hd__mux2_1
X_3385_ _3654_/CLK _3385_/D vssd1 vssd1 vccd1 vccd1 _3385_/Q sky130_fd_sc_hd__dfxtp_1
X_2336_ _3197_/A0 hold411/X _2337_/S vssd1 vssd1 vccd1 vccd1 _2336_/X sky130_fd_sc_hd__mux2_1
X_2267_ _3058_/A _2245_/C _2022_/A vssd1 vssd1 vccd1 vccd1 _2278_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_27_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2198_ _2656_/A0 hold739/X _2202_/S vssd1 vssd1 vccd1 vccd1 _2198_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2193__B _2480_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_416 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout98_A _2987_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold31 hold31/A vssd1 vssd1 vccd1 vccd1 hold31/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold20 hold20/A vssd1 vssd1 vccd1 vccd1 hold20/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 hold53/A vssd1 vssd1 vccd1 vccd1 hold53/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 hold64/A vssd1 vssd1 vccd1 vccd1 hold64/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 hold42/A vssd1 vssd1 vccd1 vccd1 hold42/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 hold97/A vssd1 vssd1 vccd1 vccd1 hold97/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold86 hold86/A vssd1 vssd1 vccd1 vccd1 hold86/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 hold75/A vssd1 vssd1 vccd1 vccd1 hold75/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2087__C _2480_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2267__A2 _2245_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_28_wb_clk_i_A clkbuf_3_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_54_wb_clk_i clkbuf_leaf_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3637_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3170_ hold858/X _3158_/Y hold870/X _3172_/C1 vssd1 vssd1 vccd1 vccd1 _3170_/X sky130_fd_sc_hd__o211a_1
X_2121_ _3718_/Q _2149_/B vssd1 vssd1 vccd1 vccd1 _2146_/A sky130_fd_sc_hd__and2_1
X_2052_ _3118_/A _3048_/B vssd1 vssd1 vccd1 vccd1 _3157_/B sky130_fd_sc_hd__nor2_4
XANTENNA__2112__D1 _2014_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2954_ _2954_/A _2954_/B vssd1 vssd1 vccd1 vccd1 _2954_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_17_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2885_ _2885_/A _2885_/B hold801/X vssd1 vssd1 vccd1 vccd1 _2886_/A sky130_fd_sc_hd__or3b_4
X_1905_ _2244_/A _1900_/X _2087_/A vssd1 vssd1 vccd1 vccd1 _1905_/Y sky130_fd_sc_hd__o21ai_1
X_1836_ _1889_/A _1832_/Y _1834_/Y _1835_/Y vssd1 vssd1 vccd1 vccd1 _1836_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_32_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold501 _3357_/Q vssd1 vssd1 vccd1 vccd1 hold501/X sky130_fd_sc_hd__dlygate4sd3_1
X_1767_ _2819_/A _3130_/A vssd1 vssd1 vccd1 vccd1 _1767_/Y sky130_fd_sc_hd__nand2_2
Xhold545 _3367_/Q vssd1 vssd1 vccd1 vccd1 hold545/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold534 _2602_/X vssd1 vssd1 vccd1 vccd1 _3537_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3506_ _3545_/CLK _3506_/D vssd1 vssd1 vccd1 vccd1 _3506_/Q sky130_fd_sc_hd__dfxtp_1
Xhold512 _2639_/X vssd1 vssd1 vccd1 vccd1 _3569_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold523 _3739_/Q vssd1 vssd1 vccd1 vccd1 hold523/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold556 _2217_/X vssd1 vssd1 vccd1 vccd1 _3254_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold567 _3255_/Q vssd1 vssd1 vccd1 vccd1 hold567/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold578 _2287_/X vssd1 vssd1 vccd1 vccd1 _3302_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1698_ _1698_/A _2854_/B _1922_/B _1698_/D vssd1 vssd1 vccd1 vccd1 _1698_/X sky130_fd_sc_hd__or4_1
X_3437_ _3741_/CLK hold54/X vssd1 vssd1 vccd1 vccd1 hold53/A sky130_fd_sc_hd__dfxtp_1
Xhold589 _3665_/Q vssd1 vssd1 vccd1 vccd1 hold589/X sky130_fd_sc_hd__dlygate4sd3_1
X_3368_ _3543_/CLK _3368_/D vssd1 vssd1 vccd1 vccd1 _3368_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2319_ _3096_/A _2317_/X _2318_/B _2308_/Y vssd1 vssd1 vccd1 vccd1 _2320_/C sky130_fd_sc_hd__a211o_1
X_3299_ _3436_/CLK _3299_/D vssd1 vssd1 vccd1 vccd1 _3299_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2103__D1 _2228_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2957__A0 _2076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput21 _3770_/A vssd1 vssd1 vccd1 vccd1 io_oeb[12] sky130_fd_sc_hd__buf_12
Xoutput32 _3623_/Q vssd1 vssd1 vccd1 vccd1 io_oeb[33] sky130_fd_sc_hd__buf_12
Xoutput43 _3403_/Q vssd1 vssd1 vccd1 vccd1 io_out[12] sky130_fd_sc_hd__buf_12
XANTENNA__2379__A _2570_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput65 _3314_/Q vssd1 vssd1 vccd1 vccd1 io_out[5] sky130_fd_sc_hd__buf_12
Xoutput54 _3632_/Q vssd1 vssd1 vccd1 vccd1 io_out[22] sky130_fd_sc_hd__buf_12
XANTENNA__1791__S0 _2000_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2670_ _3626_/Q _3627_/Q _3628_/Q vssd1 vssd1 vccd1 vccd1 _2710_/A sky130_fd_sc_hd__or3_1
X_1621_ _1824_/A vssd1 vssd1 vccd1 vccd1 _2071_/A sky130_fd_sc_hd__inv_2
XFILLER_0_78_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_452 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2289__A _2289_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3222_ _3666_/CLK _3222_/D vssd1 vssd1 vccd1 vccd1 _3222_/Q sky130_fd_sc_hd__dfxtp_1
X_3153_ hold888/X _2886_/A _3137_/C vssd1 vssd1 vccd1 vccd1 _3153_/X sky130_fd_sc_hd__a21o_1
XANTENNA__1687__B1 _2854_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2104_ _2365_/A vssd1 vssd1 vccd1 vccd1 _3192_/A sky130_fd_sc_hd__inv_2
XFILLER_0_89_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3084_ _3677_/Q _3183_/B _3083_/X vssd1 vssd1 vccd1 vccd1 _3084_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_27_84 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1640__B _3048_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2035_ hold519/X _2731_/A2 _2701_/B _2034_/X vssd1 vssd1 vccd1 vccd1 _2035_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_49_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2100__A1 _2653_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1837__S1 _2185_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2937_ _2937_/A vssd1 vssd1 vccd1 vccd1 _2937_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2868_ _3630_/Q _2868_/B _2868_/C _2868_/D vssd1 vssd1 vccd1 vccd1 _2868_/X sky130_fd_sc_hd__or4_1
Xhold320 _2226_/X vssd1 vssd1 vccd1 vccd1 _3261_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1819_ _1819_/A _1819_/B vssd1 vssd1 vccd1 vccd1 _1819_/Y sky130_fd_sc_hd__nand2_1
X_2799_ _2861_/B _2730_/Y _2797_/Y _2798_/X _2859_/A vssd1 vssd1 vccd1 vccd1 _2799_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA__1914__A1 _2479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold342 _2582_/X vssd1 vssd1 vccd1 vccd1 _3520_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold353 _3435_/Q vssd1 vssd1 vccd1 vccd1 hold353/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold331 _3288_/Q vssd1 vssd1 vccd1 vccd1 hold331/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold375 _3674_/Q vssd1 vssd1 vccd1 vccd1 hold375/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold386 _2996_/X vssd1 vssd1 vccd1 vccd1 _3671_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold364 _2389_/X vssd1 vssd1 vccd1 vccd1 _3360_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold397 _3581_/Q vssd1 vssd1 vccd1 vccd1 hold397/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1042 _2320_/X vssd1 vssd1 vccd1 vccd1 _3313_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1031 _3052_/X vssd1 vssd1 vccd1 vccd1 _3055_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1020 _3625_/Q vssd1 vssd1 vccd1 vccd1 _2948_/A sky130_fd_sc_hd__buf_1
XANTENNA__2875__C1 _2859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1773__S0 _1981_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1075 _3614_/Q vssd1 vssd1 vccd1 vccd1 _2962_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1053 _3678_/Q vssd1 vssd1 vccd1 vccd1 _3027_/A sky130_fd_sc_hd__buf_1
Xhold1064 _3226_/Q vssd1 vssd1 vccd1 vccd1 _1707_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1086 _3597_/Q vssd1 vssd1 vccd1 vccd1 _2979_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1828__S1 _1760_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1905__A1 _2244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3771_ _3771_/A vssd1 vssd1 vccd1 vccd1 _3771_/X sky130_fd_sc_hd__buf_1
XFILLER_0_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2722_ _3626_/Q _3627_/Q _2741_/A vssd1 vssd1 vccd1 vccd1 _2723_/A sky130_fd_sc_hd__or3_2
XFILLER_0_14_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2653_ _2653_/A0 hold397/X _2653_/S vssd1 vssd1 vccd1 vccd1 _2653_/X sky130_fd_sc_hd__mux2_1
X_2584_ _2647_/A _2598_/B vssd1 vssd1 vccd1 vccd1 _2590_/S sky130_fd_sc_hd__nand2_2
X_1604_ _2876_/A vssd1 vssd1 vccd1 vccd1 _2885_/B sky130_fd_sc_hd__clkinv_4
Xfanout107 _1630_/X vssd1 vssd1 vccd1 vccd1 _3118_/A sky130_fd_sc_hd__clkbuf_4
Xfanout118 hold1071/X vssd1 vssd1 vccd1 vccd1 _2480_/A sky130_fd_sc_hd__buf_4
Xfanout129 _1849_/S1 vssd1 vssd1 vccd1 vccd1 _2014_/A sky130_fd_sc_hd__clkbuf_8
X_3205_ hold343/X _2363_/A _3205_/S vssd1 vssd1 vccd1 vccd1 _3205_/X sky130_fd_sc_hd__mux2_1
X_3136_ hold936/X _3131_/X hold953/X _3166_/C1 vssd1 vssd1 vccd1 vccd1 _3136_/X sky130_fd_sc_hd__o211a_1
X_3067_ _3097_/B _3063_/X _3064_/X _3124_/A vssd1 vssd1 vccd1 vccd1 _3067_/X sky130_fd_sc_hd__a31o_1
X_2018_ _2479_/A _2003_/X _2228_/B vssd1 vssd1 vccd1 vccd1 _2018_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__2185__C _2185_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold161 _3258_/Q vssd1 vssd1 vccd1 vccd1 hold161/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold150 _2516_/X vssd1 vssd1 vccd1 vccd1 _3463_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2560__A1 _3203_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold194 _2508_/X vssd1 vssd1 vccd1 vccd1 _3456_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold183 _3498_/Q vssd1 vssd1 vccd1 vccd1 hold183/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold172 _2475_/X vssd1 vssd1 vccd1 vccd1 _3432_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout80_A _2359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2848__C1 _2859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3000__B _3058_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1985__S0 _1988_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output61_A _2195_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1737__S0 _2000_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_9_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3737_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_3685_ _3695_/CLK _3685_/D vssd1 vssd1 vccd1 vccd1 _3685_/Q sky130_fd_sc_hd__dfxtp_1
X_2705_ _2755_/B _2705_/B _2705_/C vssd1 vssd1 vccd1 vccd1 _2707_/B sky130_fd_sc_hd__nand3_1
Xscrapcpu_174 vssd1 vssd1 vccd1 vccd1 scrapcpu_174/HI io_out[32] sky130_fd_sc_hd__conb_1
X_2636_ _3195_/A0 hold247/X _2639_/S vssd1 vssd1 vccd1 vccd1 _2636_/X sky130_fd_sc_hd__mux2_1
Xscrapcpu_163 vssd1 vssd1 vccd1 vccd1 scrapcpu_163/HI io_oeb[21] sky130_fd_sc_hd__conb_1
X_2567_ _2658_/A0 hold427/X _2569_/S vssd1 vssd1 vccd1 vccd1 _2567_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2498_ _2074_/A hold823/X _2499_/S vssd1 vssd1 vccd1 vccd1 _2498_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_3_5__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_3_5__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
X_3119_ hold817/X _3183_/B _3118_/X vssd1 vssd1 vccd1 vccd1 _3120_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_65_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3101__A _3103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1900__S0 _1954_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2533__A1 _2652_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3771__A _3771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1719__S0 _1981_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2221__A0 _2648_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold908 _3594_/Q vssd1 vssd1 vccd1 vccd1 hold908/X sky130_fd_sc_hd__buf_2
Xhold919 _2750_/X vssd1 vssd1 vccd1 vccd1 _3595_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_51_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3470_ _3743_/CLK _3470_/D vssd1 vssd1 vccd1 vccd1 _3470_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2524__A1 _2357_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2421_ _2633_/B _2612_/B vssd1 vssd1 vccd1 vccd1 _2427_/S sky130_fd_sc_hd__nor2_2
X_2352_ _2640_/A _2372_/A vssd1 vssd1 vccd1 vccd1 _2363_/B sky130_fd_sc_hd__or2_1
X_2283_ _2648_/A0 hold437/X _2288_/S vssd1 vssd1 vccd1 vccd1 _2283_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2288__A0 _2653_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout130_A _2185_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1998_ _2185_/A _1995_/Y _1997_/Y _2428_/C _1993_/Y vssd1 vssd1 vccd1 vccd1 _1998_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_0_42_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3737_ _3737_/CLK _3737_/D vssd1 vssd1 vccd1 vccd1 _3737_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3668_ _3668_/CLK _3668_/D vssd1 vssd1 vccd1 vccd1 _3668_/Q sky130_fd_sc_hd__dfxtp_1
X_2619_ _2619_/A _2654_/A vssd1 vssd1 vccd1 vccd1 _2625_/S sky130_fd_sc_hd__nand2_4
X_3599_ _3662_/CLK _3599_/D vssd1 vssd1 vccd1 vccd1 _3599_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__1949__S0 _2000_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2515__A1 _2655_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1823__B _2955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_18_wb_clk_i_A clkbuf_3_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_53_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2194__A_N _2479_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_57_wb_clk_i_A clkbuf_leaf_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_88_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2970_ hold313/X _3622_/Q _2999_/S vssd1 vssd1 vccd1 vccd1 _2970_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_29_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1921_ _1920_/B _1919_/X _1920_/Y _1922_/B vssd1 vssd1 vccd1 vccd1 _2682_/B sky130_fd_sc_hd__o211ai_4
XANTENNA__2993__A1 _2195_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1852_ _3328_/Q _2005_/S vssd1 vssd1 vccd1 vccd1 _1852_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_4_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1783_ _1889_/A _1778_/X _1782_/X _2087_/A vssd1 vssd1 vccd1 vccd1 _1783_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_0_52_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold727 _3487_/Q vssd1 vssd1 vccd1 vccd1 hold727/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold716 _2579_/X vssd1 vssd1 vccd1 vccd1 _3517_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3522_ _3558_/CLK _3522_/D vssd1 vssd1 vccd1 vccd1 _3522_/Q sky130_fd_sc_hd__dfxtp_1
Xhold705 _3221_/Q vssd1 vssd1 vccd1 vccd1 hold705/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold738 _2462_/X vssd1 vssd1 vccd1 vccd1 _3421_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold749 _3247_/Q vssd1 vssd1 vccd1 vccd1 hold749/X sky130_fd_sc_hd__dlygate4sd3_1
X_3453_ _3496_/CLK _3453_/D vssd1 vssd1 vccd1 vccd1 _3453_/Q sky130_fd_sc_hd__dfxtp_1
X_2404_ _3196_/A0 hold695/X _2406_/S vssd1 vssd1 vccd1 vccd1 _2404_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_20_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3384_ _3419_/CLK _3384_/D vssd1 vssd1 vccd1 vccd1 _3384_/Q sky130_fd_sc_hd__dfxtp_1
X_2335_ _3196_/A0 hold305/X _2337_/S vssd1 vssd1 vccd1 vccd1 _2335_/X sky130_fd_sc_hd__mux2_1
X_2266_ _3198_/A0 hold405/X _2266_/S vssd1 vssd1 vccd1 vccd1 _2266_/X sky130_fd_sc_hd__mux2_1
X_2197_ _2089_/X hold601/X _2202_/S vssd1 vssd1 vccd1 vccd1 _2197_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_87_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1834__A _2245_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold10 hold10/A vssd1 vssd1 vccd1 vccd1 hold10/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 hold32/A vssd1 vssd1 vccd1 vccd1 hold32/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 hold21/A vssd1 vssd1 vccd1 vccd1 hold21/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 hold43/A vssd1 vssd1 vccd1 vccd1 hold43/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 hold54/A vssd1 vssd1 vccd1 vccd1 hold54/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 hold65/A vssd1 vssd1 vccd1 vccd1 hold65/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold98 hold98/A vssd1 vssd1 vccd1 vccd1 hold98/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 hold87/A vssd1 vssd1 vccd1 vccd1 hold87/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 hold76/A vssd1 vssd1 vccd1 vccd1 hold76/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2975__A1 _3613_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2360__C1 _3172_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_23_wb_clk_i clkbuf_3_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3743_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_2120_ _3717_/Q _3716_/Q _3715_/Q vssd1 vssd1 vccd1 vccd1 _2149_/B sky130_fd_sc_hd__and3_1
XFILLER_0_83_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2051_ _2031_/Y _2049_/X _2050_/X _2495_/A vssd1 vssd1 vccd1 vccd1 _3349_/D sky130_fd_sc_hd__o211a_1
XANTENNA__2112__C1 _2085_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2953_ hold860/X _1685_/B _2876_/X _1979_/A vssd1 vssd1 vccd1 vccd1 _2954_/B sky130_fd_sc_hd__o31a_1
XFILLER_0_84_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1769__A2 _2731_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1904_ _3770_/A _2005_/S _2085_/C _1903_/Y vssd1 vssd1 vccd1 vccd1 _1904_/X sky130_fd_sc_hd__a211o_1
X_2884_ hold249/X _2940_/B2 _2701_/B _1712_/A vssd1 vssd1 vccd1 vccd1 _2884_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_0_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1835_ _1889_/A _1830_/X _2087_/A vssd1 vssd1 vccd1 vccd1 _1835_/Y sky130_fd_sc_hd__o21ai_1
Xhold502 _2385_/X vssd1 vssd1 vccd1 vccd1 _3357_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1766_ _2876_/B _2846_/B vssd1 vssd1 vccd1 vccd1 _1766_/Y sky130_fd_sc_hd__nor2_1
Xhold535 _3239_/Q vssd1 vssd1 vccd1 vccd1 hold535/X sky130_fd_sc_hd__dlygate4sd3_1
X_3505_ _3543_/CLK _3505_/D vssd1 vssd1 vccd1 vccd1 _3505_/Q sky130_fd_sc_hd__dfxtp_1
Xhold513 _3265_/Q vssd1 vssd1 vccd1 vccd1 hold513/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold524 _3198_/X vssd1 vssd1 vccd1 vccd1 _3739_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold557 _3538_/Q vssd1 vssd1 vccd1 vccd1 hold557/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold579 _3559_/Q vssd1 vssd1 vccd1 vccd1 hold579/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold546 _2397_/X vssd1 vssd1 vccd1 vccd1 _3367_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold568 _2218_/X vssd1 vssd1 vccd1 vccd1 _3255_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1697_ _1653_/C _1713_/B _1696_/Y vssd1 vssd1 vccd1 vccd1 _1698_/D sky130_fd_sc_hd__o21ai_1
XFILLER_0_40_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3436_ _3436_/CLK _3436_/D vssd1 vssd1 vccd1 vccd1 _3436_/Q sky130_fd_sc_hd__dfxtp_1
X_3367_ _3585_/CLK _3367_/D vssd1 vssd1 vccd1 vccd1 _3367_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2318_ hold1040/X _2318_/B vssd1 vssd1 vccd1 vccd1 _2318_/Y sky130_fd_sc_hd__nand2b_1
X_3298_ _3581_/CLK _3298_/D vssd1 vssd1 vccd1 vccd1 _3298_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2249_ hold45/X _2650_/A0 _2252_/S vssd1 vssd1 vccd1 vccd1 hold46/A sky130_fd_sc_hd__mux2_1
XANTENNA__2103__C1 _2195_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2406__A0 _3198_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput22 _3771_/X vssd1 vssd1 vccd1 vccd1 io_oeb[13] sky130_fd_sc_hd__buf_12
Xoutput33 _3624_/Q vssd1 vssd1 vccd1 vccd1 io_oeb[34] sky130_fd_sc_hd__buf_12
Xoutput55 _3328_/Q vssd1 vssd1 vccd1 vccd1 io_out[23] sky130_fd_sc_hd__buf_12
XFILLER_0_9_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput66 _3315_/Q vssd1 vssd1 vccd1 vccd1 io_out[6] sky130_fd_sc_hd__buf_12
Xoutput44 _3404_/Q vssd1 vssd1 vccd1 vccd1 io_out[13] sky130_fd_sc_hd__buf_12
XANTENNA__1791__S1 _2219_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1620_ _3058_/A vssd1 vssd1 vccd1 vccd1 _1620_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_22_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3221_ _3308_/CLK _3221_/D vssd1 vssd1 vccd1 vccd1 _3221_/Q sky130_fd_sc_hd__dfxtp_1
X_3152_ _3152_/A1 _3131_/X _3151_/X _3103_/A vssd1 vssd1 vccd1 vccd1 _3152_/X sky130_fd_sc_hd__o211a_1
XANTENNA__1687__A1 _2797_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2884__B1 _2701_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2103_ _2084_/A _2084_/B _2479_/A _2195_/B _2228_/C vssd1 vssd1 vccd1 vccd1 _2365_/A
+ sky130_fd_sc_hd__o2111a_4
XFILLER_0_89_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3083_ _3076_/Y _3082_/X _3118_/A vssd1 vssd1 vccd1 vccd1 _3083_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_27_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2636__A0 _3195_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2034_ _2854_/A _2034_/B _2082_/C _2789_/S vssd1 vssd1 vccd1 vccd1 _2034_/X sky130_fd_sc_hd__or4_4
XFILLER_0_9_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2936_ _2885_/B _2934_/X _2935_/Y _2941_/A vssd1 vssd1 vccd1 vccd1 _2937_/A sky130_fd_sc_hd__o2bb2a_1
X_2867_ _2867_/A _2867_/B _2867_/C vssd1 vssd1 vccd1 vccd1 _2867_/X sky130_fd_sc_hd__or3_1
XFILLER_0_32_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1818_ _2999_/A1 _1769_/Y _1817_/X _2854_/B vssd1 vssd1 vccd1 vccd1 _1819_/B sky130_fd_sc_hd__o22ai_1
XFILLER_0_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold310 _2426_/X vssd1 vssd1 vccd1 vccd1 _3392_/D sky130_fd_sc_hd__dlygate4sd3_1
X_2798_ _2797_/A hold565/X _2731_/X vssd1 vssd1 vccd1 vccd1 _2798_/X sky130_fd_sc_hd__a21o_1
Xhold343 _3745_/Q vssd1 vssd1 vccd1 vccd1 hold343/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold321 _3497_/Q vssd1 vssd1 vccd1 vccd1 hold321/X sky130_fd_sc_hd__dlygate4sd3_1
X_1749_ _2085_/A _1749_/B vssd1 vssd1 vccd1 vccd1 _1749_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_13_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold332 _2263_/X vssd1 vssd1 vccd1 vccd1 _3288_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold387 _3591_/Q vssd1 vssd1 vccd1 vccd1 hold387/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold376 _2999_/X vssd1 vssd1 vccd1 vccd1 _3674_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold354 _2478_/X vssd1 vssd1 vccd1 vccd1 _3435_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold365 _3219_/Q vssd1 vssd1 vccd1 vccd1 hold365/X sky130_fd_sc_hd__dlygate4sd3_1
X_3419_ _3419_/CLK _3419_/D vssd1 vssd1 vccd1 vccd1 _3419_/Q sky130_fd_sc_hd__dfxtp_1
Xhold398 _2653_/X vssd1 vssd1 vccd1 vccd1 _3581_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1032 _3055_/X vssd1 vssd1 vccd1 vccd1 _3687_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1010 _3225_/Q vssd1 vssd1 vccd1 vccd1 _2153_/A sky130_fd_sc_hd__buf_2
Xhold1021 _3351_/Q vssd1 vssd1 vccd1 vccd1 hold1021/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1773__S1 _2219_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1065 _3609_/Q vssd1 vssd1 vccd1 vccd1 _2997_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1076 _3603_/Q vssd1 vssd1 vccd1 vccd1 _2985_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1054 _3027_/Y vssd1 vssd1 vccd1 vccd1 _3028_/C sky130_fd_sc_hd__dlygate4sd3_1
Xhold1043 _3295_/Q vssd1 vssd1 vccd1 vccd1 _2274_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1087 _3311_/Q vssd1 vssd1 vccd1 vccd1 hold932/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_67_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3774__A _3774_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2866__B1 _3613_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2094__A1 _2650_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3770_ _3770_/A vssd1 vssd1 vccd1 vccd1 _3770_/X sky130_fd_sc_hd__buf_1
X_2721_ _2759_/B _2736_/B vssd1 vssd1 vccd1 vccd1 _2721_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_14_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2652_ _2652_/A0 hold383/X _2653_/S vssd1 vssd1 vccd1 vccd1 _2652_/X sky130_fd_sc_hd__mux2_1
X_2583_ _2660_/A0 hold443/X _2583_/S vssd1 vssd1 vccd1 vccd1 _2583_/X sky130_fd_sc_hd__mux2_1
X_1603_ _2309_/A vssd1 vssd1 vccd1 vccd1 _3014_/A sky130_fd_sc_hd__inv_2
XFILLER_0_10_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout108 wire109/X vssd1 vssd1 vccd1 vccd1 _3183_/B sky130_fd_sc_hd__buf_4
Xfanout119 hold1033/X vssd1 vssd1 vccd1 vccd1 _2228_/C sky130_fd_sc_hd__buf_6
X_3204_ hold593/X _2361_/A _3205_/S vssd1 vssd1 vccd1 vccd1 _3204_/X sky130_fd_sc_hd__mux2_1
X_3135_ _2892_/A _2886_/A _3137_/C vssd1 vssd1 vccd1 vccd1 _3135_/X sky130_fd_sc_hd__a21o_1
Xclkbuf_3_4__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_9_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__2609__A0 _2658_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3066_ _3037_/D _3075_/B _3018_/X vssd1 vssd1 vccd1 vccd1 _3066_/X sky130_fd_sc_hd__o21a_1
XANTENNA__2185__D _2480_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2017_ _2289_/A _2014_/Y _2016_/Y _2087_/A _2012_/Y vssd1 vssd1 vccd1 vccd1 _2017_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_0_54_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2919_ _2924_/B _2924_/C vssd1 vssd1 vccd1 vccd1 _2919_/X sky130_fd_sc_hd__and2_1
XFILLER_0_45_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold151 _3574_/Q vssd1 vssd1 vccd1 vccd1 hold151/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold162 _2223_/X vssd1 vssd1 vccd1 vccd1 _3258_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold140 _2476_/X vssd1 vssd1 vccd1 vccd1 _3433_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 _3532_/Q vssd1 vssd1 vccd1 vccd1 hold173/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold184 _2557_/X vssd1 vssd1 vccd1 vccd1 _3498_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 _3256_/Q vssd1 vssd1 vccd1 vccd1 hold195/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1842__A _2006_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout73_A _2653_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1988__S _1988_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3769__A _3769_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2784__C1 _2859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1985__S1 _2185_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1737__S1 _2219_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output54_A _3632_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2067__A1 _2074_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1814__A1 input11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3684_ _3695_/CLK _3684_/D vssd1 vssd1 vccd1 vccd1 _3684_/Q sky130_fd_sc_hd__dfxtp_1
X_2704_ _2755_/B _2704_/B _2755_/C vssd1 vssd1 vccd1 vccd1 _2762_/A sky130_fd_sc_hd__and3_1
XFILLER_0_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2635_ _2656_/A0 hold795/X _2639_/S vssd1 vssd1 vccd1 vccd1 _2635_/X sky130_fd_sc_hd__mux2_1
Xscrapcpu_164 vssd1 vssd1 vccd1 vccd1 scrapcpu_164/HI io_oeb[22] sky130_fd_sc_hd__conb_1
Xscrapcpu_175 vssd1 vssd1 vccd1 vccd1 scrapcpu_175/HI io_out[33] sky130_fd_sc_hd__conb_1
X_2566_ _3195_/A0 hold627/X _2569_/S vssd1 vssd1 vccd1 vccd1 _2566_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_10_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2497_ _2497_/A _2955_/B vssd1 vssd1 vccd1 vccd1 _2499_/S sky130_fd_sc_hd__or2_1
XFILLER_0_4_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3118_ _3118_/A _3118_/B vssd1 vssd1 vccd1 vccd1 _3118_/X sky130_fd_sc_hd__or2_1
X_3049_ _3118_/A _3124_/B _3047_/X _3037_/C _3055_/A vssd1 vssd1 vccd1 vccd1 _3049_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_0_92_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1900__S1 _2014_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_47_wb_clk_i_A clkbuf_3_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__2297__A1 _3048_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1719__S1 _1981_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2049__A1 _2228_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_48_wb_clk_i clkbuf_3_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3646_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_28_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout90 _2091_/X vssd1 vssd1 vccd1 vccd1 _2355_/A sky130_fd_sc_hd__buf_4
XFILLER_0_10_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold909 _2733_/X vssd1 vssd1 vccd1 vccd1 _3594_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_51_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2420_ hold217/X _3198_/A0 _2420_/S vssd1 vssd1 vccd1 vccd1 _2420_/X sky130_fd_sc_hd__mux2_1
X_2351_ _2640_/A _2372_/A vssd1 vssd1 vccd1 vccd1 _2351_/Y sky130_fd_sc_hd__nor2_2
X_2282_ _2654_/B _2647_/B vssd1 vssd1 vccd1 vccd1 _2288_/S sky130_fd_sc_hd__nand2_2
XFILLER_0_59_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1799__B1 _2085_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1997_ _2006_/A _1997_/B vssd1 vssd1 vccd1 vccd1 _1997_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_34_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout123_A _2289_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3736_ _3739_/CLK _3736_/D vssd1 vssd1 vccd1 vccd1 _3736_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3667_ _3676_/CLK _3667_/D vssd1 vssd1 vccd1 vccd1 _3667_/Q sky130_fd_sc_hd__dfxtp_1
X_2618_ hold71/X _2099_/X _2618_/S vssd1 vssd1 vccd1 vccd1 hold72/A sky130_fd_sc_hd__mux2_1
X_3598_ _3655_/CLK _3598_/D vssd1 vssd1 vccd1 vccd1 _3598_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1949__S1 _2219_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2549_ _2549_/A _2612_/B vssd1 vssd1 vccd1 vccd1 _2555_/S sky130_fd_sc_hd__nor2_2
XANTENNA__2488__A _2570_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2279__A1 _1716_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2951__A _3103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_3_wb_clk_i_A clkbuf_leaf_5_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2442__A1 _2652_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1876__S0 _1760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1920_ input1/X _1920_/B vssd1 vssd1 vccd1 vccd1 _1920_/Y sky130_fd_sc_hd__nand2_1
X_1851_ _2085_/C _1851_/B vssd1 vssd1 vccd1 vccd1 _1851_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_21_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1782_ _2006_/A _1779_/X _1781_/X vssd1 vssd1 vccd1 vccd1 _1782_/X sky130_fd_sc_hd__a21o_1
X_3521_ _3545_/CLK _3521_/D vssd1 vssd1 vccd1 vccd1 _3521_/Q sky130_fd_sc_hd__dfxtp_1
Xhold728 _2544_/X vssd1 vssd1 vccd1 vccd1 _3487_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold706 _2117_/X vssd1 vssd1 vccd1 vccd1 _3221_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold717 _3408_/Q vssd1 vssd1 vccd1 vccd1 hold717/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold739 _3236_/Q vssd1 vssd1 vccd1 vccd1 hold739/X sky130_fd_sc_hd__dlygate4sd3_1
X_3452_ _3570_/CLK _3452_/D vssd1 vssd1 vccd1 vccd1 _3452_/Q sky130_fd_sc_hd__dfxtp_1
X_2403_ _2475_/A1 hold653/X _2406_/S vssd1 vssd1 vccd1 vccd1 _2403_/X sky130_fd_sc_hd__mux2_1
X_3383_ _3419_/CLK _3383_/D vssd1 vssd1 vccd1 vccd1 _3383_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2101__A _2245_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2334_ _3195_/A0 hold745/X _2337_/S vssd1 vssd1 vccd1 vccd1 _2334_/X sky130_fd_sc_hd__mux2_1
X_2265_ _3197_/A0 hold479/X _2266_/S vssd1 vssd1 vccd1 vccd1 _2265_/X sky130_fd_sc_hd__mux2_1
X_2196_ _2619_/A _2407_/A vssd1 vssd1 vccd1 vccd1 _2202_/S sky130_fd_sc_hd__nand2_2
XFILLER_0_46_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2433__A1 _2357_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2197__A0 _2089_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3719_ _3721_/CLK _3719_/D vssd1 vssd1 vccd1 vccd1 _3719_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold11 hold11/A vssd1 vssd1 vccd1 vccd1 hold11/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold22 hold22/A vssd1 vssd1 vccd1 vccd1 hold22/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 hold33/A vssd1 vssd1 vccd1 vccd1 hold33/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 hold44/A vssd1 vssd1 vccd1 vccd1 hold44/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2946__A _3103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold55 hold55/A vssd1 vssd1 vccd1 vccd1 hold55/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 hold77/A vssd1 vssd1 vccd1 vccd1 hold77/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 hold99/A vssd1 vssd1 vccd1 vccd1 hold99/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 hold88/A vssd1 vssd1 vccd1 vccd1 hold88/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 hold66/A vssd1 vssd1 vccd1 vccd1 hold66/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2424__A1 _3195_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3082__D1 _3048_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1744__B _2244_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1760__A _1760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2050_ _2050_/A _2050_/B vssd1 vssd1 vccd1 vccd1 _2050_/X sky130_fd_sc_hd__or2_1
XFILLER_0_88_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2112__B1 _2244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2663__A1 _3201_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2591__A _2640_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2952_ _1685_/B _2876_/X hold860/X vssd1 vssd1 vccd1 vccd1 _2952_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__2415__A1 _3193_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1849__S0 _1954_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1903_ _3329_/Q _2005_/S vssd1 vssd1 vccd1 vccd1 _1903_/Y sky130_fd_sc_hd__nor2_1
X_2883_ _3130_/B hold998/X _2877_/X vssd1 vssd1 vccd1 vccd1 _2883_/Y sky130_fd_sc_hd__a21boi_4
XFILLER_0_32_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1834_ _2245_/B _1834_/B vssd1 vssd1 vccd1 vccd1 _1834_/Y sky130_fd_sc_hd__nand2_1
X_1765_ hold823/X _1922_/B _1763_/X _1764_/X vssd1 vssd1 vccd1 vccd1 _2868_/C sky130_fd_sc_hd__o22a_4
Xhold536 _2201_/X vssd1 vssd1 vccd1 vccd1 _3239_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold525 _3468_/Q vssd1 vssd1 vccd1 vccd1 hold525/X sky130_fd_sc_hd__dlygate4sd3_1
X_3504_ _3739_/CLK _3504_/D vssd1 vssd1 vccd1 vccd1 _3504_/Q sky130_fd_sc_hd__dfxtp_1
Xhold514 _2234_/X vssd1 vssd1 vccd1 vccd1 _3265_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold503 _3300_/Q vssd1 vssd1 vccd1 vccd1 hold503/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold558 _2603_/X vssd1 vssd1 vccd1 vccd1 _3538_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold547 _3512_/Q vssd1 vssd1 vccd1 vccd1 hold547/X sky130_fd_sc_hd__dlygate4sd3_1
X_1696_ _2876_/B _3130_/A vssd1 vssd1 vccd1 vccd1 _1696_/Y sky130_fd_sc_hd__nor2_4
Xhold569 _3654_/Q vssd1 vssd1 vccd1 vccd1 hold569/X sky130_fd_sc_hd__dlygate4sd3_1
X_3435_ _3665_/CLK _3435_/D vssd1 vssd1 vccd1 vccd1 _3435_/Q sky130_fd_sc_hd__dfxtp_1
X_3366_ _3575_/CLK _3366_/D vssd1 vssd1 vccd1 vccd1 _3366_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2317_ hold936/X _3089_/B _2316_/Y _3152_/A1 _2314_/X vssd1 vssd1 vccd1 vccd1 _2317_/X
+ sky130_fd_sc_hd__a221o_1
X_3297_ _3447_/CLK _3297_/D vssd1 vssd1 vccd1 vccd1 _3297_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1670__A _2885_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2248_ hold75/X _2355_/A _2252_/S vssd1 vssd1 vccd1 vccd1 hold76/A sky130_fd_sc_hd__mux2_1
XANTENNA__2103__B1 _2479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2179_ _2173_/Y _2177_/Y _2178_/X _2169_/B vssd1 vssd1 vccd1 vccd1 _2179_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_63_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2006__A _2006_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2590__A0 _2363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput23 _3771_/A vssd1 vssd1 vccd1 vccd1 io_oeb[14] sky130_fd_sc_hd__buf_12
Xoutput34 _3625_/Q vssd1 vssd1 vccd1 vccd1 io_oeb[35] sky130_fd_sc_hd__buf_12
XFILLER_0_31_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput56 _3329_/Q vssd1 vssd1 vccd1 vccd1 io_out[24] sky130_fd_sc_hd__buf_12
Xoutput67 _3690_/Q vssd1 vssd1 vccd1 vccd1 io_out[7] sky130_fd_sc_hd__buf_12
Xoutput45 _3405_/Q vssd1 vssd1 vccd1 vccd1 io_out[14] sky130_fd_sc_hd__buf_12
XANTENNA__2893__A1 _2876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2645__A1 _2659_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1755__A _2479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2581__A0 _2658_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3220_ _3666_/CLK _3220_/D vssd1 vssd1 vccd1 vccd1 _3220_/Q sky130_fd_sc_hd__dfxtp_1
X_3151_ _3623_/Q _2886_/A _3137_/C vssd1 vssd1 vccd1 vccd1 _3151_/X sky130_fd_sc_hd__a21o_1
Xclkbuf_3_3__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_3_3__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
X_2102_ _3348_/Q _2244_/B _2244_/C vssd1 vssd1 vccd1 vccd1 _2570_/A sky130_fd_sc_hd__and3_4
XANTENNA__1687__A2 _2960_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2884__B2 _1712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3082_ _1638_/A _1821_/X _3158_/B _2301_/C _3048_/B vssd1 vssd1 vccd1 vccd1 _3082_/X
+ sky130_fd_sc_hd__a2111o_1
X_2033_ _2741_/A _2742_/B vssd1 vssd1 vccd1 vccd1 _2789_/S sky130_fd_sc_hd__or2_2
XFILLER_0_43_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2935_ _2935_/A _2935_/B vssd1 vssd1 vccd1 vccd1 _2935_/Y sky130_fd_sc_hd__nand2_1
X_2866_ _3630_/Q _2868_/B _3613_/Q vssd1 vssd1 vccd1 vccd1 _2866_/Y sky130_fd_sc_hd__o21ai_1
X_1817_ hold375/X _2731_/A2 _2868_/D _1713_/X vssd1 vssd1 vccd1 vccd1 _1817_/X sky130_fd_sc_hd__o22a_1
Xhold300 _2646_/X vssd1 vssd1 vccd1 vccd1 _3575_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2797_ _2797_/A _2797_/B vssd1 vssd1 vccd1 vccd1 _2797_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold311 _3210_/Q vssd1 vssd1 vccd1 vccd1 hold311/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2572__A0 _3201_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold344 _3205_/X vssd1 vssd1 vccd1 vccd1 _3745_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold322 _2555_/X vssd1 vssd1 vccd1 vccd1 _3497_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1748_ hold89/A hold1/A _3210_/Q _3222_/Q _2085_/B _2014_/A vssd1 vssd1 vccd1 vccd1
+ _1749_/B sky130_fd_sc_hd__mux4_1
Xhold333 _3419_/Q vssd1 vssd1 vccd1 vccd1 hold333/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold355 _3380_/Q vssd1 vssd1 vccd1 vccd1 hold355/X sky130_fd_sc_hd__dlygate4sd3_1
X_1679_ _2846_/B _2876_/C _1679_/C vssd1 vssd1 vccd1 vccd1 _2878_/B sky130_fd_sc_hd__and3_1
Xhold377 _3263_/Q vssd1 vssd1 vccd1 vccd1 hold377/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold366 _2115_/X vssd1 vssd1 vccd1 vccd1 _3219_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold388 _2665_/X vssd1 vssd1 vccd1 vccd1 _3591_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold399 _3371_/Q vssd1 vssd1 vccd1 vccd1 hold399/X sky130_fd_sc_hd__dlygate4sd3_1
X_3418_ _3636_/CLK _3418_/D vssd1 vssd1 vccd1 vccd1 _3418_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1000 _3227_/Q vssd1 vssd1 vccd1 vccd1 _3059_/B sky130_fd_sc_hd__clkbuf_2
X_3349_ _3636_/CLK _3349_/D vssd1 vssd1 vccd1 vccd1 _3349_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1022 _2072_/X vssd1 vssd1 vccd1 vccd1 _3351_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1011 _2170_/Y vssd1 vssd1 vccd1 vccd1 _2171_/B1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1033 _3349_/Q vssd1 vssd1 vccd1 vccd1 hold1033/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1066 _2938_/X vssd1 vssd1 vccd1 vccd1 _2939_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1055 _3028_/X vssd1 vssd1 vccd1 vccd1 _3678_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1044 _2275_/X vssd1 vssd1 vccd1 vccd1 _3295_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2627__A1 _2089_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1077 _3605_/Q vssd1 vssd1 vccd1 vccd1 _2987_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1088 _3615_/Q vssd1 vssd1 vccd1 vccd1 hold952/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2618__A1 _2099_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2720_ _3594_/Q _2720_/B _2720_/C vssd1 vssd1 vccd1 vccd1 _2736_/B sky130_fd_sc_hd__and3_1
X_2651_ _2651_/A0 hold455/X _2653_/S vssd1 vssd1 vccd1 vccd1 _2651_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1602_ _3053_/B vssd1 vssd1 vccd1 vccd1 _3097_/A sky130_fd_sc_hd__inv_2
X_2582_ _2659_/A0 hold341/X _2583_/S vssd1 vssd1 vccd1 vccd1 _2582_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_22_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3203_ hold421/X _3203_/A1 _3205_/S vssd1 vssd1 vccd1 vccd1 _3203_/X sky130_fd_sc_hd__mux2_1
X_3134_ hold898/X _3131_/X _3133_/X _3166_/C1 vssd1 vssd1 vccd1 vccd1 _3134_/X sky130_fd_sc_hd__o211a_1
X_3065_ _3065_/A _3687_/Q _3686_/Q vssd1 vssd1 vccd1 vccd1 _3075_/B sky130_fd_sc_hd__or3_1
X_2016_ _2085_/C _2016_/B vssd1 vssd1 vccd1 vccd1 _2016_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__2255__S _2259_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout153_A _3172_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2918_ _1712_/A _3606_/Q hold199/X _2940_/B2 vssd1 vssd1 vccd1 vccd1 _2918_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_0_9_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2849_ _2803_/A _2711_/Y _2805_/X vssd1 vssd1 vccd1 vccd1 _2849_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__2545__A0 _2357_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold130 _2255_/X vssd1 vssd1 vccd1 vccd1 _3281_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold141 _3499_/Q vssd1 vssd1 vccd1 vccd1 hold141/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold152 _2645_/X vssd1 vssd1 vccd1 vccd1 _3574_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_37_wb_clk_i_A clkbuf_3_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold174 _2596_/X vssd1 vssd1 vccd1 vccd1 _3532_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold163 _3592_/Q vssd1 vssd1 vccd1 vccd1 hold163/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold185 _3280_/Q vssd1 vssd1 vccd1 vccd1 hold185/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold196 _2221_/X vssd1 vssd1 vccd1 vccd1 _3256_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1814__A2 _2022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3683_ _3695_/CLK _3683_/D vssd1 vssd1 vccd1 vccd1 _3683_/Q sky130_fd_sc_hd__dfxtp_1
X_2703_ _2754_/A _2735_/A _2703_/C vssd1 vssd1 vccd1 vccd1 _2755_/C sky130_fd_sc_hd__or3_1
XFILLER_0_71_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2634_ _2655_/A0 hold631/X _2639_/S vssd1 vssd1 vccd1 vccd1 _2634_/X sky130_fd_sc_hd__mux2_1
Xscrapcpu_165 vssd1 vssd1 vccd1 vccd1 scrapcpu_165/HI io_oeb[23] sky130_fd_sc_hd__conb_1
Xscrapcpu_176 vssd1 vssd1 vccd1 vccd1 scrapcpu_176/HI io_out[34] sky130_fd_sc_hd__conb_1
X_2565_ _2656_/A0 hold643/X _2569_/S vssd1 vssd1 vccd1 vccd1 _2565_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_10_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2496_ _3243_/Q _3045_/B _2496_/C _2495_/X vssd1 vssd1 vccd1 vccd1 _2955_/B sky130_fd_sc_hd__or4b_1
XFILLER_0_65_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3117_ hold817/X _3120_/A _3116_/X _3055_/A vssd1 vssd1 vccd1 vccd1 _3117_/X sky130_fd_sc_hd__o211a_1
X_3048_ _3183_/B _3048_/B _3053_/C vssd1 vssd1 vccd1 vccd1 _3048_/X sky130_fd_sc_hd__and3_1
XFILLER_0_92_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2766__B1 _2731_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2014__A _2014_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout91 _2091_/X vssd1 vssd1 vccd1 vccd1 _3201_/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout80 _2359_/A vssd1 vssd1 vccd1 vccd1 _3196_/A0 sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_17_wb_clk_i clkbuf_3_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3585_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__2859__A _2859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_390 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2350_ _3108_/A _2350_/B vssd1 vssd1 vccd1 vccd1 _3327_/D sky130_fd_sc_hd__or2_1
X_2281_ _2647_/B vssd1 vssd1 vccd1 vccd1 _2372_/A sky130_fd_sc_hd__inv_2
XFILLER_0_19_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1799__A1 _3774_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1938__A _2245_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1996_ _3459_/Q _3591_/Q _1996_/S vssd1 vssd1 vccd1 vccd1 _1997_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_70_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3735_ _3735_/CLK _3735_/D vssd1 vssd1 vccd1 vccd1 _3735_/Q sky130_fd_sc_hd__dfxtp_1
X_3666_ _3666_/CLK _3666_/D vssd1 vssd1 vccd1 vccd1 _3666_/Q sky130_fd_sc_hd__dfxtp_1
X_2617_ hold7/X _2659_/A0 _2618_/S vssd1 vssd1 vccd1 vccd1 hold8/A sky130_fd_sc_hd__mux2_1
XFILLER_0_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3597_ _3655_/CLK _3597_/D vssd1 vssd1 vccd1 vccd1 _3597_/Q sky130_fd_sc_hd__dfxtp_2
X_2548_ _2363_/A hold669/X _2548_/S vssd1 vssd1 vccd1 vccd1 _2548_/X sky130_fd_sc_hd__mux2_1
X_2479_ _2479_/A _2479_/B _2479_/C vssd1 vssd1 vccd1 vccd1 _2598_/B sky130_fd_sc_hd__and3_4
XANTENNA__2279__A2 _2480_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1876__S1 _1981_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1850_ _3340_/Q _3298_/Q _1954_/S vssd1 vssd1 vccd1 vccd1 _1851_/B sky130_fd_sc_hd__mux2_1
X_1781_ _2245_/B _1780_/X _2289_/A vssd1 vssd1 vccd1 vccd1 _1781_/X sky130_fd_sc_hd__a21o_1
X_3520_ _3545_/CLK _3520_/D vssd1 vssd1 vccd1 vccd1 _3520_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold707 _3653_/Q vssd1 vssd1 vccd1 vccd1 hold707/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold718 _2447_/X vssd1 vssd1 vccd1 vccd1 _3408_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold729 _3490_/Q vssd1 vssd1 vccd1 vccd1 hold729/X sky130_fd_sc_hd__dlygate4sd3_1
X_3451_ _3735_/CLK _3451_/D vssd1 vssd1 vccd1 vccd1 _3451_/Q sky130_fd_sc_hd__dfxtp_1
X_3382_ _3419_/CLK _3382_/D vssd1 vssd1 vccd1 vccd1 _3382_/Q sky130_fd_sc_hd__dfxtp_1
X_2402_ _3194_/A0 hold399/X _2406_/S vssd1 vssd1 vccd1 vccd1 _2402_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2101__B _2480_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2902__B1 _2867_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2333_ _3194_/A0 hold415/X _2337_/S vssd1 vssd1 vccd1 vccd1 _2333_/X sky130_fd_sc_hd__mux2_1
X_2264_ _3196_/A0 hold645/X _2266_/S vssd1 vssd1 vccd1 vccd1 _2264_/X sky130_fd_sc_hd__mux2_1
X_2195_ _2479_/A _2195_/B _2479_/B _2480_/C vssd1 vssd1 vccd1 vccd1 _2640_/B sky130_fd_sc_hd__or4_4
XFILLER_0_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1979_ _1979_/A _1979_/B vssd1 vssd1 vccd1 vccd1 _3608_/D sky130_fd_sc_hd__and2_1
X_3718_ _3718_/CLK _3718_/D vssd1 vssd1 vccd1 vccd1 _3718_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3649_ _3649_/CLK _3649_/D vssd1 vssd1 vccd1 vccd1 _3649_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold12 hold12/A vssd1 vssd1 vccd1 vccd1 hold12/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 hold23/A vssd1 vssd1 vccd1 vccd1 hold23/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 hold34/A vssd1 vssd1 vccd1 vccd1 hold34/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 hold45/A vssd1 vssd1 vccd1 vccd1 hold45/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 hold56/A vssd1 vssd1 vccd1 vccd1 hold56/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 hold78/A vssd1 vssd1 vccd1 vccd1 hold78/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold89 hold89/A vssd1 vssd1 vccd1 vccd1 hold89/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 hold67/A vssd1 vssd1 vccd1 vccd1 hold67/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_85_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2681__B _2867_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2188__A1 _2355_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_452 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1699__B1 _2961_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_3_2__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_3_2__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__1794__S0 _2289_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1760__B _1760_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2112__A1 _2084_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2951_ _3103_/A _2951_/B vssd1 vssd1 vccd1 vccd1 _3625_/D sky130_fd_sc_hd__and2_1
XANTENNA__1849__S1 _1849_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_32_wb_clk_i clkbuf_3_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3447_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_1902_ _2085_/C _1902_/B vssd1 vssd1 vccd1 vccd1 _1902_/Y sky130_fd_sc_hd__nand2_1
X_2882_ hold997/X _2881_/X _2876_/A vssd1 vssd1 vccd1 vccd1 _2882_/Y sky130_fd_sc_hd__a21oi_1
X_1833_ _3468_/Q _3486_/Q _1937_/S vssd1 vssd1 vccd1 vccd1 _1834_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_25_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1764_ input4/X _1920_/B _1677_/X vssd1 vssd1 vccd1 vccd1 _1764_/X sky130_fd_sc_hd__a21o_1
X_3503_ _3539_/CLK _3503_/D vssd1 vssd1 vccd1 vccd1 _3503_/Q sky130_fd_sc_hd__dfxtp_1
Xhold515 _3457_/Q vssd1 vssd1 vccd1 vccd1 hold515/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold526 _2522_/X vssd1 vssd1 vccd1 vccd1 _3468_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1926__B2 _2854_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold504 _2285_/X vssd1 vssd1 vccd1 vccd1 _3300_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold548 _2573_/X vssd1 vssd1 vccd1 vccd1 _3512_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold559 _3273_/Q vssd1 vssd1 vccd1 vccd1 hold559/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1695_ _1680_/X _1694_/Y _1824_/B vssd1 vssd1 vccd1 vccd1 _1695_/Y sky130_fd_sc_hd__o21ai_1
Xhold537 _3370_/Q vssd1 vssd1 vccd1 vccd1 hold537/X sky130_fd_sc_hd__dlygate4sd3_1
X_3434_ _3665_/CLK _3434_/D vssd1 vssd1 vccd1 vccd1 _3434_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3365_ _3583_/CLK _3365_/D vssd1 vssd1 vccd1 vccd1 _3365_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2316_ _2316_/A _2316_/B vssd1 vssd1 vccd1 vccd1 _2316_/Y sky130_fd_sc_hd__nor2_1
X_3296_ _3581_/CLK _3296_/D vssd1 vssd1 vccd1 vccd1 _3296_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2258__S _2259_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1670__B _2960_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2247_ hold263/X _2648_/A0 _2252_/S vssd1 vssd1 vccd1 vccd1 _2247_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_25_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2103__A1 _2084_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2178_ _3225_/Q _3224_/Q _3226_/Q _3059_/B vssd1 vssd1 vccd1 vccd1 _2178_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_67_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2782__A _2797_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1862__B1 _2228_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput24 _3772_/X vssd1 vssd1 vccd1 vccd1 io_oeb[15] sky130_fd_sc_hd__buf_12
XANTENNA__2022__A _2022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput57 _3330_/Q vssd1 vssd1 vccd1 vccd1 io_out[25] sky130_fd_sc_hd__buf_12
Xoutput35 _3767_/X vssd1 vssd1 vccd1 vccd1 io_oeb[3] sky130_fd_sc_hd__buf_12
Xoutput46 _3292_/Q vssd1 vssd1 vccd1 vccd1 io_out[15] sky130_fd_sc_hd__buf_12
XANTENNA_fanout96_A _2245_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput68 _3691_/Q vssd1 vssd1 vccd1 vccd1 io_out[8] sky130_fd_sc_hd__buf_12
XANTENNA__1861__A _2085_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2676__B _2868_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1776__S0 _1981_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1853__B1 _2085_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3070__A2 _3048_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2289__D _2480_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2867__A _2867_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3150_ _3150_/A1 _3131_/X _3149_/X _3103_/A vssd1 vssd1 vccd1 vccd1 _3150_/X sky130_fd_sc_hd__o211a_1
X_2101_ _2245_/B _2480_/C vssd1 vssd1 vccd1 vccd1 _2244_/C sky130_fd_sc_hd__nor2_1
XANTENNA__2884__A2 _2940_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3081_ _3225_/Q _3081_/B vssd1 vssd1 vccd1 vccd1 _3158_/B sky130_fd_sc_hd__nor2_2
X_2032_ _2741_/A _2742_/B vssd1 vssd1 vccd1 vccd1 _2803_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_11_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2934_ _1712_/A _2997_/A1 hold409/X _2940_/B2 vssd1 vssd1 vccd1 vccd1 _2934_/X sky130_fd_sc_hd__a22o_1
X_2865_ _3613_/Q _2080_/C hold860/X vssd1 vssd1 vccd1 vccd1 _2865_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__1946__A _2006_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1816_ hold833/X _1922_/B _1814_/X _1815_/X vssd1 vssd1 vccd1 vccd1 _2868_/D sky130_fd_sc_hd__o22a_4
Xhold301 _3587_/Q vssd1 vssd1 vccd1 vccd1 hold301/X sky130_fd_sc_hd__dlygate4sd3_1
X_2796_ _2786_/Y _2839_/B _2811_/A vssd1 vssd1 vccd1 vccd1 _2797_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_25_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_27_wb_clk_i_A clkbuf_3_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_1747_ _2244_/A _1743_/Y _1745_/X _1746_/Y vssd1 vssd1 vccd1 vccd1 _1747_/X sky130_fd_sc_hd__a31o_1
Xhold312 _2098_/X vssd1 vssd1 vccd1 vccd1 _3210_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold334 _2460_/X vssd1 vssd1 vccd1 vccd1 _3419_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold323 _3335_/Q vssd1 vssd1 vccd1 vccd1 hold323/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold356 _2412_/X vssd1 vssd1 vccd1 vccd1 _3380_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold345 _3398_/Q vssd1 vssd1 vccd1 vccd1 hold345/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold367 _3563_/Q vssd1 vssd1 vccd1 vccd1 hold367/X sky130_fd_sc_hd__dlygate4sd3_1
X_1678_ _1678_/A _1922_/B vssd1 vssd1 vccd1 vccd1 _1679_/C sky130_fd_sc_hd__and2_1
Xhold378 _2232_/X vssd1 vssd1 vccd1 vccd1 _3263_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3417_ _3733_/CLK _3417_/D vssd1 vssd1 vccd1 vccd1 _3417_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold389 _3641_/Q vssd1 vssd1 vccd1 vccd1 hold389/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2496__B _3045_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3348_ _3666_/CLK _3348_/D vssd1 vssd1 vccd1 vccd1 _3348_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1001 _2180_/X vssd1 vssd1 vccd1 vccd1 _3227_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1012 _2171_/X vssd1 vssd1 vccd1 vccd1 _3225_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1023 _3296_/Q vssd1 vssd1 vccd1 vccd1 _2276_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1067 _3622_/Q vssd1 vssd1 vccd1 vccd1 _2929_/A sky130_fd_sc_hd__buf_1
Xhold1056 _3685_/Q vssd1 vssd1 vccd1 vccd1 _2309_/A sky130_fd_sc_hd__buf_1
Xhold1045 _3626_/Q vssd1 vssd1 vccd1 vccd1 _2717_/A sky130_fd_sc_hd__dlygate4sd3_1
X_3279_ _3721_/CLK hold66/X vssd1 vssd1 vccd1 vccd1 hold65/A sky130_fd_sc_hd__dfxtp_1
Xhold1034 _3294_/Q vssd1 vssd1 vccd1 vccd1 _2272_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1078 _3604_/Q vssd1 vssd1 vccd1 vccd1 _2986_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1835__B1 _2087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1930__S0 _1981_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold890 _3154_/X vssd1 vssd1 vccd1 vccd1 _3713_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2687__A _3595_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2650_ _2650_/A0 hold357/X _2653_/S vssd1 vssd1 vccd1 vccd1 _2650_/X sky130_fd_sc_hd__mux2_1
X_1601_ _2305_/A vssd1 vssd1 vccd1 vccd1 _3065_/A sky130_fd_sc_hd__inv_2
X_2581_ _2658_/A0 hold507/X _2583_/S vssd1 vssd1 vccd1 vccd1 _2581_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2554__A1 _2659_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3202_ hold677/X _2357_/A _3205_/S vssd1 vssd1 vccd1 vccd1 _3202_/X sky130_fd_sc_hd__mux2_1
X_3133_ _2892_/B _2886_/A _3137_/C vssd1 vssd1 vccd1 vccd1 _3133_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_89_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3064_ _3037_/C _3037_/D _2308_/C vssd1 vssd1 vccd1 vccd1 _3064_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_89_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1817__B1 _2868_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2015_ _3232_/Q _3247_/Q _2085_/B vssd1 vssd1 vccd1 vccd1 _2016_/B sky130_fd_sc_hd__mux2_1
XANTENNA__2490__A0 _2355_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2242__A0 _2652_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2917_ _2914_/A _2944_/B _2916_/X _3166_/C1 vssd1 vssd1 vccd1 vccd1 _2917_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_92_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2848_ hold925/X _2824_/X _2844_/X _2847_/X _2859_/A vssd1 vssd1 vccd1 vccd1 _2848_/X
+ sky130_fd_sc_hd__o221a_1
X_2779_ _2779_/A _2809_/B _2779_/C vssd1 vssd1 vccd1 vccd1 _2779_/X sky130_fd_sc_hd__or3_1
Xhold142 _2558_/X vssd1 vssd1 vccd1 vccd1 _3499_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold153 _3589_/Q vssd1 vssd1 vccd1 vccd1 hold153/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold120 _2552_/X vssd1 vssd1 vccd1 vccd1 _3494_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold131 _3304_/Q vssd1 vssd1 vccd1 vccd1 hold131/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold164 _2666_/X vssd1 vssd1 vccd1 vccd1 _3592_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold186 _2254_/X vssd1 vssd1 vccd1 vccd1 _3280_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold175 _3231_/Q vssd1 vssd1 vccd1 vccd1 hold175/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold197 _3340_/Q vssd1 vssd1 vccd1 vccd1 hold197/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1808__B1 _2428_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2233__A0 _2475_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2536__A1 _2655_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2224__A0 _2651_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2702_ _2736_/A _2714_/B vssd1 vssd1 vccd1 vccd1 _2704_/B sky130_fd_sc_hd__and2_1
XFILLER_0_27_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3682_ _3695_/CLK _3682_/D vssd1 vssd1 vccd1 vccd1 _3682_/Q sky130_fd_sc_hd__dfxtp_1
X_2633_ _2640_/A _2633_/B vssd1 vssd1 vccd1 vccd1 _2639_/S sky130_fd_sc_hd__or2_4
XANTENNA_clkbuf_3_2__f_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xscrapcpu_177 vssd1 vssd1 vccd1 vccd1 scrapcpu_177/HI io_out[35] sky130_fd_sc_hd__conb_1
XANTENNA__2527__A1 _2363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2564_ _2655_/A0 hold713/X _2569_/S vssd1 vssd1 vccd1 vccd1 _2564_/X sky130_fd_sc_hd__mux2_1
Xscrapcpu_166 vssd1 vssd1 vccd1 vccd1 scrapcpu_166/HI io_oeb[24] sky130_fd_sc_hd__conb_1
XFILLER_0_2_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2495_ _2495_/A _3242_/Q _3096_/B vssd1 vssd1 vccd1 vccd1 _2495_/X sky130_fd_sc_hd__and3_1
XFILLER_0_10_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3116_ _3697_/Q _3118_/A _3126_/A _3115_/X vssd1 vssd1 vccd1 vccd1 _3116_/X sky130_fd_sc_hd__a211o_1
X_3047_ _3063_/B _3040_/A _3183_/B _3063_/A vssd1 vssd1 vccd1 vccd1 _3047_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_77_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2463__A0 _3197_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2215__A0 _3195_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2766__A1 _2797_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2518__A1 _3196_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3191__A1 _2363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2206__A0 _2357_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout81 _2651_/A0 vssd1 vssd1 vccd1 vccd1 _3203_/A1 sky130_fd_sc_hd__buf_4
Xfanout70 _2883_/Y vssd1 vssd1 vccd1 vccd1 _2944_/B sky130_fd_sc_hd__buf_4
XFILLER_0_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout92 _3193_/A0 vssd1 vssd1 vccd1 vccd1 _2655_/A0 sky130_fd_sc_hd__buf_4
XFILLER_0_24_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2509__A1 _3201_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_57_wb_clk_i clkbuf_leaf_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3662_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2280_ _2480_/A _2195_/B _2087_/A _2480_/C vssd1 vssd1 vccd1 vccd1 _2647_/B sky130_fd_sc_hd__a31o_4
XFILLER_0_59_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2445__A0 _3193_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1995_ _2185_/C _1995_/B vssd1 vssd1 vccd1 vccd1 _1995_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_27_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3734_ _3737_/CLK _3734_/D vssd1 vssd1 vccd1 vccd1 _3734_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3665_ _3665_/CLK _3665_/D vssd1 vssd1 vccd1 vccd1 _3665_/Q sky130_fd_sc_hd__dfxtp_1
X_2616_ hold491/X _2359_/A _2618_/S vssd1 vssd1 vccd1 vccd1 _2616_/X sky130_fd_sc_hd__mux2_1
X_3596_ _3655_/CLK _3596_/D vssd1 vssd1 vccd1 vccd1 _3596_/Q sky130_fd_sc_hd__dfxtp_4
X_2547_ _2361_/A hold729/X _2548_/S vssd1 vssd1 vccd1 vccd1 _2547_/X sky130_fd_sc_hd__mux2_1
X_2478_ hold353/X _3198_/A0 _2478_/S vssd1 vssd1 vccd1 vccd1 _2478_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2279__A3 _2653_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2679__B _2867_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_3_1__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_5_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_88_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1780_ _3473_/Q _3491_/Q _1937_/S vssd1 vssd1 vccd1 vccd1 _1780_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_64_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold708 _2978_/X vssd1 vssd1 vccd1 vccd1 _3653_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold719 _3411_/Q vssd1 vssd1 vccd1 vccd1 hold719/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3450_ _3496_/CLK _3450_/D vssd1 vssd1 vccd1 vccd1 _3450_/Q sky130_fd_sc_hd__dfxtp_1
X_3381_ _3543_/CLK _3381_/D vssd1 vssd1 vccd1 vccd1 _3381_/Q sky130_fd_sc_hd__dfxtp_1
X_2401_ _3193_/A0 hold537/X _2406_/S vssd1 vssd1 vccd1 vccd1 _2401_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2902__B2 _1712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2332_ _3193_/A0 hold623/X _2337_/S vssd1 vssd1 vccd1 vccd1 _2332_/X sky130_fd_sc_hd__mux2_1
X_2263_ _2475_/A1 hold331/X _2266_/S vssd1 vssd1 vccd1 vccd1 _2263_/X sky130_fd_sc_hd__mux2_1
X_2194_ _2479_/B _2479_/C _2228_/A vssd1 vssd1 vccd1 vccd1 _2407_/A sky130_fd_sc_hd__and3b_4
XANTENNA__3091__B1 _3048_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1978_ _2046_/A _1977_/X _2028_/S vssd1 vssd1 vccd1 vccd1 _1979_/B sky130_fd_sc_hd__mux2_1
X_3717_ _3718_/CLK _3717_/D vssd1 vssd1 vccd1 vccd1 _3717_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3648_ _3674_/CLK _3648_/D vssd1 vssd1 vccd1 vccd1 _3648_/Q sky130_fd_sc_hd__dfxtp_1
X_3579_ _3724_/CLK _3579_/D vssd1 vssd1 vccd1 vccd1 _3579_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2354__C1 _3058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold13 hold13/A vssd1 vssd1 vccd1 vccd1 hold13/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 hold35/A vssd1 vssd1 vccd1 vccd1 hold35/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_2_wb_clk_i clkbuf_leaf_5_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3654_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold46 hold46/A vssd1 vssd1 vccd1 vccd1 hold46/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 hold24/A vssd1 vssd1 vccd1 vccd1 hold24/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2657__A0 _3195_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold57 hold57/A vssd1 vssd1 vccd1 vccd1 hold57/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 hold79/A vssd1 vssd1 vccd1 vccd1 hold79/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold68 hold68/A vssd1 vssd1 vccd1 vccd1 hold68/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2409__A0 _2656_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1859__A _2014_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1794__S1 _2479_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2648__A0 _2648_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2112__A2 _2084_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2950_ _2948_/A _2944_/Y _2949_/X _2944_/B vssd1 vssd1 vccd1 vccd1 _2951_/B sky130_fd_sc_hd__a22o_1
XANTENNA__3073__B1 _3157_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2881_ _3613_/Q _2712_/A _3627_/Q _1672_/B _1711_/X vssd1 vssd1 vccd1 vccd1 _2881_/X
+ sky130_fd_sc_hd__o311a_1
X_1901_ hold37/A _3299_/Q _2005_/S vssd1 vssd1 vccd1 vccd1 _1902_/B sky130_fd_sc_hd__mux2_1
X_1832_ _2085_/C _1832_/B vssd1 vssd1 vccd1 vccd1 _1832_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_25_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_17_wb_clk_i_A clkbuf_3_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_1763_ input10/X _2022_/A _1759_/Y _1762_/X vssd1 vssd1 vccd1 vccd1 _1763_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_52_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3502_ _3744_/CLK _3502_/D vssd1 vssd1 vccd1 vccd1 _3502_/Q sky130_fd_sc_hd__dfxtp_1
Xhold516 _2509_/X vssd1 vssd1 vccd1 vccd1 _3457_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold505 _3542_/Q vssd1 vssd1 vccd1 vccd1 hold505/X sky130_fd_sc_hd__dlygate4sd3_1
X_1694_ _2876_/A _1694_/B vssd1 vssd1 vccd1 vccd1 _1694_/Y sky130_fd_sc_hd__nor2_1
Xhold527 _3736_/Q vssd1 vssd1 vccd1 vccd1 hold527/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold538 _2401_/X vssd1 vssd1 vccd1 vccd1 _3370_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3433_ _3665_/CLK _3433_/D vssd1 vssd1 vccd1 vccd1 _3433_/Q sky130_fd_sc_hd__dfxtp_1
Xhold549 _3410_/Q vssd1 vssd1 vccd1 vccd1 hold549/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3364_ _3570_/CLK _3364_/D vssd1 vssd1 vccd1 vccd1 _3364_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2315_ _2315_/A _2316_/B vssd1 vssd1 vccd1 vccd1 _3089_/B sky130_fd_sc_hd__nor2_1
X_3295_ _3725_/CLK _3295_/D vssd1 vssd1 vccd1 vccd1 _3295_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2639__A0 _2660_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2246_ _2290_/A _3199_/A vssd1 vssd1 vccd1 vccd1 _2252_/S sky130_fd_sc_hd__nor2_2
XFILLER_0_79_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2103__A2 _2084_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2177_ _2182_/B vssd1 vssd1 vccd1 vccd1 _2177_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_79_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1862__A1 _2289_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_56_wb_clk_i_A clkbuf_leaf_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_75_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput25 _3772_/A vssd1 vssd1 vccd1 vccd1 io_oeb[16] sky130_fd_sc_hd__buf_12
Xoutput58 _3331_/Q vssd1 vssd1 vccd1 vccd1 io_out[26] sky130_fd_sc_hd__buf_12
Xoutput36 _1705_/X vssd1 vssd1 vccd1 vccd1 io_oeb[4] sky130_fd_sc_hd__buf_12
Xoutput47 _3293_/Q vssd1 vssd1 vccd1 vccd1 io_out[16] sky130_fd_sc_hd__buf_12
XANTENNA_fanout89_A _2091_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput69 _3400_/Q vssd1 vssd1 vccd1 vccd1 io_out[9] sky130_fd_sc_hd__buf_12
XANTENNA__1776__S1 _1981_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2692__B _2867_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1853__A1 _3769_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2867__B _2867_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3080_ _3080_/A _3080_/B _3080_/C vssd1 vssd1 vccd1 vccd1 _3085_/S sky130_fd_sc_hd__and3_1
X_2100_ hold25/X _2653_/A0 _2100_/S vssd1 vssd1 vccd1 vccd1 hold26/A sky130_fd_sc_hd__mux2_1
X_2031_ _2050_/B vssd1 vssd1 vccd1 vccd1 _2031_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_76_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3046__B1 _3108_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2933_ _3103_/A _2933_/B vssd1 vssd1 vccd1 vccd1 _3622_/D sky130_fd_sc_hd__and2_1
XFILLER_0_57_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2864_ _3594_/Q _2861_/X _2080_/C vssd1 vssd1 vccd1 vccd1 _2864_/X sky130_fd_sc_hd__o21a_1
X_2795_ _2790_/X _2791_/Y _2794_/X vssd1 vssd1 vccd1 vccd1 _2839_/B sky130_fd_sc_hd__a21oi_2
X_1815_ input5/X _1920_/B _1677_/X vssd1 vssd1 vccd1 vccd1 _1815_/X sky130_fd_sc_hd__a21o_1
Xhold302 _2660_/X vssd1 vssd1 vccd1 vccd1 _3587_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1746_ _2244_/A _1741_/X _2087_/A vssd1 vssd1 vccd1 vccd1 _1746_/Y sky130_fd_sc_hd__o21ai_1
Xhold313 _3645_/Q vssd1 vssd1 vccd1 vccd1 hold313/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold335 _3661_/Q vssd1 vssd1 vccd1 vccd1 hold335/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold324 _2367_/X vssd1 vssd1 vccd1 vccd1 _3335_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold346 _2435_/X vssd1 vssd1 vccd1 vccd1 _3398_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold368 _2632_/X vssd1 vssd1 vccd1 vccd1 _3563_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1677_ _1677_/A _1677_/B _1683_/B vssd1 vssd1 vccd1 vccd1 _1677_/X sky130_fd_sc_hd__or3b_2
XFILLER_0_40_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold357 _3578_/Q vssd1 vssd1 vccd1 vccd1 hold357/X sky130_fd_sc_hd__dlygate4sd3_1
X_3416_ _3733_/CLK hold36/X vssd1 vssd1 vccd1 vccd1 hold35/A sky130_fd_sc_hd__dfxtp_1
Xhold379 _3222_/Q vssd1 vssd1 vccd1 vccd1 hold379/X sky130_fd_sc_hd__dlygate4sd3_1
X_3347_ _3668_/CLK _3347_/D vssd1 vssd1 vccd1 vccd1 _3347_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1013 _3693_/Q vssd1 vssd1 vccd1 vccd1 _1599_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1002 _3711_/Q vssd1 vssd1 vccd1 vccd1 _3150_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1024 _2277_/X vssd1 vssd1 vccd1 vccd1 _3296_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1057 _3049_/X vssd1 vssd1 vccd1 vccd1 _3685_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1046 _3681_/Q vssd1 vssd1 vccd1 vccd1 _3035_/A sky130_fd_sc_hd__buf_1
X_3278_ _3308_/CLK hold2/X vssd1 vssd1 vccd1 vccd1 hold1/A sky130_fd_sc_hd__dfxtp_1
Xhold1035 _3297_/Q vssd1 vssd1 vccd1 vccd1 _2278_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1068 _2932_/X vssd1 vssd1 vccd1 vccd1 _2933_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1079 _3619_/Q vssd1 vssd1 vccd1 vccd1 _2967_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_2229_ _2289_/A _1954_/S _2014_/A _2480_/C vssd1 vssd1 vccd1 vccd1 _2598_/A sky130_fd_sc_hd__a31o_4
XANTENNA__1835__A1 _1889_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1930__S1 _1981_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1771__A0 _2074_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold891 _3323_/Q vssd1 vssd1 vccd1 vccd1 hold891/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold880 _3324_/Q vssd1 vssd1 vccd1 vccd1 hold880/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2251__A1 _2652_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1600_ _1600_/A vssd1 vssd1 vccd1 vccd1 _1600_/Y sky130_fd_sc_hd__inv_2
X_2580_ _3195_/A0 hold361/X _2583_/S vssd1 vssd1 vccd1 vccd1 _2580_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_22_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3201_ hold125/X _3201_/A1 _3205_/S vssd1 vssd1 vccd1 vccd1 _3201_/X sky130_fd_sc_hd__mux2_1
X_3132_ hold992/X _3130_/Y _2877_/X vssd1 vssd1 vccd1 vccd1 _3137_/C sky130_fd_sc_hd__o21ai_4
X_3063_ _3063_/A _3063_/B _3682_/Q vssd1 vssd1 vccd1 vccd1 _3063_/X sky130_fd_sc_hd__or3b_1
X_2014_ _2014_/A _2014_/B vssd1 vssd1 vccd1 vccd1 _2014_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_77_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2916_ _2885_/B _2912_/X _2915_/X vssd1 vssd1 vccd1 vccd1 _2916_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_57_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2847_ _2797_/A _2845_/X _2846_/X _2825_/Y vssd1 vssd1 vccd1 vccd1 _2847_/X sky130_fd_sc_hd__a31o_1
XANTENNA_fanout139_A _3346_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold110 _2560_/X vssd1 vssd1 vccd1 vccd1 _3501_/D sky130_fd_sc_hd__dlygate4sd3_1
X_2778_ _2707_/B _2707_/C _2762_/A vssd1 vssd1 vccd1 vccd1 _2779_/C sky130_fd_sc_hd__a21oi_1
X_1729_ hold81/A _3478_/Q hold35/A _3428_/Q _2244_/B _2185_/C vssd1 vssd1 vccd1 vccd1
+ _1730_/B sky130_fd_sc_hd__mux4_1
Xhold121 _3459_/Q vssd1 vssd1 vccd1 vccd1 hold121/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold143 _3388_/Q vssd1 vssd1 vccd1 vccd1 hold143/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold132 _2291_/X vssd1 vssd1 vccd1 vccd1 _3304_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold154 _2663_/X vssd1 vssd1 vccd1 vccd1 _3589_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold165 _3207_/Q vssd1 vssd1 vccd1 vccd1 hold165/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold176 _2189_/X vssd1 vssd1 vccd1 vccd1 _3231_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold198 _2373_/X vssd1 vssd1 vccd1 vccd1 _3340_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold187 _3737_/Q vssd1 vssd1 vccd1 vccd1 hold187/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1808__A1 _3348_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1867__A _2022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1806__S _1937_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2210__B _2479_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2701_ _3594_/Q _2701_/B vssd1 vssd1 vccd1 vccd1 _2714_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_40_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3681_ _3725_/CLK _3681_/D vssd1 vssd1 vccd1 vccd1 _3681_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2632_ hold367/X _3198_/A0 _2632_/S vssd1 vssd1 vccd1 vccd1 _2632_/X sky130_fd_sc_hd__mux2_1
X_2563_ _2654_/A _2598_/A vssd1 vssd1 vccd1 vccd1 _2569_/S sky130_fd_sc_hd__nand2_4
Xscrapcpu_167 vssd1 vssd1 vccd1 vccd1 scrapcpu_167/HI io_oeb[25] sky130_fd_sc_hd__conb_1
Xscrapcpu_178 vssd1 vssd1 vccd1 vccd1 io_oeb[29] scrapcpu_178/LO sky130_fd_sc_hd__conb_1
XANTENNA__1735__B1 _2428_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1830__S0 _1937_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2494_ _2653_/A0 hold687/X _2494_/S vssd1 vssd1 vccd1 vccd1 _2494_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_65_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3115_ _3010_/Y _3118_/B _3183_/B vssd1 vssd1 vccd1 vccd1 _3115_/X sky130_fd_sc_hd__o21a_1
XANTENNA__2160__B1 _3157_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3046_ hold946/X _3045_/X _3108_/A vssd1 vssd1 vccd1 vccd1 _3046_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__1897__S0 _2000_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3176__C1 _3058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_3_0__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_1_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_41_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2030__B _3045_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout71_A _3198_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2454__A1 _2650_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout71 _3198_/A0 vssd1 vssd1 vccd1 vccd1 _2660_/A0 sky130_fd_sc_hd__buf_4
Xfanout82 _2359_/A vssd1 vssd1 vccd1 vccd1 _2651_/A0 sky130_fd_sc_hd__buf_4
XFILLER_0_64_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout93 _2089_/X vssd1 vssd1 vccd1 vccd1 _3193_/A0 sky130_fd_sc_hd__buf_4
XFILLER_0_36_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2390__A0 _3196_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_26_wb_clk_i clkbuf_3_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3744_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_59_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1879__S0 _1981_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1994_ hold43/A _3397_/Q _1996_/S vssd1 vssd1 vccd1 vccd1 _1995_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_55_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3733_ _3733_/CLK hold60/X vssd1 vssd1 vccd1 vccd1 hold59/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3664_ _3668_/CLK _3664_/D vssd1 vssd1 vccd1 vccd1 _3664_/Q sky130_fd_sc_hd__dfxtp_1
X_2615_ hold107/X _2643_/A1 _2618_/S vssd1 vssd1 vccd1 vccd1 _2615_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_70_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3595_ _3662_/CLK _3595_/D vssd1 vssd1 vccd1 vccd1 _3595_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_23_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2546_ _3203_/A1 hold439/X _2548_/S vssd1 vssd1 vccd1 vccd1 _2546_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2381__A0 _2656_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2477_ hold471/X _3197_/A0 _2478_/S vssd1 vssd1 vccd1 vccd1 _2477_/X sky130_fd_sc_hd__mux2_1
XANTENNA_hold1021_A _3351_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2436__A1 _2363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3029_ _3678_/Q _3677_/Q _3080_/A _3030_/A vssd1 vssd1 vccd1 vccd1 _3029_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_73_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1947__B1 _2428_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2427__A1 _2660_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold709 _3379_/Q vssd1 vssd1 vccd1 vccd1 hold709/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2400_ _3192_/A _3199_/A vssd1 vssd1 vccd1 vccd1 _2406_/S sky130_fd_sc_hd__or2_4
X_3380_ _3543_/CLK _3380_/D vssd1 vssd1 vccd1 vccd1 _3380_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2902__A2 _2940_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2331_ _2365_/A _2647_/A vssd1 vssd1 vccd1 vccd1 _2337_/S sky130_fd_sc_hd__nand2_2
X_2262_ _3194_/A0 hold679/X _2266_/S vssd1 vssd1 vccd1 vccd1 _2262_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2115__A0 _2355_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2666__A1 _2361_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2193_ _2195_/B _2480_/C vssd1 vssd1 vccd1 vccd1 _2479_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_79_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2418__A1 _3196_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_46_wb_clk_i_A clkbuf_3_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__1965__A _2085_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1977_ _2996_/A1 _1769_/Y _1976_/X _2854_/B vssd1 vssd1 vccd1 vccd1 _1977_/X sky130_fd_sc_hd__o22a_1
X_3716_ _3718_/CLK _3716_/D vssd1 vssd1 vccd1 vccd1 _3716_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2051__C1 _2495_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout121_A _3349_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3647_ _3674_/CLK _3647_/D vssd1 vssd1 vccd1 vccd1 _3647_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3578_ _3581_/CLK _3578_/D vssd1 vssd1 vccd1 vccd1 _3578_/Q sky130_fd_sc_hd__dfxtp_1
X_2529_ hold17/X _2353_/A _2534_/S vssd1 vssd1 vccd1 vccd1 hold18/A sky130_fd_sc_hd__mux2_1
Xhold14 hold14/A vssd1 vssd1 vccd1 vccd1 hold14/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 hold36/A vssd1 vssd1 vccd1 vccd1 hold36/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 hold47/A vssd1 vssd1 vccd1 vccd1 hold47/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 hold25/A vssd1 vssd1 vccd1 vccd1 hold25/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2106__A0 _3193_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold69 hold69/A vssd1 vssd1 vccd1 vccd1 hold69/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 hold58/A vssd1 vssd1 vccd1 vccd1 hold58/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1875__A _1979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2345__A0 _2651_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2880_ hold996/X _3630_/Q _2741_/B _2879_/Y vssd1 vssd1 vccd1 vccd1 _2880_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_29_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1900_ _3293_/Q _3443_/Q _3577_/Q _3401_/Q _1954_/S _2014_/A vssd1 vssd1 vccd1 vccd1
+ _1900_/X sky130_fd_sc_hd__mux4_1
X_1831_ _3436_/Q _3740_/Q _1937_/S vssd1 vssd1 vccd1 vccd1 _1832_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_32_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1762_ _2087_/B _1762_/B _1762_/C vssd1 vssd1 vccd1 vccd1 _1762_/X sky130_fd_sc_hd__or3_4
XFILLER_0_52_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3501_ _3741_/CLK _3501_/D vssd1 vssd1 vccd1 vccd1 _3501_/Q sky130_fd_sc_hd__dfxtp_1
Xhold506 _2608_/X vssd1 vssd1 vccd1 vccd1 _3542_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1693_ _2080_/A _2960_/A _1692_/X _1979_/A vssd1 vssd1 vccd1 vccd1 _1693_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_40_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold517 _3262_/Q vssd1 vssd1 vccd1 vccd1 hold517/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold539 _3238_/Q vssd1 vssd1 vccd1 vccd1 hold539/X sky130_fd_sc_hd__dlygate4sd3_1
X_3432_ _3496_/CLK _3432_/D vssd1 vssd1 vccd1 vccd1 _3432_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2336__A0 _3197_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold528 _3195_/X vssd1 vssd1 vccd1 vccd1 _3736_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_41_wb_clk_i clkbuf_3_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3725_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_3363_ _3387_/CLK _3363_/D vssd1 vssd1 vccd1 vccd1 _3363_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2887__A1 _2876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2314_ hold858/X _2316_/A _3089_/A _3059_/B vssd1 vssd1 vccd1 vccd1 _2314_/X sky130_fd_sc_hd__o211a_1
X_3294_ _3581_/CLK _3294_/D vssd1 vssd1 vccd1 vccd1 _3294_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2245_ _2289_/A _2245_/B _2245_/C _1937_/S vssd1 vssd1 vccd1 vccd1 _3199_/A sky130_fd_sc_hd__or4b_4
X_2176_ _3225_/Q _3224_/Q _3059_/B _3226_/Q vssd1 vssd1 vccd1 vccd1 _2182_/B sky130_fd_sc_hd__and4_1
XFILLER_0_79_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_2_wb_clk_i_A clkbuf_leaf_5_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__3049__D1 _3055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2575__A0 _2361_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput26 _3773_/X vssd1 vssd1 vccd1 vccd1 io_oeb[17] sky130_fd_sc_hd__buf_12
Xoutput37 _3768_/X vssd1 vssd1 vccd1 vccd1 io_oeb[5] sky130_fd_sc_hd__buf_12
Xoutput48 _3294_/Q vssd1 vssd1 vccd1 vccd1 io_out[17] sky130_fd_sc_hd__buf_12
Xoutput59 _3332_/Q vssd1 vssd1 vccd1 vccd1 io_out[27] sky130_fd_sc_hd__buf_12
XFILLER_0_85_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2566__A0 _3195_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2867__C _2867_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2869__A1 _2701_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2030_ _2071_/A _3045_/B _2042_/D vssd1 vssd1 vccd1 vccd1 _2050_/B sky130_fd_sc_hd__or3_2
XANTENNA__2097__A2 _2084_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2932_ _2944_/B _2930_/X _2931_/Y _2929_/A vssd1 vssd1 vccd1 vccd1 _2932_/X sky130_fd_sc_hd__a22o_1
X_2863_ _2863_/A _2863_/B _2863_/C vssd1 vssd1 vccd1 vccd1 _2863_/X sky130_fd_sc_hd__and3_1
XFILLER_0_57_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1814_ input11/X _2022_/A _1762_/X _1813_/Y vssd1 vssd1 vccd1 vccd1 _1814_/X sky130_fd_sc_hd__o211a_1
X_2794_ _2723_/Y _2788_/Y _2793_/X _2708_/Y _2792_/X vssd1 vssd1 vccd1 vccd1 _2794_/X
+ sky130_fd_sc_hd__a221o_1
X_1745_ _3773_/A _2005_/S _2085_/C _1744_/Y vssd1 vssd1 vccd1 vccd1 _1745_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_40_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold325 _3473_/Q vssd1 vssd1 vccd1 vccd1 hold325/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold303 _3585_/Q vssd1 vssd1 vccd1 vccd1 hold303/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold314 _2970_/X vssd1 vssd1 vccd1 vccd1 _3645_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold369 _3583_/Q vssd1 vssd1 vccd1 vccd1 hold369/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold347 _3395_/Q vssd1 vssd1 vccd1 vccd1 hold347/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold336 _2986_/X vssd1 vssd1 vccd1 vccd1 _3661_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1676_ _1677_/A _1676_/B _1683_/B vssd1 vssd1 vccd1 vccd1 _1922_/B sky130_fd_sc_hd__and3b_4
XFILLER_0_40_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold358 _2650_/X vssd1 vssd1 vccd1 vccd1 _3578_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3415_ _3732_/CLK _3415_/D vssd1 vssd1 vccd1 vccd1 _3415_/Q sky130_fd_sc_hd__dfxtp_1
X_3346_ _3666_/CLK _3346_/D vssd1 vssd1 vccd1 vccd1 _3346_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1014 _3100_/X vssd1 vssd1 vccd1 vccd1 _3101_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1003 _3150_/X vssd1 vssd1 vccd1 vccd1 _3711_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1036 _2279_/X vssd1 vssd1 vccd1 vccd1 _3297_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1058 _3623_/Q vssd1 vssd1 vccd1 vccd1 _2941_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1025 _3691_/Q vssd1 vssd1 vccd1 vccd1 _3085_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1047 _3036_/X vssd1 vssd1 vccd1 vccd1 _3681_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3277_ _3721_/CLK hold22/X vssd1 vssd1 vccd1 vccd1 hold21/A sky130_fd_sc_hd__dfxtp_1
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1069 _3606_/Q vssd1 vssd1 vccd1 vccd1 _2994_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_2228_ _2228_/A _2228_/B _2228_/C _2480_/C vssd1 vssd1 vccd1 vccd1 _2549_/A sky130_fd_sc_hd__or4_4
X_2159_ _1679_/C _2159_/B _2819_/A _2159_/D vssd1 vssd1 vccd1 vccd1 _2159_/X sky130_fd_sc_hd__and4b_1
XFILLER_0_67_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2548__A0 _2363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold881 _3403_/Q vssd1 vssd1 vccd1 vccd1 hold881/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold870 _3169_/X vssd1 vssd1 vccd1 vccd1 hold870/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold892 _2341_/X vssd1 vssd1 vccd1 vccd1 _2342_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3200__A1 _2353_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3200_ hold269/X _2353_/A _3205_/S vssd1 vssd1 vccd1 vccd1 _3200_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3055__A _3055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3131_ hold992/X _3130_/Y _2877_/X vssd1 vssd1 vccd1 vccd1 _3131_/X sky130_fd_sc_hd__o21a_4
XFILLER_0_89_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3062_ _2167_/C _3061_/X _2298_/A vssd1 vssd1 vccd1 vccd1 _3062_/X sky130_fd_sc_hd__o21a_1
XANTENNA__1817__A2 _2731_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2013_ _3259_/Q _3271_/Q _2085_/B vssd1 vssd1 vccd1 vccd1 _2014_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_49_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2915_ _2948_/B _2913_/Y _2924_/C _2944_/B vssd1 vssd1 vccd1 vccd1 _2915_/X sky130_fd_sc_hd__o31a_1
XFILLER_0_45_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2846_ hold79/X _2846_/B vssd1 vssd1 vccd1 vccd1 _2846_/X sky130_fd_sc_hd__or2_1
XFILLER_0_5_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold100 _3189_/X vssd1 vssd1 vccd1 vccd1 _3731_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2777_ _2723_/Y _2773_/B _2776_/X vssd1 vssd1 vccd1 vccd1 _2777_/Y sky130_fd_sc_hd__a21oi_1
X_1728_ _1889_/A _1724_/Y _1726_/Y _1727_/Y vssd1 vssd1 vccd1 vccd1 _1728_/X sky130_fd_sc_hd__a31o_1
Xhold111 _3529_/Q vssd1 vssd1 vccd1 vccd1 hold111/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold122 _2511_/X vssd1 vssd1 vccd1 vccd1 _3459_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold144 _2422_/X vssd1 vssd1 vccd1 vccd1 _3388_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold133 _3342_/Q vssd1 vssd1 vccd1 vccd1 hold133/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold155 _3547_/Q vssd1 vssd1 vccd1 vccd1 hold155/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold177 _3260_/Q vssd1 vssd1 vccd1 vccd1 hold177/X sky130_fd_sc_hd__dlygate4sd3_1
X_1659_ _1663_/B _1659_/B _1672_/B vssd1 vssd1 vccd1 vccd1 _1678_/A sky130_fd_sc_hd__or3_1
Xhold166 _2092_/X vssd1 vssd1 vccd1 vccd1 _3207_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold199 _3643_/Q vssd1 vssd1 vccd1 vccd1 hold199/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold188 _3196_/X vssd1 vssd1 vccd1 vccd1 _3737_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3329_ _3728_/CLK _3329_/D vssd1 vssd1 vccd1 vccd1 _3329_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1883__A _2006_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2700_ _2788_/A _2700_/B vssd1 vssd1 vccd1 vccd1 _2709_/C sky130_fd_sc_hd__xor2_2
X_3680_ _3725_/CLK _3680_/D vssd1 vssd1 vccd1 vccd1 _3680_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2631_ hold209/X _2659_/A0 _2632_/S vssd1 vssd1 vccd1 vccd1 _2631_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_35_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2562_ hold425/X _2363_/A _2562_/S vssd1 vssd1 vccd1 vccd1 _2562_/X sky130_fd_sc_hd__mux2_1
Xscrapcpu_168 vssd1 vssd1 vccd1 vccd1 scrapcpu_168/HI io_oeb[26] sky130_fd_sc_hd__conb_1
XANTENNA__1735__A1 _1889_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1830__S1 _2245_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2493_ _2652_/A0 hold329/X _2494_/S vssd1 vssd1 vccd1 vccd1 _2493_/X sky130_fd_sc_hd__mux2_1
X_3114_ hold825/X _3120_/A _3113_/X _3055_/A vssd1 vssd1 vccd1 vccd1 _3114_/X sky130_fd_sc_hd__o211a_1
X_3045_ _3045_/A _3045_/B _3096_/A _3045_/D vssd1 vssd1 vccd1 vccd1 _3045_/X sky130_fd_sc_hd__or4_1
XANTENNA__1897__S1 _2219_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout151_A input18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2829_ hold923/X _1696_/Y _2940_/B2 hold647/X _2825_/Y vssd1 vssd1 vccd1 vccd1 _2829_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_5_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1888__S1 _2185_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout72 _2099_/X vssd1 vssd1 vccd1 vccd1 _3198_/A0 sky130_fd_sc_hd__buf_4
Xfanout83 _2475_/A1 vssd1 vssd1 vccd1 vccd1 _3195_/A0 sky130_fd_sc_hd__buf_4
Xfanout94 _2089_/X vssd1 vssd1 vccd1 vccd1 _2648_/A0 sky130_fd_sc_hd__buf_4
XFILLER_0_91_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1879__S1 _1981_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_36_wb_clk_i_A clkbuf_3_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_59_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1993_ _2185_/A _1993_/B vssd1 vssd1 vccd1 vccd1 _1993_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_27_132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3732_ _3732_/CLK hold82/X vssd1 vssd1 vccd1 vccd1 hold81/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3663_ _3666_/CLK _3663_/D vssd1 vssd1 vccd1 vccd1 _3663_/Q sky130_fd_sc_hd__dfxtp_1
X_2614_ hold155/X _2656_/A0 _2618_/S vssd1 vssd1 vccd1 vccd1 _2614_/X sky130_fd_sc_hd__mux2_1
X_3594_ _3662_/CLK _3594_/D vssd1 vssd1 vccd1 vccd1 _3594_/Q sky130_fd_sc_hd__dfxtp_2
X_2545_ _2357_/A hold651/X _2548_/S vssd1 vssd1 vccd1 vccd1 _2545_/X sky130_fd_sc_hd__mux2_1
X_2476_ hold139/X _3196_/A0 _2478_/S vssd1 vssd1 vccd1 vccd1 _2476_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_76_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3028_ _3086_/A _3036_/B _3028_/C vssd1 vssd1 vccd1 vccd1 _3028_/X sky130_fd_sc_hd__and3_1
XFILLER_0_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2330_ hold842/X _2318_/B _2329_/X _3108_/A vssd1 vssd1 vccd1 vccd1 _2330_/X sky130_fd_sc_hd__a211o_1
X_2261_ _3193_/A0 hold755/X _2266_/S vssd1 vssd1 vccd1 vccd1 _2261_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_46_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2192_ hold3/X _2653_/A0 _2192_/S vssd1 vssd1 vccd1 vccd1 hold4/A sky130_fd_sc_hd__mux2_1
XANTENNA__1874__A0 _2074_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1721__S0 _2085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1976_ hold385/X _2731_/A2 _2867_/B _1713_/X vssd1 vssd1 vccd1 vccd1 _1976_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_55_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3715_ _3723_/CLK _3715_/D vssd1 vssd1 vccd1 vccd1 _3715_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3646_ _3646_/CLK _3646_/D vssd1 vssd1 vccd1 vccd1 _3646_/Q sky130_fd_sc_hd__dfxtp_1
X_3577_ _3724_/CLK _3577_/D vssd1 vssd1 vccd1 vccd1 _3577_/Q sky130_fd_sc_hd__dfxtp_1
X_2528_ _2570_/A _2528_/B vssd1 vssd1 vccd1 vccd1 _2534_/S sky130_fd_sc_hd__and2_2
XFILLER_0_11_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold15 hold15/A vssd1 vssd1 vccd1 vccd1 hold15/X sky130_fd_sc_hd__dlygate4sd3_1
X_2459_ _3193_/A0 hold281/X _2464_/S vssd1 vssd1 vccd1 vccd1 _2459_/X sky130_fd_sc_hd__mux2_1
Xhold26 hold26/A vssd1 vssd1 vccd1 vccd1 hold26/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 hold37/A vssd1 vssd1 vccd1 vccd1 hold37/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 hold59/A vssd1 vssd1 vccd1 vccd1 hold59/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold48 hold48/A vssd1 vssd1 vccd1 vccd1 hold48/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1865__B1 _2195_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1960__S0 _2085_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2593__A1 _3201_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1891__A _2185_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1830_ _3498_/Q _3510_/Q _3522_/Q _3534_/Q _1937_/S _2245_/B vssd1 vssd1 vccd1 vccd1
+ _1830_/X sky130_fd_sc_hd__mux4_1
X_3500_ _3539_/CLK _3500_/D vssd1 vssd1 vccd1 vccd1 _3500_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3058__A _3058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1761_ _2087_/B _1762_/B _1762_/C vssd1 vssd1 vccd1 vccd1 _1920_/B sky130_fd_sc_hd__nor3_4
Xhold507 _3519_/Q vssd1 vssd1 vccd1 vccd1 hold507/X sky130_fd_sc_hd__dlygate4sd3_1
X_1692_ _1683_/B _1694_/B _1685_/B vssd1 vssd1 vccd1 vccd1 _1692_/X sky130_fd_sc_hd__a21o_1
Xhold518 _2231_/X vssd1 vssd1 vccd1 vccd1 _3262_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold529 _3467_/Q vssd1 vssd1 vccd1 vccd1 hold529/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3431_ _3665_/CLK _3431_/D vssd1 vssd1 vccd1 vccd1 _3431_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3362_ _3654_/CLK _3362_/D vssd1 vssd1 vccd1 vccd1 _3362_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2887__A2 _1696_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2313_ _3227_/Q _2315_/A _3089_/A vssd1 vssd1 vccd1 vccd1 _2313_/X sky130_fd_sc_hd__and3_1
XFILLER_0_57_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3293_ _3724_/CLK _3293_/D vssd1 vssd1 vccd1 vccd1 _3293_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2244_ _2244_/A _2244_/B _2244_/C vssd1 vssd1 vccd1 vccd1 _2654_/B sky130_fd_sc_hd__and3_2
X_2175_ _3157_/B _2174_/Y _2175_/B1 _3108_/A vssd1 vssd1 vccd1 vccd1 _2175_/Y sky130_fd_sc_hd__a211oi_1
Xclkbuf_leaf_10_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3738_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_7_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1959_ _2244_/A _1955_/Y _1957_/X _1958_/Y vssd1 vssd1 vccd1 vccd1 _1959_/X sky130_fd_sc_hd__a31o_1
XANTENNA__1783__C1 _2087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3629_ _3668_/CLK _3629_/D vssd1 vssd1 vccd1 vccd1 _3629_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput38 _3768_/A vssd1 vssd1 vccd1 vccd1 io_oeb[6] sky130_fd_sc_hd__buf_12
Xoutput27 _3773_/A vssd1 vssd1 vccd1 vccd1 io_oeb[18] sky130_fd_sc_hd__buf_12
Xoutput49 _3295_/Q vssd1 vssd1 vccd1 vccd1 io_out[18] sky130_fd_sc_hd__buf_12
XANTENNA__1933__S0 _2085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2263__A0 _2475_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2931_ _2948_/B _2935_/B _2944_/B vssd1 vssd1 vccd1 vccd1 _2931_/Y sky130_fd_sc_hd__o21ai_1
X_2862_ _1627_/Y _2846_/B _2845_/X _2861_/X _2797_/A vssd1 vssd1 vccd1 vccd1 _2862_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA__2557__A1 _2353_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1813_ _1809_/X _1810_/Y _1812_/X _2022_/A vssd1 vssd1 vccd1 vccd1 _1813_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_0_4_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2793_ _2709_/C _2779_/A _2809_/B vssd1 vssd1 vccd1 vccd1 _2793_/X sky130_fd_sc_hd__o21ba_1
X_1744_ _3332_/Q _2244_/B vssd1 vssd1 vccd1 vccd1 _1744_/Y sky130_fd_sc_hd__nor2_1
Xhold326 _2527_/X vssd1 vssd1 vccd1 vccd1 _3473_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold304 _2658_/X vssd1 vssd1 vccd1 vccd1 _3585_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold315 _3415_/Q vssd1 vssd1 vccd1 vccd1 hold315/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold348 _2432_/X vssd1 vssd1 vccd1 vccd1 _3395_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3414_ _3592_/CLK hold6/X vssd1 vssd1 vccd1 vccd1 hold5/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1675_ _1653_/C _1713_/B _1662_/B vssd1 vssd1 vccd1 vccd1 _1683_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_40_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold337 _3577_/Q vssd1 vssd1 vccd1 vccd1 hold337/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold359 _3213_/Q vssd1 vssd1 vccd1 vccd1 hold359/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3345_ _3728_/CLK hold58/X vssd1 vssd1 vccd1 vccd1 hold57/A sky130_fd_sc_hd__dfxtp_1
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1015 _3712_/Q vssd1 vssd1 vccd1 vccd1 _3152_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1004 _3224_/Q vssd1 vssd1 vccd1 vccd1 _3059_/A sky130_fd_sc_hd__buf_2
X_3276_ _3676_/CLK hold46/X vssd1 vssd1 vccd1 vccd1 hold45/A sky130_fd_sc_hd__dfxtp_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1048 _3627_/Q vssd1 vssd1 vccd1 vccd1 _2058_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1026 _3085_/X vssd1 vssd1 vccd1 vccd1 _3086_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1037 _3293_/Q vssd1 vssd1 vccd1 vccd1 _2270_/A sky130_fd_sc_hd__dlygate4sd3_1
X_2227_ _2228_/A _2228_/B _2228_/C _2480_/C vssd1 vssd1 vccd1 vccd1 _2500_/B sky130_fd_sc_hd__nor4_4
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1059 _2941_/X vssd1 vssd1 vccd1 vccd1 _2949_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2493__A0 _2652_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2158_ _3096_/A _3096_/B vssd1 vssd1 vccd1 vccd1 _2167_/C sky130_fd_sc_hd__nand2_2
X_2089_ hold908/X _2084_/A _2099_/B1 hold978/X vssd1 vssd1 vccd1 vccd1 _2089_/X sky130_fd_sc_hd__a22o_4
XFILLER_0_48_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold860 _3632_/Q vssd1 vssd1 vccd1 vccd1 hold860/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout94_A _2089_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold882 _2441_/X vssd1 vssd1 vccd1 vccd1 _3403_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold871 _3170_/X vssd1 vssd1 vccd1 vccd1 _3720_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold893 _3597_/Q vssd1 vssd1 vccd1 vccd1 hold893/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_58_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2236__A0 _3198_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2539__A1 _2658_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3130_ _3130_/A _3130_/B vssd1 vssd1 vccd1 vccd1 _3130_/Y sky130_fd_sc_hd__nor2_2
X_3061_ _2153_/Y _3060_/Y _2166_/X vssd1 vssd1 vccd1 vccd1 _3061_/X sky130_fd_sc_hd__o21ba_1
X_2012_ _2289_/A _2012_/B vssd1 vssd1 vccd1 vccd1 _2012_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_70_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2914_ _2914_/A _2914_/B _2914_/C vssd1 vssd1 vccd1 vccd1 _2924_/C sky130_fd_sc_hd__and3_1
X_2845_ hold996/X _1646_/Y _2079_/B _3130_/A vssd1 vssd1 vccd1 vccd1 _2845_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_5_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2776_ _2082_/D _2771_/A _2759_/B _2690_/X vssd1 vssd1 vccd1 vccd1 _2776_/X sky130_fd_sc_hd__a2bb2o_1
Xhold101 _3466_/Q vssd1 vssd1 vccd1 vccd1 hold101/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold123 _3729_/Q vssd1 vssd1 vccd1 vccd1 hold123/X sky130_fd_sc_hd__dlygate4sd3_1
X_1727_ _1889_/A _1722_/X _2087_/A vssd1 vssd1 vccd1 vccd1 _1727_/Y sky130_fd_sc_hd__o21ai_1
Xhold112 _2593_/X vssd1 vssd1 vccd1 vccd1 _3529_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold134 _2375_/X vssd1 vssd1 vccd1 vccd1 _3342_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold156 _2614_/X vssd1 vssd1 vccd1 vccd1 _3547_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold167 _3730_/Q vssd1 vssd1 vccd1 vccd1 hold167/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1658_ _3630_/Q _2741_/B _2669_/C vssd1 vssd1 vccd1 vccd1 _1672_/B sky130_fd_sc_hd__a21oi_1
Xhold145 _3229_/Q vssd1 vssd1 vccd1 vccd1 hold145/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold178 _2225_/X vssd1 vssd1 vccd1 vccd1 _3260_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold189 _3215_/Q vssd1 vssd1 vccd1 vccd1 hold189/X sky130_fd_sc_hd__dlygate4sd3_1
X_3328_ _3447_/CLK _3328_/D vssd1 vssd1 vccd1 vccd1 _3328_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3259_ _3322_/CLK _3259_/D vssd1 vssd1 vccd1 vccd1 _3259_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2466__A0 _2648_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2218__A0 _2660_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold690 _2236_/X vssd1 vssd1 vccd1 vccd1 _3267_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_26_wb_clk_i_A clkbuf_3_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_59_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2209__A0 _2653_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2630_ hold27/X _2658_/A0 _2632_/S vssd1 vssd1 vccd1 vccd1 hold28/A sky130_fd_sc_hd__mux2_1
XFILLER_0_40_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2561_ hold243/X _2361_/A _2562_/S vssd1 vssd1 vccd1 vccd1 _2561_/X sky130_fd_sc_hd__mux2_1
Xscrapcpu_158 vssd1 vssd1 vccd1 vccd1 scrapcpu_158/HI io_oeb[0] sky130_fd_sc_hd__conb_1
Xscrapcpu_169 vssd1 vssd1 vccd1 vccd1 scrapcpu_169/HI io_oeb[27] sky130_fd_sc_hd__conb_1
XFILLER_0_2_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2492_ _2651_/A0 hold441/X _2494_/S vssd1 vssd1 vccd1 vccd1 _2492_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_49_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3113_ _3126_/A _3113_/B vssd1 vssd1 vccd1 vccd1 _3113_/X sky130_fd_sc_hd__or2_1
XFILLER_0_65_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3044_ _3045_/B _3045_/D _3045_/A vssd1 vssd1 vccd1 vccd1 _3044_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__2448__A0 _3196_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2620__A0 _2655_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1974__A2 _1922_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2828_ hold918/X _2871_/A _2746_/Y _2876_/B vssd1 vssd1 vccd1 vccd1 _2828_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_5_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2759_ _2759_/A _2759_/B vssd1 vssd1 vccd1 vccd1 _2759_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_60_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2923__B2 _2940_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2923__A1 _1712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2055__A _2955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout73 _2653_/A0 vssd1 vssd1 vccd1 vccd1 _2363_/A sky130_fd_sc_hd__buf_4
XANTENNA__2611__A0 _2660_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout95 _2089_/X vssd1 vssd1 vccd1 vccd1 _2353_/A sky130_fd_sc_hd__clkbuf_4
Xfanout84 _2475_/A1 vssd1 vssd1 vccd1 vccd1 _2643_/A1 sky130_fd_sc_hd__buf_2
XANTENNA__1833__S _1937_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output38_A _3768_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2602__A0 _3203_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3731_ _3732_/CLK _3731_/D vssd1 vssd1 vccd1 vccd1 hold99/A sky130_fd_sc_hd__dfxtp_1
X_1992_ hold99/A _3477_/Q _3415_/Q _3427_/Q _1996_/S _2185_/C vssd1 vssd1 vccd1 vccd1
+ _1993_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_27_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_35_wb_clk_i clkbuf_3_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3436_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_15_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3662_ _3662_/CLK hold80/X vssd1 vssd1 vccd1 vccd1 hold79/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3593_ _3745_/CLK _3593_/D vssd1 vssd1 vccd1 vccd1 _3593_/Q sky130_fd_sc_hd__dfxtp_1
X_2613_ hold47/X _3193_/A0 _2618_/S vssd1 vssd1 vccd1 vccd1 hold48/A sky130_fd_sc_hd__mux2_1
XFILLER_0_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2544_ _3201_/A1 hold727/X _2548_/S vssd1 vssd1 vccd1 vccd1 _2544_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_50_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2475_ hold171/X _2475_/A1 _2478_/S vssd1 vssd1 vccd1 vccd1 _2475_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_76_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1979__A _1979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3027_ _3027_/A _3027_/B vssd1 vssd1 vccd1 vccd1 _3027_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__2841__B1 _2940_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1698__B _2854_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_394 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1889__A _1889_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2260_ _2365_/A _2619_/A vssd1 vssd1 vccd1 vccd1 _2266_/S sky130_fd_sc_hd__nand2_4
X_2191_ hold207/X _2652_/A0 _2192_/S vssd1 vssd1 vccd1 vccd1 _2191_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3076__B1 _3048_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2407__B _2598_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1721__S1 _2228_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1975_ _2867_/B vssd1 vssd1 vccd1 vccd1 _2689_/B sky130_fd_sc_hd__inv_2
XFILLER_0_55_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3714_ _3714_/CLK _3714_/D vssd1 vssd1 vccd1 vccd1 _3714_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3645_ _3646_/CLK _3645_/D vssd1 vssd1 vccd1 vccd1 _3645_/Q sky130_fd_sc_hd__dfxtp_1
X_3576_ _3724_/CLK _3576_/D vssd1 vssd1 vccd1 vccd1 _3576_/Q sky130_fd_sc_hd__dfxtp_1
X_2527_ hold325/X _2363_/A _2527_/S vssd1 vssd1 vccd1 vccd1 _2527_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_11_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2458_ _2570_/A _2500_/B vssd1 vssd1 vccd1 vccd1 _2464_/S sky130_fd_sc_hd__nand2_4
XFILLER_0_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold27 hold27/A vssd1 vssd1 vccd1 vccd1 hold27/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold16 hold16/A vssd1 vssd1 vccd1 vccd1 hold16/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold38 hold38/A vssd1 vssd1 vccd1 vccd1 hold38/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 hold49/A vssd1 vssd1 vccd1 vccd1 hold49/X sky130_fd_sc_hd__dlygate4sd3_1
X_2389_ _2475_/A1 hold363/X _2392_/S vssd1 vssd1 vccd1 vccd1 _2389_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1960__S1 _2014_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2814__B1 _2731_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2052__B _3048_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2750__C1 _2859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2480__D_N _2428_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1760_ _1760_/A _1760_/B vssd1 vssd1 vccd1 vccd1 _1762_/C sky130_fd_sc_hd__nand2_1
XANTENNA__3058__B _3058_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold508 _2581_/X vssd1 vssd1 vccd1 vccd1 _3519_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1691_ _1701_/A _1691_/B vssd1 vssd1 vccd1 vccd1 _1694_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold519 _3663_/Q vssd1 vssd1 vccd1 vccd1 hold519/X sky130_fd_sc_hd__dlygate4sd3_1
X_3430_ _3665_/CLK _3430_/D vssd1 vssd1 vccd1 vccd1 _3430_/Q sky130_fd_sc_hd__dfxtp_1
X_3361_ _3654_/CLK _3361_/D vssd1 vssd1 vccd1 vccd1 _3361_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2312_ _2167_/C _2303_/X _2311_/Y _2298_/A vssd1 vssd1 vccd1 vccd1 _2318_/B sky130_fd_sc_hd__o211ai_4
XFILLER_0_57_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3292_ _3724_/CLK _3292_/D vssd1 vssd1 vccd1 vccd1 _3292_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2243_ _2653_/A0 hold559/X _2243_/S vssd1 vssd1 vccd1 vccd1 _2243_/X sky130_fd_sc_hd__mux2_1
X_2174_ _2315_/A _1707_/C _2173_/Y vssd1 vssd1 vccd1 vccd1 _2174_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_73_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_50_wb_clk_i clkbuf_3_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3718_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_75_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2024__A1 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1958_ _2244_/A _1953_/X _2087_/A vssd1 vssd1 vccd1 vccd1 _1958_/Y sky130_fd_sc_hd__o21ai_1
X_1889_ _1889_/A _1889_/B vssd1 vssd1 vccd1 vccd1 _1889_/Y sky130_fd_sc_hd__nor2_1
X_3628_ _3668_/CLK _3628_/D vssd1 vssd1 vccd1 vccd1 _3628_/Q sky130_fd_sc_hd__dfxtp_2
Xoutput39 _3769_/X vssd1 vssd1 vccd1 vccd1 io_oeb[9] sky130_fd_sc_hd__buf_12
Xoutput28 _3774_/X vssd1 vssd1 vccd1 vccd1 io_oeb[19] sky130_fd_sc_hd__buf_12
X_3559_ _3585_/CLK _3559_/D vssd1 vssd1 vccd1 vccd1 _3559_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1933__S1 _2228_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2799__C1 _2859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1841__S _2244_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2254__A1 _2089_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2930_ _1605_/Y _2935_/A _2941_/C _2928_/X _2885_/B vssd1 vssd1 vccd1 vccd1 _2930_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2861_ _3599_/Q _2861_/B _2861_/C vssd1 vssd1 vccd1 vccd1 _2861_/X sky130_fd_sc_hd__or3_1
X_1812_ _2228_/A _1801_/X _1808_/X _1811_/Y vssd1 vssd1 vccd1 vccd1 _1812_/X sky130_fd_sc_hd__a31o_1
X_2792_ _2082_/D _2788_/A _2759_/B _2675_/X vssd1 vssd1 vccd1 vccd1 _2792_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_25_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1743_ _2085_/C _1743_/B vssd1 vssd1 vccd1 vccd1 _1743_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_40_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold316 _2455_/X vssd1 vssd1 vccd1 vccd1 _3415_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1674_ _1677_/B vssd1 vssd1 vccd1 vccd1 _1676_/B sky130_fd_sc_hd__inv_2
XANTENNA__2701__A _3594_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold305 _3319_/Q vssd1 vssd1 vccd1 vccd1 hold305/X sky130_fd_sc_hd__dlygate4sd3_1
X_3413_ _3733_/CLK hold34/X vssd1 vssd1 vccd1 vccd1 hold33/A sky130_fd_sc_hd__dfxtp_1
Xhold327 _3659_/Q vssd1 vssd1 vccd1 vccd1 hold327/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold349 _3648_/Q vssd1 vssd1 vccd1 vccd1 hold349/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold338 _2649_/X vssd1 vssd1 vccd1 vccd1 _3577_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3344_ _3344_/CLK hold88/X vssd1 vssd1 vccd1 vccd1 hold87/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1005 _2168_/X vssd1 vssd1 vccd1 vccd1 _3224_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3275_ _3308_/CLK hold76/X vssd1 vssd1 vccd1 vccd1 hold75/A sky130_fd_sc_hd__dfxtp_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2226_ _2653_/A0 hold319/X _2226_/S vssd1 vssd1 vccd1 vccd1 _2226_/X sky130_fd_sc_hd__mux2_1
Xhold1016 _3152_/X vssd1 vssd1 vccd1 vccd1 _3712_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1027 _3226_/Q vssd1 vssd1 vccd1 vccd1 _2316_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1038 _3347_/Q vssd1 vssd1 vccd1 vccd1 hold1038/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1049 _3292_/Q vssd1 vssd1 vccd1 vccd1 _2268_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2157_ _3225_/Q _1821_/X _3059_/A vssd1 vssd1 vccd1 vccd1 _2167_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_88_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2088_ _2640_/A _2290_/A vssd1 vssd1 vccd1 vccd1 _2100_/S sky130_fd_sc_hd__nor2_2
XANTENNA__1987__A _2006_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1756__B1 _2195_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold861 _2952_/Y vssd1 vssd1 vccd1 vccd1 _2954_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold850 _3602_/Q vssd1 vssd1 vccd1 vccd1 hold850/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold872 _3721_/Q vssd1 vssd1 vccd1 vccd1 _3171_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold894 _2784_/X vssd1 vssd1 vccd1 vccd1 _3597_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout87_A _2093_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold883 _3325_/Q vssd1 vssd1 vccd1 vccd1 hold883/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_16_wb_clk_i_A clkbuf_3_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__2484__A1 _2357_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2521__A _2640_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_55_wb_clk_i_A clkbuf_leaf_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__2711__A2 _2868_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3060_ _3228_/Q _3096_/C vssd1 vssd1 vccd1 vccd1 _3060_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__3121__C1 _3055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2011_ hold73/A hold21/A hold85/A _3221_/Q _2085_/B _2014_/A vssd1 vssd1 vccd1 vccd1
+ _2012_/B sky130_fd_sc_hd__mux4_1
XANTENNA__2475__A1 _2475_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2913_ _3618_/Q _2914_/C _2914_/A vssd1 vssd1 vccd1 vccd1 _2913_/Y sky130_fd_sc_hd__a21oi_1
X_2844_ _3599_/Q _2871_/A _2843_/Y _2876_/B vssd1 vssd1 vccd1 vccd1 _2844_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_72_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2775_ _2775_/A _2775_/B _2775_/C vssd1 vssd1 vccd1 vccd1 _2790_/A sky130_fd_sc_hd__and3_1
Xhold124 _3187_/X vssd1 vssd1 vccd1 vccd1 _3729_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold135 _3283_/Q vssd1 vssd1 vccd1 vccd1 hold135/X sky130_fd_sc_hd__dlygate4sd3_1
X_1726_ _2245_/B _1726_/B vssd1 vssd1 vccd1 vccd1 _1726_/Y sky130_fd_sc_hd__nand2_1
Xhold113 _3584_/Q vssd1 vssd1 vccd1 vccd1 hold113/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold102 _2519_/X vssd1 vssd1 vccd1 vccd1 _3466_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 _3188_/X vssd1 vssd1 vccd1 vccd1 _3730_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold157 _3393_/Q vssd1 vssd1 vccd1 vccd1 hold157/X sky130_fd_sc_hd__dlygate4sd3_1
X_1657_ _2712_/A _3627_/Q vssd1 vssd1 vccd1 vccd1 _2741_/B sky130_fd_sc_hd__nand2_2
Xhold146 _2187_/X vssd1 vssd1 vccd1 vccd1 _3229_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold179 _3511_/Q vssd1 vssd1 vccd1 vccd1 hold179/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3327_ _3724_/CLK _3327_/D vssd1 vssd1 vccd1 vccd1 _3327_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3258_ _3270_/CLK _3258_/D vssd1 vssd1 vccd1 vccd1 _3258_/Q sky130_fd_sc_hd__dfxtp_1
X_3189_ hold99/X _3203_/A1 _3191_/S vssd1 vssd1 vccd1 vccd1 _3189_/X sky130_fd_sc_hd__mux2_1
X_2209_ _2653_/A0 hold775/X _2209_/S vssd1 vssd1 vccd1 vccd1 _2209_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_68_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold680 _2262_/X vssd1 vssd1 vccd1 vccd1 _3287_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold691 _3738_/Q vssd1 vssd1 vccd1 vccd1 hold691/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2457__A1 _2363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2219__C _2219_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2560_ hold109/X _3203_/A1 _2562_/S vssd1 vssd1 vccd1 vccd1 _2560_/X sky130_fd_sc_hd__mux2_1
Xscrapcpu_159 vssd1 vssd1 vccd1 vccd1 scrapcpu_159/HI io_oeb[1] sky130_fd_sc_hd__conb_1
XFILLER_0_2_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2491_ _2650_/A0 hold681/X _2494_/S vssd1 vssd1 vccd1 vccd1 _2491_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_10_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3112_ hold803/X _3016_/X _3183_/B vssd1 vssd1 vccd1 vccd1 _3113_/B sky130_fd_sc_hd__mux2_1
X_3043_ _3063_/B _3039_/X _3042_/Y vssd1 vssd1 vccd1 vccd1 _3043_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_85_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout137_A _1954_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2827_ hold978/X _2824_/X _2826_/X _2817_/X _2859_/A vssd1 vssd1 vccd1 vccd1 _2827_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_26_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2384__A0 _2659_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2758_ _2755_/Y _2756_/X _2738_/A _2738_/B vssd1 vssd1 vccd1 vccd1 _2775_/A sky130_fd_sc_hd__a211oi_2
X_1709_ _2497_/A _2496_/C vssd1 vssd1 vccd1 vccd1 _2071_/D sky130_fd_sc_hd__or2_1
X_2689_ _3596_/Q _2689_/B vssd1 vssd1 vccd1 vccd1 _2705_/B sky130_fd_sc_hd__nand2_1
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2439__A1 _2355_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_5_wb_clk_i clkbuf_leaf_5_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3665_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_49_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2072__C1 _2495_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout74 _2099_/X vssd1 vssd1 vccd1 vccd1 _2653_/A0 sky130_fd_sc_hd__buf_4
XFILLER_0_64_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout85 _2093_/X vssd1 vssd1 vccd1 vccd1 _2475_/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout96 _2245_/C vssd1 vssd1 vccd1 vccd1 _2480_/C sky130_fd_sc_hd__buf_6
XFILLER_0_36_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1991_ _1889_/A _1987_/Y _1989_/Y _1990_/Y vssd1 vssd1 vccd1 vccd1 _1991_/X sky130_fd_sc_hd__a31o_1
X_3730_ _3732_/CLK _3730_/D vssd1 vssd1 vccd1 vccd1 _3730_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2063__C1 _1979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3661_ _3661_/CLK _3661_/D vssd1 vssd1 vccd1 vccd1 _3661_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3592_ _3592_/CLK _3592_/D vssd1 vssd1 vccd1 vccd1 _3592_/Q sky130_fd_sc_hd__dfxtp_1
X_2612_ _2640_/B _2612_/B vssd1 vssd1 vccd1 vccd1 _2618_/S sky130_fd_sc_hd__nor2_2
XANTENNA__2366__A0 _3193_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2543_ _2353_/A hold641/X _2548_/S vssd1 vssd1 vccd1 vccd1 _2543_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_50_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2118__A0 _2652_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2474_ hold205/X _3194_/A0 _2478_/S vssd1 vssd1 vccd1 vccd1 _2474_/X sky130_fd_sc_hd__mux2_1
X_3026_ _3027_/A _3026_/B _3027_/B _3035_/A vssd1 vssd1 vccd1 vccd1 _3036_/B sky130_fd_sc_hd__or4b_1
XANTENNA__1698__C _1922_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1995__A _2185_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwire109 _1629_/Y vssd1 vssd1 vccd1 vccd1 wire109/X sky130_fd_sc_hd__buf_1
XFILLER_0_61_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2109__A0 _3196_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2899__A1 _2876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2190_ hold241/X _2651_/A0 _2192_/S vssd1 vssd1 vccd1 vccd1 _2190_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_1_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2587__A0 _3195_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1974_ hold815/X _1922_/B _1972_/X _1973_/X vssd1 vssd1 vccd1 vccd1 _2867_/B sky130_fd_sc_hd__o22a_4
X_3713_ _3714_/CLK _3713_/D vssd1 vssd1 vccd1 vccd1 _3713_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3644_ _3674_/CLK _3644_/D vssd1 vssd1 vccd1 vccd1 _3644_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2339__B1 _3108_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3575_ _3575_/CLK _3575_/D vssd1 vssd1 vccd1 vccd1 _3575_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2526_ hold295/X _2361_/A _2527_/S vssd1 vssd1 vccd1 vccd1 _2526_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_11_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2457_ hold105/X _2363_/A _2457_/S vssd1 vssd1 vccd1 vccd1 _2457_/X sky130_fd_sc_hd__mux2_1
Xhold28 hold28/A vssd1 vssd1 vccd1 vccd1 hold28/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold17 hold17/A vssd1 vssd1 vccd1 vccd1 hold17/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold39 hold39/A vssd1 vssd1 vccd1 vccd1 hold39/X sky130_fd_sc_hd__dlygate4sd3_1
X_2388_ _3194_/A0 hold753/X _2392_/S vssd1 vssd1 vccd1 vccd1 _2388_/X sky130_fd_sc_hd__mux2_1
X_3009_ _2310_/B _3063_/A _3124_/B vssd1 vssd1 vccd1 vccd1 _3010_/B sky130_fd_sc_hd__o21a_1
XANTENNA__2814__A1 _2797_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2275__C1 _3058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2578__A0 _2655_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2227__C _2228_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1839__S _2244_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2569__A0 _2660_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold509 _3356_/Q vssd1 vssd1 vccd1 vccd1 hold509/X sky130_fd_sc_hd__dlygate4sd3_1
X_1690_ _2846_/B _1690_/B vssd1 vssd1 vccd1 vccd1 _1691_/B sky130_fd_sc_hd__nand2_1
X_3360_ _3387_/CLK _3360_/D vssd1 vssd1 vccd1 vccd1 _3360_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2311_ _2308_/Y _2311_/B _2311_/C vssd1 vssd1 vccd1 vccd1 _2311_/Y sky130_fd_sc_hd__nand3b_2
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3291_ _3387_/CLK _3291_/D vssd1 vssd1 vccd1 vccd1 _3291_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2242_ _2652_/A0 hold699/X _2243_/S vssd1 vssd1 vccd1 vccd1 _2242_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_73_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2173_ _2153_/A _2301_/C _1821_/X _2153_/Y vssd1 vssd1 vccd1 vccd1 _2173_/Y sky130_fd_sc_hd__a31oi_2
XFILLER_0_75_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1957_ _3771_/A _2005_/S _2006_/A _1956_/Y vssd1 vssd1 vccd1 vccd1 _1957_/X sky130_fd_sc_hd__a211o_1
X_1888_ _3729_/Q hold97/A hold33/A _3425_/Q _1996_/S _2185_/C vssd1 vssd1 vccd1 vccd1
+ _1889_/B sky130_fd_sc_hd__mux4_1
XANTENNA__1783__A1 _1889_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3627_ _3637_/CLK _3627_/D vssd1 vssd1 vccd1 vccd1 _3627_/Q sky130_fd_sc_hd__dfxtp_2
X_3558_ _3558_/CLK hold64/X vssd1 vssd1 vccd1 vccd1 hold63/A sky130_fd_sc_hd__dfxtp_1
Xoutput29 _3774_/A vssd1 vssd1 vccd1 vccd1 io_oeb[20] sky130_fd_sc_hd__buf_12
X_2509_ hold515/X _3201_/A1 _2513_/S vssd1 vssd1 vccd1 vccd1 _2509_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2732__B1 _2731_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3489_ _3744_/CLK _3489_/D vssd1 vssd1 vccd1 vccd1 _3489_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2344__A _3108_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_45_wb_clk_i_A clkbuf_3_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_27_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2860_ _3597_/Q _3596_/Q _3595_/Q vssd1 vssd1 vccd1 vccd1 _2861_/C sky130_fd_sc_hd__or3_1
X_1811_ _2228_/A _1777_/X _2195_/B vssd1 vssd1 vccd1 vccd1 _1811_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__3203__A1 _3203_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2791_ _2790_/A _2790_/B _2718_/B vssd1 vssd1 vccd1 vccd1 _2791_/Y sky130_fd_sc_hd__a21oi_1
X_1742_ hold87/A _3302_/Q _2244_/B vssd1 vssd1 vccd1 vccd1 _1743_/B sky130_fd_sc_hd__mux2_1
Xhold317 _3389_/Q vssd1 vssd1 vccd1 vccd1 hold317/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1673_ _2669_/C _2742_/B _1673_/C vssd1 vssd1 vccd1 vccd1 _1677_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_13_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2701__B _2701_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold306 _2335_/X vssd1 vssd1 vccd1 vccd1 _3319_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3412_ _3592_/CLK hold10/X vssd1 vssd1 vccd1 vccd1 hold9/A sky130_fd_sc_hd__dfxtp_1
Xhold328 _2984_/X vssd1 vssd1 vccd1 vccd1 _3659_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold339 _3266_/Q vssd1 vssd1 vccd1 vccd1 hold339/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2190__A1 _2651_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3343_ _3344_/CLK _3343_/D vssd1 vssd1 vccd1 vccd1 _3343_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1006 _3630_/Q vssd1 vssd1 vccd1 vccd1 _2034_/B sky130_fd_sc_hd__clkbuf_2
X_3274_ _3666_/CLK _3274_/D vssd1 vssd1 vccd1 vccd1 _3274_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2225_ _2652_/A0 hold177/X _2226_/S vssd1 vssd1 vccd1 vccd1 _2225_/X sky130_fd_sc_hd__mux2_1
Xhold1017 _3225_/Q vssd1 vssd1 vccd1 vccd1 _1638_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1028 _2172_/X vssd1 vssd1 vccd1 vccd1 _2175_/B1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1039 _2043_/X vssd1 vssd1 vccd1 vccd1 _3347_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2156_ _3709_/Q _2156_/B vssd1 vssd1 vccd1 vccd1 _2164_/B sky130_fd_sc_hd__xnor2_1
X_2087_ _2087_/A _2087_/B _2480_/C vssd1 vssd1 vccd1 vccd1 _2290_/A sky130_fd_sc_hd__or3_4
XFILLER_0_8_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2989_ hold489/X _1760_/B _2992_/S vssd1 vssd1 vccd1 vccd1 _2989_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1756__A1 _2479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2953__B1 _1979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold862 _2954_/Y vssd1 vssd1 vccd1 vccd1 _3632_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold840 _3314_/Q vssd1 vssd1 vccd1 vccd1 hold840/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold851 _2834_/X vssd1 vssd1 vccd1 vccd1 _3602_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold873 _3171_/X vssd1 vssd1 vccd1 vccd1 hold873/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold884 _2345_/X vssd1 vssd1 vccd1 vccd1 _2346_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold895 _3326_/Q vssd1 vssd1 vccd1 vccd1 hold895/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2074__A _2074_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3197__A0 _3197_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1747__A1 _2244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_1_wb_clk_i_A clkbuf_leaf_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__2013__S _2085_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2010_ _2244_/A _2006_/Y _2008_/X _2009_/Y vssd1 vssd1 vccd1 vccd1 _2010_/X sky130_fd_sc_hd__a31o_1
Xclkbuf_leaf_29_wb_clk_i clkbuf_3_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3732_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_2912_ hold497/X _2940_/B2 _2868_/D _1712_/A vssd1 vssd1 vccd1 vccd1 _2912_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_45_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2843_ _2871_/A _2843_/B vssd1 vssd1 vccd1 vccd1 _2843_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_57_198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2774_ _2775_/B _2775_/C _2775_/A vssd1 vssd1 vccd1 vccd1 _2774_/Y sky130_fd_sc_hd__a21oi_1
X_1725_ _3472_/Q _3490_/Q _1988_/S vssd1 vssd1 vccd1 vccd1 _1726_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_5_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold125 _3741_/Q vssd1 vssd1 vccd1 vccd1 hold125/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold114 _2657_/X vssd1 vssd1 vccd1 vccd1 _3584_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold103 _3383_/Q vssd1 vssd1 vccd1 vccd1 hold103/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold147 _3284_/Q vssd1 vssd1 vccd1 vccd1 hold147/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold136 _2257_/X vssd1 vssd1 vccd1 vccd1 _3283_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold158 _2427_/X vssd1 vssd1 vccd1 vccd1 _3393_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1656_ _2717_/B _2854_/A vssd1 vssd1 vccd1 vccd1 _2669_/C sky130_fd_sc_hd__nand2_1
Xhold169 _3382_/Q vssd1 vssd1 vccd1 vccd1 hold169/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3326_ _3721_/CLK _3326_/D vssd1 vssd1 vccd1 vccd1 _3326_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3257_ _3270_/CLK _3257_/D vssd1 vssd1 vccd1 vccd1 _3257_/Q sky130_fd_sc_hd__dfxtp_1
X_3188_ hold167/X _2357_/A _3191_/S vssd1 vssd1 vccd1 vccd1 _3188_/X sky130_fd_sc_hd__mux2_1
X_2208_ _2652_/A0 hold457/X _2209_/S vssd1 vssd1 vccd1 vccd1 _2208_/X sky130_fd_sc_hd__mux2_1
X_2139_ _3722_/Q _2155_/A vssd1 vssd1 vccd1 vccd1 _2161_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_48_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1937__S _1937_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1977__B2 _2854_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold670 _2548_/X vssd1 vssd1 vccd1 vccd1 _3491_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold681 _3444_/Q vssd1 vssd1 vccd1 vccd1 hold681/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold692 _3197_/X vssd1 vssd1 vccd1 vccd1 _3738_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2219__D _3348_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2862__C1 _2797_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1968__A1 _2479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2490_ _2355_/A hold449/X _2494_/S vssd1 vssd1 vccd1 vccd1 _2490_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_50_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3111_ hold803/X _3120_/A _3110_/X _3055_/A vssd1 vssd1 vccd1 vccd1 _3111_/X sky130_fd_sc_hd__o211a_1
X_3042_ _3063_/B _3039_/X _3055_/A vssd1 vssd1 vccd1 vccd1 _3042_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_73_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_327 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1959__A1 _2244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2826_ hold918/X _1696_/Y _2940_/B2 hold621/X _2825_/Y vssd1 vssd1 vccd1 vccd1 _2826_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_5_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2908__B1 _2940_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2757_ _2738_/A _2738_/B _2755_/Y _2756_/X vssd1 vssd1 vccd1 vccd1 _2757_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_30_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1708_ _2054_/A _3048_/B vssd1 vssd1 vccd1 vccd1 _2496_/C sky130_fd_sc_hd__or2_1
X_2688_ _2735_/A _2703_/C _2754_/A vssd1 vssd1 vccd1 vccd1 _2755_/B sky130_fd_sc_hd__o21ai_2
X_1639_ _3081_/B _2302_/A vssd1 vssd1 vccd1 vccd1 _3096_/B sky130_fd_sc_hd__or2_4
XFILLER_0_41_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3309_ _3721_/CLK hold42/X vssd1 vssd1 vccd1 vccd1 hold41/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2352__A _2640_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout86 _2650_/A0 vssd1 vssd1 vccd1 vccd1 _2357_/A sky130_fd_sc_hd__buf_4
Xfanout97 _2987_/S vssd1 vssd1 vccd1 vccd1 _2999_/S sky130_fd_sc_hd__clkbuf_8
Xfanout75 _2659_/A0 vssd1 vssd1 vccd1 vccd1 _3197_/A0 sky130_fd_sc_hd__buf_4
XANTENNA__2375__A1 _2650_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2071__B _2076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1886__B1 _2087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1981__S0 _1981_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2246__B _3199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1990_ _1889_/A _1985_/X _2428_/C vssd1 vssd1 vccd1 vccd1 _1990_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_55_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3660_ _3661_/CLK _3660_/D vssd1 vssd1 vccd1 vccd1 _3660_/Q sky130_fd_sc_hd__dfxtp_1
X_3591_ _3745_/CLK _3591_/D vssd1 vssd1 vccd1 vccd1 _3591_/Q sky130_fd_sc_hd__dfxtp_1
X_2611_ _2660_/A0 hold431/X _2611_/S vssd1 vssd1 vccd1 vccd1 _2611_/X sky130_fd_sc_hd__mux2_1
X_2542_ _2619_/A _2598_/B vssd1 vssd1 vccd1 vccd1 _2548_/S sky130_fd_sc_hd__nand2_4
X_2473_ hold307/X _3193_/A0 _2478_/S vssd1 vssd1 vccd1 vccd1 _2473_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_44_wb_clk_i clkbuf_3_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3695_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_3025_ _3086_/A _3025_/B _3027_/B vssd1 vssd1 vccd1 vccd1 _3677_/D sky130_fd_sc_hd__and3_1
XANTENNA__2841__A2 _1696_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_168 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2809_ _2809_/A _2809_/B _2808_/X vssd1 vssd1 vccd1 vccd1 _2809_/X sky130_fd_sc_hd__or3b_1
XFILLER_0_69_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2596__A1 _2361_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1860__S _2085_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2520__A1 _3198_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2284__A0 _2355_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1973_ input2/X _1920_/B _1677_/X vssd1 vssd1 vccd1 vccd1 _1973_/X sky130_fd_sc_hd__a21o_1
X_3712_ _3714_/CLK _3712_/D vssd1 vssd1 vccd1 vccd1 _3712_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3643_ _3646_/CLK _3643_/D vssd1 vssd1 vccd1 vccd1 _3643_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2720__A _3594_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2339__A1 _2648_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3574_ _3575_/CLK _3574_/D vssd1 vssd1 vccd1 vccd1 _3574_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2525_ hold77/X _3203_/A1 _2527_/S vssd1 vssd1 vccd1 vccd1 hold78/A sky130_fd_sc_hd__mux2_1
XFILLER_0_87_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2456_ hold35/X _2361_/A _2457_/S vssd1 vssd1 vccd1 vccd1 hold36/A sky130_fd_sc_hd__mux2_1
Xhold29 hold29/A vssd1 vssd1 vccd1 vccd1 hold29/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold18 hold18/A vssd1 vssd1 vccd1 vccd1 hold18/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2511__A1 _3203_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2387_ _3193_/A0 hold751/X _2392_/S vssd1 vssd1 vccd1 vccd1 _2387_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2167__A _3045_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3008_ _3014_/A _3045_/A vssd1 vssd1 vccd1 vccd1 _3063_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_19_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1945__S _2244_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_35_wb_clk_i_A clkbuf_3_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__2750__A1 hold918/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2266__A0 _3198_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2227__D _2480_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_3_7__f_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2310_ _3053_/B _2310_/B _3097_/C _3007_/A vssd1 vssd1 vccd1 vccd1 _2311_/B sky130_fd_sc_hd__or4_2
X_3290_ _3654_/CLK _3290_/D vssd1 vssd1 vccd1 vccd1 _3290_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2241_ _2651_/A0 hold771/X _2243_/S vssd1 vssd1 vccd1 vccd1 _2241_/X sky130_fd_sc_hd__mux2_1
X_2172_ _1707_/C _2169_/B _2315_/A vssd1 vssd1 vccd1 vccd1 _2172_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_75_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2715__A _3612_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2009__B1 _2087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1956_ _3330_/Q _2005_/S vssd1 vssd1 vccd1 vccd1 _1956_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_16_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1887_ _1889_/A _1883_/Y _1885_/Y _1886_/Y vssd1 vssd1 vccd1 vccd1 _1887_/X sky130_fd_sc_hd__a31o_1
XANTENNA_fanout112_A _2244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3626_ _3637_/CLK _3626_/D vssd1 vssd1 vccd1 vccd1 _3626_/Q sky130_fd_sc_hd__dfxtp_2
X_3557_ _3587_/CLK _3557_/D vssd1 vssd1 vccd1 vccd1 _3557_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput19 _3769_/A vssd1 vssd1 vccd1 vccd1 io_oeb[10] sky130_fd_sc_hd__buf_12
X_2508_ hold193/X _2353_/A _2513_/S vssd1 vssd1 vccd1 vccd1 _2508_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2732__A1 _2797_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3488_ _3539_/CLK _3488_/D vssd1 vssd1 vccd1 vccd1 _3488_/Q sky130_fd_sc_hd__dfxtp_1
X_2439_ hold968/X _2355_/A _2443_/S vssd1 vssd1 vccd1 vccd1 _3401_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_66_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_252 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1759__C1 _2022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold860_A _3632_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2184__C1 _3055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2239__A0 _2355_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1810_ _2479_/A _1794_/X _2228_/B vssd1 vssd1 vccd1 vccd1 _1810_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__2411__A0 _2658_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2790_ _2790_/A _2790_/B vssd1 vssd1 vccd1 vccd1 _2790_/X sky130_fd_sc_hd__or2_1
XFILLER_0_25_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1741_ _3296_/Q _3446_/Q _3580_/Q _3404_/Q _2005_/S _2014_/A vssd1 vssd1 vccd1 vccd1
+ _1741_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_7_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1672_ _3631_/Q _1672_/B vssd1 vssd1 vccd1 vccd1 _1677_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_40_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold307 _3430_/Q vssd1 vssd1 vccd1 vccd1 hold307/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1765__A2 _1922_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold318 _2423_/X vssd1 vssd1 vccd1 vccd1 _3389_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold329 _3446_/Q vssd1 vssd1 vccd1 vccd1 hold329/X sky130_fd_sc_hd__dlygate4sd3_1
X_3411_ _3419_/CLK _3411_/D vssd1 vssd1 vccd1 vccd1 _3411_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2175__C1 _3108_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3342_ _3344_/CLK _3342_/D vssd1 vssd1 vccd1 vccd1 _3342_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3273_ _3743_/CLK _3273_/D vssd1 vssd1 vccd1 vccd1 _3273_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1018 _3096_/B vssd1 vssd1 vccd1 vccd1 _1640_/C sky130_fd_sc_hd__buf_1
Xhold1007 _2075_/X vssd1 vssd1 vccd1 vccd1 _3630_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1029 _2175_/Y vssd1 vssd1 vccd1 vccd1 _3226_/D sky130_fd_sc_hd__dlygate4sd3_1
X_2224_ _2651_/A0 hold403/X _2226_/S vssd1 vssd1 vccd1 vccd1 _2224_/X sky130_fd_sc_hd__mux2_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2155_ _2155_/A _2155_/B vssd1 vssd1 vccd1 vccd1 _2156_/B sky130_fd_sc_hd__or2_1
X_2086_ _2087_/A _2087_/B _2480_/C vssd1 vssd1 vccd1 vccd1 _2237_/A sky130_fd_sc_hd__nor3_4
XFILLER_0_48_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2650__A0 _2650_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2988_ hold519/X _1760_/A _2992_/S vssd1 vssd1 vccd1 vccd1 _2988_/X sky130_fd_sc_hd__mux2_1
X_1939_ _1889_/A _1934_/X _2428_/C vssd1 vssd1 vccd1 vccd1 _1939_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_8_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold830 _3043_/Y vssd1 vssd1 vccd1 vccd1 _3683_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3609_ _3672_/CLK _3609_/D vssd1 vssd1 vccd1 vccd1 _3609_/Q sky130_fd_sc_hd__dfxtp_1
Xhold852 _3604_/Q vssd1 vssd1 vccd1 vccd1 hold852/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold841 _2325_/X vssd1 vssd1 vccd1 vccd1 _3314_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold863 _3718_/Q vssd1 vssd1 vccd1 vccd1 _3165_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold896 _3710_/Q vssd1 vssd1 vccd1 vccd1 _2161_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold874 _3172_/X vssd1 vssd1 vccd1 vccd1 _3721_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold885 _3723_/Q vssd1 vssd1 vccd1 vccd1 _3175_/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2469__A0 _3203_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2355__A _2355_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2911_ _2914_/B _2883_/Y _2910_/Y _3166_/C1 vssd1 vssd1 vccd1 vccd1 _2911_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_57_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3188__A1 _2357_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2842_ hold852/X _2824_/X _2840_/X _2841_/X _2859_/A vssd1 vssd1 vccd1 vccd1 _2842_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_5_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2773_ _2803_/A _2773_/B vssd1 vssd1 vccd1 vccd1 _2775_/C sky130_fd_sc_hd__or2_1
X_1724_ _2006_/A _1724_/B vssd1 vssd1 vccd1 vccd1 _1724_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_79_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold126 _3201_/X vssd1 vssd1 vccd1 vccd1 _3741_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold104 _2416_/X vssd1 vssd1 vccd1 vccd1 _3383_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold115 _3343_/Q vssd1 vssd1 vccd1 vccd1 hold115/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold148 _2258_/X vssd1 vssd1 vccd1 vccd1 _3284_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold137 _3469_/Q vssd1 vssd1 vccd1 vccd1 hold137/X sky130_fd_sc_hd__dlygate4sd3_1
X_1655_ _2669_/A _1713_/B vssd1 vssd1 vccd1 vccd1 _1659_/B sky130_fd_sc_hd__nor2_1
Xhold159 _3480_/Q vssd1 vssd1 vccd1 vccd1 hold159/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3325_ _3723_/CLK _3325_/D vssd1 vssd1 vccd1 vccd1 _3325_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3256_ _3270_/CLK _3256_/D vssd1 vssd1 vccd1 vccd1 _3256_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2207_ _2651_/A0 hold749/X _2209_/S vssd1 vssd1 vccd1 vccd1 _2207_/X sky130_fd_sc_hd__mux2_1
X_3187_ hold123/X _3201_/A1 _3191_/S vssd1 vssd1 vccd1 vccd1 _3187_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2138_ _3711_/Q _2138_/B vssd1 vssd1 vccd1 vccd1 _2164_/A sky130_fd_sc_hd__xnor2_1
X_2069_ hold473/X _2731_/A2 _2868_/D _2034_/X vssd1 vssd1 vccd1 vccd1 _2069_/X sky130_fd_sc_hd__o22a_1
XANTENNA__2623__A0 _2658_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold671 _3540_/Q vssd1 vssd1 vccd1 vccd1 hold671/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold660 _2286_/X vssd1 vssd1 vccd1 vccd1 _3301_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout92_A _3193_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold693 _3420_/Q vssd1 vssd1 vccd1 vccd1 hold693/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold682 _2491_/X vssd1 vssd1 vccd1 vccd1 _3444_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2085__A _2085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2090__A1 _3193_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3110_ _3126_/A _3110_/B vssd1 vssd1 vccd1 vccd1 _3110_/X sky130_fd_sc_hd__or2_1
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3041_ _3039_/X _3040_/Y _3055_/A vssd1 vssd1 vccd1 vccd1 _3041_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_73_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2825_ _2825_/A _2874_/B vssd1 vssd1 vccd1 vccd1 _2825_/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_45_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2908__A1 _1712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2756_ _2803_/A _2756_/B vssd1 vssd1 vccd1 vccd1 _2756_/X sky130_fd_sc_hd__or2_1
X_1707_ _2301_/A _1707_/B _1707_/C _3059_/B vssd1 vssd1 vccd1 vccd1 _2497_/A sky130_fd_sc_hd__or4b_2
X_2687_ _3595_/Q _2687_/B vssd1 vssd1 vccd1 vccd1 _2703_/C sky130_fd_sc_hd__and2_1
XFILLER_0_41_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1638_ _1638_/A _3059_/A vssd1 vssd1 vccd1 vccd1 _2302_/A sky130_fd_sc_hd__or2_1
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3308_ _3308_/CLK hold90/X vssd1 vssd1 vccd1 vccd1 hold89/A sky130_fd_sc_hd__dfxtp_1
X_3239_ _3585_/CLK _3239_/D vssd1 vssd1 vccd1 vccd1 _3239_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2633__A _2640_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout98 _2987_/S vssd1 vssd1 vccd1 vccd1 _2992_/S sky130_fd_sc_hd__clkbuf_4
Xfanout87 _2093_/X vssd1 vssd1 vccd1 vccd1 _2650_/A0 sky130_fd_sc_hd__buf_4
Xfanout76 _2097_/X vssd1 vssd1 vccd1 vccd1 _2659_/A0 sky130_fd_sc_hd__buf_4
XANTENNA__2071__C _3045_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold490 _2989_/X vssd1 vssd1 vccd1 vccd1 _3664_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1886__A1 _1889_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1981__S1 _1981_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1712__A _1712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1858__S _2085_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2063__A1 _2050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1810__A1 _2479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2610_ _2659_/A0 hold683/X _2611_/S vssd1 vssd1 vccd1 vccd1 _2610_/X sky130_fd_sc_hd__mux2_1
X_3590_ _3592_/CLK _3590_/D vssd1 vssd1 vccd1 vccd1 _3590_/Q sky130_fd_sc_hd__dfxtp_1
X_2541_ hold15/X _2660_/A0 _2541_/S vssd1 vssd1 vccd1 vccd1 hold16/A sky130_fd_sc_hd__mux2_1
X_2472_ _3192_/B _2549_/A vssd1 vssd1 vccd1 vccd1 _2478_/S sky130_fd_sc_hd__nor2_2
XFILLER_0_76_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1622__A _2480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3024_ _3024_/A _3080_/A vssd1 vssd1 vccd1 vccd1 _3027_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_92_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_13_wb_clk_i clkbuf_3_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3545_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__2826__B1 _2940_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout142_A _1988_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1801__A1 _2244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2808_ _2803_/B _2803_/C _2709_/C _2779_/A vssd1 vssd1 vccd1 vccd1 _2808_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3003__B1 _2961_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_25_wb_clk_i_A clkbuf_3_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_2739_ _2738_/A _2738_/B _2718_/B vssd1 vssd1 vccd1 vccd1 _2739_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_5_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2293__A1 _2650_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2363__A _2363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2045__A1 _2085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2082__B _2961_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output36_A _1705_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2036__A1 _2731_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1972_ input8/X _2022_/A _1762_/X _1971_/Y vssd1 vssd1 vccd1 vccd1 _1972_/X sky130_fd_sc_hd__o211a_1
X_3711_ _3714_/CLK _3711_/D vssd1 vssd1 vccd1 vccd1 _3711_/Q sky130_fd_sc_hd__dfxtp_1
X_3642_ _3672_/CLK _3642_/D vssd1 vssd1 vccd1 vccd1 _3642_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2339__A2 _2619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3573_ _3585_/CLK _3573_/D vssd1 vssd1 vccd1 vccd1 _3573_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2524_ hold181/X _2357_/A _2527_/S vssd1 vssd1 vccd1 vccd1 _2524_/X sky130_fd_sc_hd__mux2_1
X_2455_ hold315/X _3203_/A1 _2457_/S vssd1 vssd1 vccd1 vccd1 _2455_/X sky130_fd_sc_hd__mux2_1
X_2386_ _2640_/A _3192_/A vssd1 vssd1 vccd1 vccd1 _2392_/S sky130_fd_sc_hd__or2_4
Xhold19 hold19/A vssd1 vssd1 vccd1 vccd1 hold19/X sky130_fd_sc_hd__dlygate4sd3_1
X_3007_ _3007_/A _3045_/D vssd1 vssd1 vccd1 vccd1 _3124_/B sky130_fd_sc_hd__or2_1
XFILLER_0_36_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2275__A1 _1716_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2027__B2 _2854_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1881__S0 _1988_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2018__A1 _2479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2240_ _2357_/A hold543/X _2243_/S vssd1 vssd1 vccd1 vccd1 _2240_/X sky130_fd_sc_hd__mux2_1
X_2171_ _2153_/A _3158_/A _2171_/B1 _2169_/B _3055_/A vssd1 vssd1 vccd1 vccd1 _2171_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA__2257__A1 _2658_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2009__A1 _2244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1955_ _2006_/A _1955_/B vssd1 vssd1 vccd1 vccd1 _1955_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__1768__B1 _2731_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1886_ _1889_/A _1881_/X _2087_/A vssd1 vssd1 vccd1 vccd1 _1886_/Y sky130_fd_sc_hd__o21ai_1
X_3625_ _3674_/CLK _3625_/D vssd1 vssd1 vccd1 vccd1 _3625_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3556_ _3583_/CLK _3556_/D vssd1 vssd1 vccd1 vccd1 _3556_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout105_A _1716_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2507_ _2612_/B _3185_/B vssd1 vssd1 vccd1 vccd1 _2513_/S sky130_fd_sc_hd__nor2_2
XFILLER_0_11_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3487_ _3744_/CLK _3487_/D vssd1 vssd1 vccd1 vccd1 _3487_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2438_ hold941/X _2648_/A0 _2443_/S vssd1 vssd1 vccd1 vccd1 _2438_/X sky130_fd_sc_hd__mux2_1
X_2369_ _3196_/A0 hold291/X _2371_/S vssd1 vssd1 vccd1 vccd1 _2369_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2248__A1 _2355_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2420__A1 _3198_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2487__A1 _2363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2088__A _2640_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1998__B1 _2428_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2535__B _3199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1740_ _1739_/X _1738_/X _1736_/X _1737_/X _2289_/A _2479_/B vssd1 vssd1 vccd1 vccd1
+ _1755_/B sky130_fd_sc_hd__mux4_2
XANTENNA__1845__S0 _2000_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1671_ _2876_/B _1979_/A _2822_/A vssd1 vssd1 vccd1 vccd1 _2080_/B sky130_fd_sc_hd__and3_1
Xhold308 _2473_/X vssd1 vssd1 vccd1 vccd1 _3430_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold319 _3261_/Q vssd1 vssd1 vccd1 vccd1 hold319/X sky130_fd_sc_hd__dlygate4sd3_1
X_3410_ _3419_/CLK _3410_/D vssd1 vssd1 vccd1 vccd1 _3410_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3341_ _3344_/CLK hold38/X vssd1 vssd1 vccd1 vccd1 hold37/A sky130_fd_sc_hd__dfxtp_1
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3272_ _3743_/CLK _3272_/D vssd1 vssd1 vccd1 vccd1 _3272_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1008 _3611_/Q vssd1 vssd1 vccd1 vccd1 _2999_/A1 sky130_fd_sc_hd__buf_1
Xhold1019 _3607_/Q vssd1 vssd1 vccd1 vccd1 _1926_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2478__A1 _3198_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2223_ _2357_/A hold161/X _2226_/S vssd1 vssd1 vccd1 vccd1 _2223_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_84_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2154_ _3721_/Q _2154_/B vssd1 vssd1 vccd1 vccd1 _2155_/B sky130_fd_sc_hd__nor2_1
X_2085_ _2085_/A _2085_/B _2085_/C _2480_/C vssd1 vssd1 vccd1 vccd1 _2640_/A sky130_fd_sc_hd__or4_4
XFILLER_0_48_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2987_ hold79/X _2987_/A1 _2987_/S vssd1 vssd1 vccd1 vccd1 hold80/A sky130_fd_sc_hd__mux2_1
XFILLER_0_16_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1938_ _2245_/B _1938_/B vssd1 vssd1 vccd1 vccd1 _1938_/Y sky130_fd_sc_hd__nand2_1
X_1869_ _1626_/Y _1762_/X _1867_/X _1868_/Y _1922_/B vssd1 vssd1 vccd1 vccd1 _2720_/B
+ sky130_fd_sc_hd__o221ai_4
Xhold820 _2975_/X vssd1 vssd1 vccd1 vccd1 _3650_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3608_ _3637_/CLK _3608_/D vssd1 vssd1 vccd1 vccd1 _3608_/Q sky130_fd_sc_hd__dfxtp_1
Xhold853 _2842_/X vssd1 vssd1 vccd1 vccd1 _3604_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold842 _3315_/Q vssd1 vssd1 vccd1 vccd1 hold842/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold831 _3727_/Q vssd1 vssd1 vccd1 vccd1 _3183_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold864 _3165_/X vssd1 vssd1 vccd1 vccd1 hold864/X sky130_fd_sc_hd__dlygate4sd3_1
X_3539_ _3539_/CLK _3539_/D vssd1 vssd1 vccd1 vccd1 _3539_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1805__A _2245_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold875 _3614_/Q vssd1 vssd1 vccd1 vccd1 _2892_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xhold897 _3174_/X vssd1 vssd1 vccd1 vccd1 _3722_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold886 _3175_/X vssd1 vssd1 vccd1 vccd1 hold886/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1913__B1 _2228_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2641__A1 _3193_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1827__S0 _1760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1715__A _2085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1904__B1 _2085_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2004__S0 _1954_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2632__A1 _3198_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2910_ _2876_/A _2908_/Y _2909_/Y _2948_/B _2883_/Y vssd1 vssd1 vccd1 vccd1 _2910_/Y
+ sky130_fd_sc_hd__o221ai_1
XANTENNA__2980__S _2987_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2841_ _3599_/Q _1696_/Y _2940_/B2 hold335/X _2825_/Y vssd1 vssd1 vccd1 vccd1 _2841_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_38_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2772_ _2707_/B _2707_/C _2789_/S vssd1 vssd1 vccd1 vccd1 _2775_/B sky130_fd_sc_hd__a21o_1
X_1723_ hold61/A _3744_/Q _1937_/S vssd1 vssd1 vccd1 vccd1 _1724_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_38_wb_clk_i clkbuf_3_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3721_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_41_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold105 _3417_/Q vssd1 vssd1 vccd1 vccd1 hold105/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold116 _2376_/X vssd1 vssd1 vccd1 vccd1 _3343_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 _2523_/X vssd1 vssd1 vccd1 vccd1 _3469_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold127 _3376_/Q vssd1 vssd1 vccd1 vccd1 hold127/X sky130_fd_sc_hd__dlygate4sd3_1
X_1654_ _2159_/B _1654_/B _2159_/D vssd1 vssd1 vccd1 vccd1 _1667_/A sky130_fd_sc_hd__and3_1
XFILLER_0_0_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold149 _3463_/Q vssd1 vssd1 vccd1 vccd1 hold149/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1625__A _2185_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3324_ _3344_/CLK _3324_/D vssd1 vssd1 vccd1 vccd1 _3324_/Q sky130_fd_sc_hd__dfxtp_1
X_3255_ _3739_/CLK _3255_/D vssd1 vssd1 vccd1 vccd1 _3255_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2206_ _2357_/A hold765/X _2209_/S vssd1 vssd1 vccd1 vccd1 _2206_/X sky130_fd_sc_hd__mux2_1
X_3186_ hold31/X _2353_/A _3191_/S vssd1 vssd1 vccd1 vccd1 hold32/A sky130_fd_sc_hd__mux2_1
X_2137_ _2137_/A _2137_/B vssd1 vssd1 vccd1 vccd1 _2138_/B sky130_fd_sc_hd__or2_1
X_2068_ _2495_/A _2068_/B vssd1 vssd1 vccd1 vccd1 _3350_/D sky130_fd_sc_hd__and2_1
XFILLER_0_88_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2387__A0 _3193_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold661 _3567_/Q vssd1 vssd1 vccd1 vccd1 hold661/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold672 _2606_/X vssd1 vssd1 vccd1 vccd1 _3540_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold650 _2417_/X vssd1 vssd1 vccd1 vccd1 _3384_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold683 _3544_/Q vssd1 vssd1 vccd1 vccd1 hold683/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold694 _2461_/X vssd1 vssd1 vccd1 vccd1 _3420_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout85_A _2093_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2085__B _2085_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2075__C1 _2495_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2614__A1 _2656_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2975__S _2987_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3040_ _3040_/A _3054_/A vssd1 vssd1 vccd1 vccd1 _3040_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_58_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1813__C1 _2022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2824_ _2825_/A _2874_/B vssd1 vssd1 vccd1 vccd1 _2824_/X sky130_fd_sc_hd__and2_2
XFILLER_0_5_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2908__A2 _2868_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2369__A0 _3196_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_15_wb_clk_i_A clkbuf_3_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_5_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2755_ _2803_/A _2755_/B _2755_/C vssd1 vssd1 vccd1 vccd1 _2755_/Y sky130_fd_sc_hd__nand3_1
X_1706_ _2153_/A _3059_/A vssd1 vssd1 vccd1 vccd1 _1707_/C sky130_fd_sc_hd__nand2_1
X_2686_ _2742_/C _2734_/B _2734_/C vssd1 vssd1 vccd1 vccd1 _2735_/A sky130_fd_sc_hd__a21oi_2
X_1637_ _3228_/Q _3227_/Q _3226_/Q vssd1 vssd1 vccd1 vccd1 _3081_/B sky130_fd_sc_hd__or3_2
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3307_ _3721_/CLK hold74/X vssd1 vssd1 vccd1 vccd1 hold73/A sky130_fd_sc_hd__dfxtp_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3238_ _3585_/CLK _3238_/D vssd1 vssd1 vccd1 vccd1 _3238_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3169_ _3169_/A _3181_/B vssd1 vssd1 vccd1 vccd1 _3169_/X sky130_fd_sc_hd__or2_1
XANTENNA_clkbuf_leaf_54_wb_clk_i_A clkbuf_leaf_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__2057__C1 _1979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout77 _2652_/A0 vssd1 vssd1 vccd1 vccd1 _2361_/A sky130_fd_sc_hd__buf_4
Xfanout99 _2961_/Y vssd1 vssd1 vccd1 vccd1 _2987_/S sky130_fd_sc_hd__buf_6
Xfanout88 _2091_/X vssd1 vssd1 vccd1 vccd1 _3194_/A0 sky130_fd_sc_hd__clkbuf_4
XANTENNA__1964__S _2085_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold480 _2265_/X vssd1 vssd1 vccd1 vccd1 _3290_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold491 _3549_/Q vssd1 vssd1 vccd1 vccd1 hold491/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2599__A0 _2655_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2063__A2 _2955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2540_ hold95/X _3197_/A0 _2541_/S vssd1 vssd1 vccd1 vccd1 hold96/A sky130_fd_sc_hd__mux2_1
X_2471_ _2363_/A hold251/X _2471_/S vssd1 vssd1 vccd1 vccd1 _2471_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_23_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2826__A1 hold918/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3023_ _3024_/A _3023_/B vssd1 vssd1 vccd1 vccd1 _3025_/B sky130_fd_sc_hd__or2_1
XANTENNA__2039__C1 _2495_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_53_wb_clk_i clkbuf_leaf_5_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3668_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_18_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout135_A _3346_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2807_ _2723_/Y _2802_/Y _2806_/X vssd1 vssd1 vccd1 vccd1 _2807_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_33_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2738_ _2738_/A _2738_/B vssd1 vssd1 vccd1 vccd1 _2738_/Y sky130_fd_sc_hd__nor2_1
X_2669_ _2669_/A _2669_/B _2669_/C vssd1 vssd1 vccd1 vccd1 _2811_/A sky130_fd_sc_hd__and3_2
XFILLER_0_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1868__A2 _2022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2817__A1 hold908/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2505__A0 _3197_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2269__C1 _3058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output29_A _3774_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1971_ _2022_/A _1971_/B _1971_/C vssd1 vssd1 vccd1 vccd1 _1971_/Y sky130_fd_sc_hd__nand3_1
X_3710_ _3714_/CLK _3710_/D vssd1 vssd1 vccd1 vccd1 _3710_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3641_ _3672_/CLK _3641_/D vssd1 vssd1 vccd1 vccd1 _3641_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3572_ _3575_/CLK _3572_/D vssd1 vssd1 vccd1 vccd1 _3572_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2523_ hold137/X _3201_/A1 _2527_/S vssd1 vssd1 vccd1 vccd1 _2523_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_11_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2454_ hold5/X _2650_/A0 _2457_/S vssd1 vssd1 vccd1 vccd1 hold6/A sky130_fd_sc_hd__mux2_1
XFILLER_0_11_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2385_ _2660_/A0 hold501/X _2385_/S vssd1 vssd1 vccd1 vccd1 _2385_/X sky130_fd_sc_hd__mux2_1
Xinput1 io_in[10] vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__buf_1
XANTENNA__1779__S _1937_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3006_ _3007_/A _3045_/D vssd1 vssd1 vccd1 vccd1 _3053_/C sky130_fd_sc_hd__nor2_1
XANTENNA__2275__A2 _2245_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1881__S1 _2245_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2170_ _3059_/A _1821_/X _2153_/A vssd1 vssd1 vccd1 vccd1 _2170_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_73_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2983__S _2987_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1954_ _3342_/Q _3300_/Q _1954_/S vssd1 vssd1 vccd1 vccd1 _1955_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1885_ _2245_/B _1885_/B vssd1 vssd1 vccd1 vccd1 _1885_/Y sky130_fd_sc_hd__nand2_1
X_3624_ _3674_/CLK _3624_/D vssd1 vssd1 vccd1 vccd1 _3624_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3555_ _3585_/CLK _3555_/D vssd1 vssd1 vccd1 vccd1 _3555_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3486_ _3539_/CLK _3486_/D vssd1 vssd1 vccd1 vccd1 _3486_/Q sky130_fd_sc_hd__dfxtp_1
X_2506_ _3198_/A0 hold663/X _2506_/S vssd1 vssd1 vccd1 vccd1 _2506_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1940__A1 _1889_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2437_ _3108_/A _2084_/A _2084_/B _2598_/A _2647_/B vssd1 vssd1 vccd1 vccd1 _2443_/S
+ sky130_fd_sc_hd__o311a_2
XFILLER_0_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2368_ _3195_/A0 hold777/X _2371_/S vssd1 vssd1 vccd1 vccd1 _2368_/X sky130_fd_sc_hd__mux2_1
X_2299_ _2301_/A _3227_/Q _3226_/Q _2302_/A vssd1 vssd1 vccd1 vccd1 _2300_/A sky130_fd_sc_hd__or4_1
XFILLER_0_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2956__A0 _2074_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1790__S0 _2000_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1845__S1 _2219_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1670_ _2885_/B _2960_/A vssd1 vssd1 vccd1 vccd1 _2083_/B sky130_fd_sc_hd__nand2_4
XFILLER_0_40_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1882__S _1988_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold309 _3392_/Q vssd1 vssd1 vccd1 vccd1 hold309/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2978__S _2987_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2175__A1 _3157_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3340_ _3581_/CLK _3340_/D vssd1 vssd1 vccd1 vccd1 _3340_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3271_ _3322_/CLK _3271_/D vssd1 vssd1 vccd1 vccd1 _3271_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1009 _1820_/X vssd1 vssd1 vccd1 vccd1 _3611_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2222_ _2355_/A hold279/X _2226_/S vssd1 vssd1 vccd1 vccd1 _2222_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1686__B1 _2961_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2153_ _2153_/A _2301_/C _3081_/B vssd1 vssd1 vccd1 vccd1 _2153_/Y sky130_fd_sc_hd__nor3_2
XFILLER_0_88_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2084_ _2084_/A _2084_/B vssd1 vssd1 vccd1 vccd1 _2245_/C sky130_fd_sc_hd__nor2_4
XFILLER_0_88_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2986_ hold335/X _2986_/A1 _2987_/S vssd1 vssd1 vccd1 vccd1 _2986_/X sky130_fd_sc_hd__mux2_1
X_1937_ _3470_/Q _3488_/Q _1937_/S vssd1 vssd1 vccd1 vccd1 _1938_/B sky130_fd_sc_hd__mux2_1
X_1868_ input6/X _2022_/A _1762_/X vssd1 vssd1 vccd1 vccd1 _1868_/Y sky130_fd_sc_hd__o21ai_2
Xhold821 _3699_/Q vssd1 vssd1 vccd1 vccd1 hold821/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold810 _3123_/X vssd1 vssd1 vccd1 vccd1 _3700_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3607_ _3670_/CLK _3607_/D vssd1 vssd1 vccd1 vccd1 _3607_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3538_ _3741_/CLK _3538_/D vssd1 vssd1 vccd1 vccd1 _3538_/Q sky130_fd_sc_hd__dfxtp_1
X_1799_ _3774_/A _2005_/S _2085_/C _1798_/Y vssd1 vssd1 vccd1 vccd1 _1799_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_12_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold854 _3619_/Q vssd1 vssd1 vccd1 vccd1 _2914_/A sky130_fd_sc_hd__buf_1
Xhold843 _2330_/X vssd1 vssd1 vccd1 vccd1 _3315_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold832 _3183_/Y vssd1 vssd1 vccd1 vccd1 hold832/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold876 _2890_/X vssd1 vssd1 vccd1 vccd1 _3614_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold898 _3703_/Q vssd1 vssd1 vccd1 vccd1 hold898/X sky130_fd_sc_hd__buf_1
Xhold865 _3166_/X vssd1 vssd1 vccd1 vccd1 _3718_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold887 _3176_/X vssd1 vssd1 vccd1 vccd1 _3723_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1913__A1 _2085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3469_ _3744_/CLK _3469_/D vssd1 vssd1 vccd1 vccd1 _3469_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_8_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3735_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__1827__S1 _1760_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1715__B _2228_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1904__A1 _3770_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2004__S1 _2014_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2840_ _3598_/Q _2871_/A _2839_/Y _2876_/B vssd1 vssd1 vccd1 vccd1 _2840_/X sky130_fd_sc_hd__o211a_1
X_2771_ _2771_/A _2771_/B vssd1 vssd1 vccd1 vccd1 _2773_/B sky130_fd_sc_hd__xnor2_1
X_1722_ _3502_/Q _3514_/Q _3526_/Q _3538_/Q _1937_/S _2245_/B vssd1 vssd1 vccd1 vccd1
+ _1722_/X sky130_fd_sc_hd__mux4_1
Xhold106 _2457_/X vssd1 vssd1 vccd1 vccd1 _3417_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1653_ _3628_/Q _3629_/Q _1653_/C _3627_/Q vssd1 vssd1 vccd1 vccd1 _2159_/D sky130_fd_sc_hd__or4b_2
Xhold117 _3386_/Q vssd1 vssd1 vccd1 vccd1 hold117/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold128 _2408_/X vssd1 vssd1 vccd1 vccd1 _3376_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold139 _3433_/Q vssd1 vssd1 vccd1 vccd1 hold139/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3323_ _3721_/CLK _3323_/D vssd1 vssd1 vccd1 vccd1 _3323_/Q sky130_fd_sc_hd__dfxtp_1
X_3254_ _3545_/CLK _3254_/D vssd1 vssd1 vccd1 vccd1 _3254_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2205_ _2355_/A hold697/X _2209_/S vssd1 vssd1 vccd1 vccd1 _2205_/X sky130_fd_sc_hd__mux2_1
X_3185_ _3192_/B _3185_/B vssd1 vssd1 vccd1 vccd1 _3191_/S sky130_fd_sc_hd__nor2_4
XANTENNA__1641__A _3045_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2136_ _3722_/Q _2155_/A _3723_/Q vssd1 vssd1 vccd1 vccd1 _2137_/B sky130_fd_sc_hd__a21oi_1
X_2067_ _2066_/X _2074_/A _2067_/S vssd1 vssd1 vccd1 vccd1 _2068_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_48_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_44_wb_clk_i_A clkbuf_3_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__1787__S _2244_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2472__A _3192_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2969_ hold297/X _3621_/Q _2999_/S vssd1 vssd1 vccd1 vccd1 _2969_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold640 _2395_/X vssd1 vssd1 vccd1 vccd1 _3365_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold662 _2637_/X vssd1 vssd1 vccd1 vccd1 _3567_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold651 _3488_/Q vssd1 vssd1 vccd1 vccd1 hold651/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold684 _2610_/X vssd1 vssd1 vccd1 vccd1 _3544_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold695 _3373_/Q vssd1 vssd1 vccd1 vccd1 hold695/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold673 _3218_/Q vssd1 vssd1 vccd1 vccd1 hold673/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout78_A _2097_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2647__A _2647_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2085__C _2085_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2378__A1 _2653_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1726__A _2245_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1984__S0 _2085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2550__A1 _2655_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1736__S0 _2000_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2838__C1 _2859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2823_ _2874_/B vssd1 vssd1 vccd1 vccd1 _2823_/Y sky130_fd_sc_hd__inv_2
X_2754_ _2754_/A _2754_/B vssd1 vssd1 vccd1 vccd1 _2756_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_83_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1705_ _3694_/Q _3693_/Q vssd1 vssd1 vccd1 vccd1 _1705_/X sky130_fd_sc_hd__or2_2
XFILLER_0_30_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2685_ _2720_/B _2720_/C _3594_/Q vssd1 vssd1 vccd1 vccd1 _2734_/C sky130_fd_sc_hd__a21bo_1
X_1636_ _3097_/B _3124_/A vssd1 vssd1 vccd1 vccd1 _3048_/B sky130_fd_sc_hd__or2_4
XANTENNA__2541__A1 _2660_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3306_ _3721_/CLK hold52/X vssd1 vssd1 vccd1 vccd1 hold51/A sky130_fd_sc_hd__dfxtp_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3237_ _3575_/CLK _3237_/D vssd1 vssd1 vccd1 vccd1 _3237_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_0_wb_clk_i_A clkbuf_leaf_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_3168_ hold927/X _3158_/Y _3167_/X _3172_/C1 vssd1 vssd1 vccd1 vccd1 _3168_/X sky130_fd_sc_hd__o211a_1
XANTENNA__2186__B _3192_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2119_ _2653_/A0 hold467/X _2119_/S vssd1 vssd1 vccd1 vccd1 _2119_/X sky130_fd_sc_hd__mux2_1
X_3099_ _2301_/A _3048_/B _3096_/C _3097_/X vssd1 vssd1 vccd1 vccd1 _3099_/X sky130_fd_sc_hd__o31a_1
XFILLER_0_49_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout89 _2091_/X vssd1 vssd1 vccd1 vccd1 _2656_/A0 sky130_fd_sc_hd__clkbuf_4
Xfanout78 _2097_/X vssd1 vssd1 vccd1 vccd1 _2652_/A0 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_17_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold470 _2398_/X vssd1 vssd1 vccd1 vccd1 _3368_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold481 _3452_/Q vssd1 vssd1 vccd1 vccd1 hold481/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold492 _2616_/X vssd1 vssd1 vccd1 vccd1 _3549_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2532__A1 _3203_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1718__S0 _1981_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2048__B1 _2867_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_300 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2470_ _2652_/A0 hold531/X _2471_/S vssd1 vssd1 vccd1 vccd1 _2470_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2986__S _2987_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2523__A1 _3201_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1890__S _2244_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2287__A0 _2361_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3022_ _3045_/B _3019_/Y _3080_/A vssd1 vssd1 vccd1 vccd1 _3023_/B sky130_fd_sc_hd__o21a_1
XANTENNA__2826__A2 _1696_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_83 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout128_A _1849_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2806_ _2082_/D _2802_/A _2759_/B _2851_/A vssd1 vssd1 vccd1 vccd1 _2806_/X sky130_fd_sc_hd__a2bb2o_1
X_2737_ _2740_/B _2736_/X _2789_/S vssd1 vssd1 vccd1 vccd1 _2738_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_22_wb_clk_i clkbuf_3_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3270_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2668_ _2669_/B _2669_/C vssd1 vssd1 vccd1 vccd1 _2871_/A sky130_fd_sc_hd__and2_4
XFILLER_0_14_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1619_ _2316_/A vssd1 vssd1 vccd1 vccd1 _2315_/A sky130_fd_sc_hd__inv_2
X_2599_ _2655_/A0 hold259/X _2604_/S vssd1 vssd1 vccd1 vccd1 _2599_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_1_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2450__A0 _3198_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2202__A0 _2660_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1970_ _2228_/A _1959_/X _1966_/X _1969_/Y vssd1 vssd1 vccd1 vccd1 _1971_/C sky130_fd_sc_hd__a31o_1
XFILLER_0_55_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2570__A _2570_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3640_ _3718_/CLK _3640_/D vssd1 vssd1 vccd1 vccd1 _3640_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2992__A1 _2480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3571_ _3585_/CLK _3571_/D vssd1 vssd1 vccd1 vccd1 _3571_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2522_ hold525/X _2353_/A _2527_/S vssd1 vssd1 vccd1 vccd1 _2522_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_87_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2453_ hold33/X _3201_/A1 _2457_/S vssd1 vssd1 vccd1 vccd1 hold34/A sky130_fd_sc_hd__mux2_1
X_2384_ _2659_/A0 hold509/X _2385_/S vssd1 vssd1 vccd1 vccd1 _2384_/X sky130_fd_sc_hd__mux2_1
Xinput2 io_in[11] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__buf_1
X_3005_ _3063_/B _3040_/A vssd1 vssd1 vccd1 vccd1 _3045_/D sky130_fd_sc_hd__nand2_2
XFILLER_0_36_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2275__A3 _2651_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2480__A _2480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3769_ _3769_/A vssd1 vssd1 vccd1 vccd1 _3769_/X sky130_fd_sc_hd__buf_1
XANTENNA__2499__A0 _2076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2974__A1 _3612_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1734__A _2006_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2549__B _2612_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1953_ _3294_/Q _3444_/Q _3578_/Q _3402_/Q _2005_/S _2014_/A vssd1 vssd1 vccd1 vccd1
+ _1953_/X sky130_fd_sc_hd__mux4_1
X_1884_ _3469_/Q _3487_/Q _1937_/S vssd1 vssd1 vccd1 vccd1 _1885_/B sky130_fd_sc_hd__mux2_1
XANTENNA__1768__A2 _2868_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3623_ _3714_/CLK _3623_/D vssd1 vssd1 vccd1 vccd1 _3623_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_24_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3554_ _3586_/CLK _3554_/D vssd1 vssd1 vccd1 vccd1 _3554_/Q sky130_fd_sc_hd__dfxtp_1
X_3485_ _3587_/CLK hold16/X vssd1 vssd1 vccd1 vccd1 hold15/A sky130_fd_sc_hd__dfxtp_1
X_2505_ _3197_/A0 hold487/X _2506_/S vssd1 vssd1 vccd1 vccd1 _2505_/X sky130_fd_sc_hd__mux2_1
X_2436_ hold573/X _2363_/A _2436_/S vssd1 vssd1 vccd1 vccd1 _2436_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2367_ _3194_/A0 hold323/X _2371_/S vssd1 vssd1 vccd1 vccd1 _2367_/X sky130_fd_sc_hd__mux2_1
X_2298_ _2298_/A vssd1 vssd1 vccd1 vccd1 _2298_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_78_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2653__A0 _2653_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2405__A0 _3197_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2184__A2 _3157_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1790__S1 _2219_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2947__A1 _1712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3270_ _3270_/CLK _3270_/D vssd1 vssd1 vccd1 vccd1 _3270_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2221_ _2648_/A0 hold195/X _2226_/S vssd1 vssd1 vccd1 vccd1 _2221_/X sky130_fd_sc_hd__mux2_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2152_ _3715_/Q _3703_/Q _2152_/S vssd1 vssd1 vccd1 vccd1 _2152_/X sky130_fd_sc_hd__mux2_1
X_2083_ _2854_/A _2083_/B _2083_/C vssd1 vssd1 vccd1 vccd1 _2083_/Y sky130_fd_sc_hd__nor3_1
XANTENNA__2635__A0 _2656_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_34_wb_clk_i_A clkbuf_3_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_8_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2985_ hold607/X _2985_/A1 _2987_/S vssd1 vssd1 vccd1 vccd1 _2985_/X sky130_fd_sc_hd__mux2_1
X_1936_ _2006_/A _1936_/B vssd1 vssd1 vccd1 vccd1 _1936_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_71_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1867_ _2022_/A _1867_/B _1867_/C vssd1 vssd1 vccd1 vccd1 _1867_/X sky130_fd_sc_hd__and3_1
X_1798_ _3333_/Q _2005_/S vssd1 vssd1 vccd1 vccd1 _1798_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_fanout110_A _2006_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3606_ _3670_/CLK _3606_/D vssd1 vssd1 vccd1 vccd1 _3606_/Q sky130_fd_sc_hd__dfxtp_1
Xhold811 _3701_/Q vssd1 vssd1 vccd1 vccd1 hold811/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold800 _2463_/X vssd1 vssd1 vccd1 vccd1 _3422_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3537_ _3561_/CLK _3537_/D vssd1 vssd1 vccd1 vccd1 _3537_/Q sky130_fd_sc_hd__dfxtp_1
Xhold822 _3121_/X vssd1 vssd1 vccd1 vccd1 _3699_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold855 _2917_/X vssd1 vssd1 vccd1 vccd1 _3619_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold844 _3617_/Q vssd1 vssd1 vccd1 vccd1 _2904_/A sky130_fd_sc_hd__buf_1
Xhold833 _3449_/Q vssd1 vssd1 vccd1 vccd1 hold833/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold888 _3624_/Q vssd1 vssd1 vccd1 vccd1 hold888/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold877 _3717_/Q vssd1 vssd1 vccd1 vccd1 _3163_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold866 _3724_/Q vssd1 vssd1 vccd1 vccd1 _3177_/A sky130_fd_sc_hd__dlygate4sd3_1
X_3468_ _3743_/CLK _3468_/D vssd1 vssd1 vccd1 vccd1 _3468_/Q sky130_fd_sc_hd__dfxtp_1
Xhold899 _3134_/X vssd1 vssd1 vccd1 vccd1 _3703_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3399_ _3744_/CLK _3399_/D vssd1 vssd1 vccd1 vccd1 _3399_/Q sky130_fd_sc_hd__dfxtp_1
X_2419_ hold117/X _3197_/A0 _2420_/S vssd1 vssd1 vccd1 vccd1 _2419_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_79_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2933__A _3103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3042__B1 _3055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2770_ _2680_/X _2754_/B _2759_/A vssd1 vssd1 vccd1 vccd1 _2771_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_79_25 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1721_ _1719_/X _1720_/X _1718_/X _1717_/X _2085_/A _2228_/C vssd1 vssd1 vccd1 vccd1
+ _1721_/X sky130_fd_sc_hd__mux4_1
Xhold107 _3548_/Q vssd1 vssd1 vccd1 vccd1 hold107/X sky130_fd_sc_hd__dlygate4sd3_1
X_1652_ _1713_/B _2034_/B _1663_/B vssd1 vssd1 vccd1 vccd1 _1654_/B sky130_fd_sc_hd__or3b_2
Xhold129 _3281_/Q vssd1 vssd1 vccd1 vccd1 hold129/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold118 _2419_/X vssd1 vssd1 vccd1 vccd1 _3386_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3322_ _3322_/CLK _3322_/D vssd1 vssd1 vccd1 vccd1 _3322_/Q sky130_fd_sc_hd__dfxtp_1
X_3253_ _3543_/CLK _3253_/D vssd1 vssd1 vccd1 vccd1 _3253_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_47_wb_clk_i clkbuf_3_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3674_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_3184_ _3080_/A hold832/X _2961_/A vssd1 vssd1 vccd1 vccd1 _3727_/D sky130_fd_sc_hd__a21oi_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2204_ _2648_/A0 hold787/X _2209_/S vssd1 vssd1 vccd1 vccd1 _2204_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1641__B _3048_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2135_ _3712_/Q _2135_/B _2135_/C vssd1 vssd1 vccd1 vccd1 _2166_/D sky130_fd_sc_hd__or3_1
XANTENNA__2608__A0 _3195_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2066_ _2480_/A _2036_/Y _2065_/X _2083_/B vssd1 vssd1 vccd1 vccd1 _2066_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_44_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2968_ hold199/X _2968_/A1 _2999_/S vssd1 vssd1 vccd1 vccd1 _2968_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_60_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1919_ _2022_/A _1915_/X _1917_/X _1918_/Y vssd1 vssd1 vccd1 vccd1 _1919_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_60_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2899_ _2876_/A _2895_/X _2898_/Y vssd1 vssd1 vccd1 vccd1 _2900_/B sky130_fd_sc_hd__o21ai_1
Xhold630 _2434_/X vssd1 vssd1 vccd1 vccd1 _3397_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold652 _2545_/X vssd1 vssd1 vccd1 vccd1 _3488_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold641 _3486_/Q vssd1 vssd1 vccd1 vccd1 hold641/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold663 _3455_/Q vssd1 vssd1 vccd1 vccd1 hold663/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold696 _2404_/X vssd1 vssd1 vccd1 vccd1 _3373_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold674 _2114_/X vssd1 vssd1 vccd1 vccd1 _3218_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold685 _3220_/Q vssd1 vssd1 vccd1 vccd1 hold685/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1832__A _2085_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2085__D _2480_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1984__S1 _2228_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1736__S1 _2219_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2066__A1 _2480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2822_ _2822_/A _2822_/B _2822_/C vssd1 vssd1 vccd1 vccd1 _2874_/B sky130_fd_sc_hd__and3_1
XFILLER_0_5_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2753_ _2734_/B _2736_/B _2742_/C vssd1 vssd1 vccd1 vccd1 _2754_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_81_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1704_ _3694_/Q _1704_/B vssd1 vssd1 vccd1 vccd1 _3768_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_30_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2684_ _2742_/C _2734_/B vssd1 vssd1 vccd1 vccd1 _2736_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1635_ _3097_/B _3124_/A vssd1 vssd1 vccd1 vccd1 _3096_/A sky130_fd_sc_hd__nor2_4
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3305_ _3308_/CLK hold56/X vssd1 vssd1 vccd1 vccd1 hold55/A sky130_fd_sc_hd__dfxtp_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3236_ _3585_/CLK _3236_/D vssd1 vssd1 vccd1 vccd1 _3236_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2829__B1 _2940_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3167_ _3719_/Q _3181_/B vssd1 vssd1 vccd1 vccd1 _3167_/X sky130_fd_sc_hd__or2_1
X_3098_ _2311_/C _3097_/X _3096_/X _2298_/Y vssd1 vssd1 vccd1 vccd1 _3100_/S sky130_fd_sc_hd__a211o_1
X_2118_ _2652_/A0 hold379/X _2119_/S vssd1 vssd1 vccd1 vccd1 _2118_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2057__A1 _2074_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2049_ _2228_/C _2036_/Y _2048_/X _2083_/B vssd1 vssd1 vccd1 vccd1 _2049_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_49_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout79 _3196_/A0 vssd1 vssd1 vccd1 vccd1 _2658_/A0 sky130_fd_sc_hd__buf_4
XFILLER_0_17_353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold460 _2213_/X vssd1 vssd1 vccd1 vccd1 _3250_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold471 _3434_/Q vssd1 vssd1 vccd1 vccd1 hold471/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout90_A _2091_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold482 _2503_/X vssd1 vssd1 vccd1 vccd1 _3452_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold493 _3338_/Q vssd1 vssd1 vccd1 vccd1 hold493/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1718__S1 _1981_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2296__A1 _2653_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3021_ _3183_/A _3183_/B vssd1 vssd1 vccd1 vccd1 _3080_/A sky130_fd_sc_hd__or2_2
XFILLER_0_25_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2805_ _2803_/A _2802_/Y _2800_/X _2790_/B _2790_/A vssd1 vssd1 vccd1 vccd1 _2805_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_0_41_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2736_ _2736_/A _2736_/B vssd1 vssd1 vccd1 vccd1 _2736_/X sky130_fd_sc_hd__xor2_1
X_2667_ hold215/X _2363_/A _2667_/S vssd1 vssd1 vccd1 vccd1 _2667_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1618_ _3059_/A vssd1 vssd1 vccd1 vccd1 _2301_/C sky130_fd_sc_hd__inv_2
X_2598_ _2598_/A _2598_/B vssd1 vssd1 vccd1 vccd1 _2604_/S sky130_fd_sc_hd__nand2_4
XANTENNA__3172__C1 _3172_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3219_ _3636_/CLK _3219_/D vssd1 vssd1 vccd1 vccd1 _3219_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3772__A _3772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold290 _2534_/X vssd1 vssd1 vccd1 vccd1 _3479_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2269__A1 _2022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2441__A1 _2651_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3570_ _3570_/CLK hold50/X vssd1 vssd1 vccd1 vccd1 hold49/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2521_ _2640_/A _3199_/B vssd1 vssd1 vccd1 vccd1 _2527_/S sky130_fd_sc_hd__nor2_2
XFILLER_0_23_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2452_ hold9/X _2648_/A0 _2457_/S vssd1 vssd1 vccd1 vccd1 hold10/A sky130_fd_sc_hd__mux2_1
XANTENNA__3154__C1 _3103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2383_ _2658_/A0 hold635/X _2385_/S vssd1 vssd1 vccd1 vccd1 _2383_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2901__C1 _3103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput3 io_in[12] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__buf_1
X_3004_ _3727_/Q _3045_/B vssd1 vssd1 vccd1 vccd1 _3004_/Y sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_3_4__f_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2432__A1 _3201_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout140_A _1988_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2480__B _3351_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3768_ _3768_/A vssd1 vssd1 vccd1 vccd1 _3768_/X sky130_fd_sc_hd__buf_1
X_2719_ _3628_/Q _2742_/B vssd1 vssd1 vccd1 vccd1 _2759_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_14_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3699_ _3714_/CLK _3699_/D vssd1 vssd1 vccd1 vccd1 _3699_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1840__A _2185_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1986__S _1988_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3767__A _3768_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2423__A1 _2656_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_24_wb_clk_i_A clkbuf_3_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__2111__A0 _2660_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2662__A1 _2353_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1952_ _1951_/X _1950_/X _1948_/X _1949_/X _2289_/A _2479_/B vssd1 vssd1 vccd1 vccd1
+ _1952_/X sky130_fd_sc_hd__mux4_1
XANTENNA__1848__S0 _2289_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1883_ _2006_/A _1883_/B vssd1 vssd1 vccd1 vccd1 _1883_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_22_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3622_ _3714_/CLK _3622_/D vssd1 vssd1 vccd1 vccd1 _3622_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_3_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3553_ _3583_/CLK _3553_/D vssd1 vssd1 vccd1 vccd1 _3553_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1925__B1 _2867_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3484_ _3496_/CLK hold96/X vssd1 vssd1 vccd1 vccd1 hold95/A sky130_fd_sc_hd__dfxtp_1
X_2504_ _3196_/A0 hold275/X _2506_/S vssd1 vssd1 vccd1 vccd1 _2504_/X sky130_fd_sc_hd__mux2_1
X_2435_ hold345/X _2361_/A _2436_/S vssd1 vssd1 vccd1 vccd1 _2435_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3127__C1 _3055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2366_ _3193_/A0 hold665/X _2371_/S vssd1 vssd1 vccd1 vccd1 _2366_/X sky130_fd_sc_hd__mux2_1
X_2297_ _3048_/B _3096_/B _3183_/B vssd1 vssd1 vccd1 vccd1 _2298_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_47_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1916__B1 _2195_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2341__A0 _2355_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2644__A1 _2658_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2580__A0 _3195_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2220_ _2237_/A _2647_/A vssd1 vssd1 vccd1 vccd1 _2226_/S sky130_fd_sc_hd__nand2_2
XANTENNA__2332__A0 _3193_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2151_ _3716_/Q _3704_/Q vssd1 vssd1 vccd1 vccd1 _2152_/S sky130_fd_sc_hd__xnor2_1
X_2082_ _3630_/Q _2961_/A _2082_/C _2082_/D vssd1 vssd1 vccd1 vccd1 _2083_/C sky130_fd_sc_hd__or4_1
XFILLER_0_48_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2399__A0 _2660_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2984_ hold327/X _2984_/A1 _2987_/S vssd1 vssd1 vccd1 vccd1 _2984_/X sky130_fd_sc_hd__mux2_1
X_1935_ hold69/A _3742_/Q _1937_/S vssd1 vssd1 vccd1 vccd1 _1936_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_8_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1866_ _2228_/A _1855_/X _1862_/X _1865_/Y vssd1 vssd1 vccd1 vccd1 _1867_/C sky130_fd_sc_hd__a31o_1
X_1797_ _2085_/C _1797_/B vssd1 vssd1 vccd1 vccd1 _1797_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_12_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold812 _3127_/X vssd1 vssd1 vccd1 vccd1 _3701_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3605_ _3662_/CLK _3605_/D vssd1 vssd1 vccd1 vccd1 _3605_/Q sky130_fd_sc_hd__dfxtp_1
Xhold801 _3675_/Q vssd1 vssd1 vccd1 vccd1 hold801/X sky130_fd_sc_hd__dlygate4sd3_1
X_3536_ _3539_/CLK _3536_/D vssd1 vssd1 vccd1 vccd1 _3536_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout103_A _1767_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold845 _2907_/X vssd1 vssd1 vccd1 vccd1 _3617_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold834 _2499_/X vssd1 vssd1 vccd1 vccd1 _3449_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold823 _3448_/Q vssd1 vssd1 vccd1 vccd1 hold823/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2571__A0 _2353_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold856 _3241_/Q vssd1 vssd1 vccd1 vccd1 _2054_/A sky130_fd_sc_hd__buf_1
Xhold889 _3153_/X vssd1 vssd1 vccd1 vccd1 hold889/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold878 _3163_/X vssd1 vssd1 vccd1 vccd1 hold878/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold867 _3177_/X vssd1 vssd1 vccd1 vccd1 hold867/X sky130_fd_sc_hd__dlygate4sd3_1
X_3467_ _3739_/CLK _3467_/D vssd1 vssd1 vccd1 vccd1 _3467_/Q sky130_fd_sc_hd__dfxtp_1
X_3398_ _3732_/CLK _3398_/D vssd1 vssd1 vccd1 vccd1 _3398_/Q sky130_fd_sc_hd__dfxtp_1
X_2418_ hold733/X _3196_/A0 _2420_/S vssd1 vssd1 vccd1 vccd1 _2418_/X sky130_fd_sc_hd__mux2_1
X_2349_ _2653_/A0 hold900/X _2349_/S vssd1 vssd1 vccd1 vccd1 _2349_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_74_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2865__A1 _3613_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3004__B _3045_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2617__A1 _2659_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2093__A2 _2084_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3020__A _3045_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_418 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1720_ _3434_/Q _3422_/Q _3410_/Q _3266_/Q _1981_/S0 _1981_/S1 vssd1 vssd1 vccd1
+ vccd1 _1720_/X sky130_fd_sc_hd__mux4_1
Xhold108 _2615_/X vssd1 vssd1 vccd1 vccd1 _3548_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1651_ _1713_/B _2669_/A _1663_/B vssd1 vssd1 vccd1 vccd1 _2878_/A sky130_fd_sc_hd__and3b_1
Xhold119 _3494_/Q vssd1 vssd1 vccd1 vccd1 hold119/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3321_ _3739_/CLK _3321_/D vssd1 vssd1 vccd1 vccd1 _3321_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3252_ _3545_/CLK _3252_/D vssd1 vssd1 vccd1 vccd1 _3252_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3183_ _3183_/A _3183_/B vssd1 vssd1 vccd1 vccd1 _3183_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__1922__B _1922_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2203_ _2237_/A _2570_/A vssd1 vssd1 vccd1 vccd1 _2209_/S sky130_fd_sc_hd__nand2_4
XFILLER_0_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2134_ _2135_/B _2135_/C _3712_/Q vssd1 vssd1 vccd1 vccd1 _2166_/C sky130_fd_sc_hd__o21ai_1
X_2065_ hold417/X _2731_/A2 _2034_/X _2868_/C vssd1 vssd1 vccd1 vccd1 _2065_/X sky130_fd_sc_hd__o22a_1
Xclkbuf_leaf_16_wb_clk_i clkbuf_3_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3586_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_63_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2967_ hold497/X _2967_/A1 _2999_/S vssd1 vssd1 vccd1 vccd1 _2967_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_44_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1918_ input7/X _2022_/A vssd1 vssd1 vccd1 vccd1 _1918_/Y sky130_fd_sc_hd__nor2_1
X_2898_ _2896_/Y _2904_/B _2935_/A vssd1 vssd1 vccd1 vccd1 _2898_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_44_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1849_ _3292_/Q _3442_/Q _3576_/Q _3400_/Q _1954_/S _1849_/S1 vssd1 vssd1 vccd1 vccd1
+ _1849_/X sky130_fd_sc_hd__mux4_1
Xhold620 _2642_/X vssd1 vssd1 vccd1 vccd1 _3571_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2544__A0 _3201_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold642 _2543_/X vssd1 vssd1 vccd1 vccd1 _3486_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold631 _3564_/Q vssd1 vssd1 vccd1 vccd1 hold631/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold653 _3372_/Q vssd1 vssd1 vccd1 vccd1 hold653/X sky130_fd_sc_hd__dlygate4sd3_1
X_3519_ _3543_/CLK _3519_/D vssd1 vssd1 vccd1 vccd1 _3519_/Q sky130_fd_sc_hd__dfxtp_1
Xhold664 _2506_/X vssd1 vssd1 vccd1 vccd1 _3455_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold675 _3339_/Q vssd1 vssd1 vccd1 vccd1 hold675/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold686 _2116_/X vssd1 vssd1 vccd1 vccd1 _3220_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold697 _3245_/Q vssd1 vssd1 vccd1 vccd1 hold697/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2847__A1 _2797_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2783__B1 _2731_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2821_ _1650_/A _2878_/A _2819_/A vssd1 vssd1 vccd1 vccd1 _2822_/C sky130_fd_sc_hd__o21ai_1
X_2752_ _2752_/A vssd1 vssd1 vccd1 vccd1 _2752_/Y sky130_fd_sc_hd__inv_2
X_1703_ _2054_/A _1700_/Y _1702_/X _2960_/A _2961_/A vssd1 vssd1 vccd1 vccd1 _1703_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_30_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2683_ _2682_/B _2682_/C _3595_/Q vssd1 vssd1 vccd1 vccd1 _2734_/B sky130_fd_sc_hd__a21o_1
X_1634_ _2305_/A _3687_/Q _3053_/B vssd1 vssd1 vccd1 vccd1 _3124_/A sky130_fd_sc_hd__or3_4
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3304_ _3666_/CLK _3304_/D vssd1 vssd1 vccd1 vccd1 _3304_/Q sky130_fd_sc_hd__dfxtp_1
X_3235_ _3575_/CLK _3235_/D vssd1 vssd1 vccd1 vccd1 _3235_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3166_ _3706_/Q _3158_/Y hold864/X _3166_/C1 vssd1 vssd1 vccd1 vccd1 _3166_/X sky130_fd_sc_hd__o211a_1
X_3097_ _3097_/A _3097_/B _3097_/C vssd1 vssd1 vccd1 vccd1 _3097_/X sky130_fd_sc_hd__or3_1
X_2117_ _2651_/A0 hold705/X _2119_/S vssd1 vssd1 vccd1 vccd1 _2117_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2057__A2 _2955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2048_ hold435/X _2731_/A2 _2867_/C _2034_/X vssd1 vssd1 vccd1 vccd1 _2048_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_76_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold461 _3237_/Q vssd1 vssd1 vccd1 vccd1 hold461/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2939__A _3103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold472 _2477_/X vssd1 vssd1 vccd1 vccd1 _3434_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold450 _2490_/X vssd1 vssd1 vccd1 vccd1 _3443_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold483 _3543_/Q vssd1 vssd1 vccd1 vccd1 hold483/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold494 _2370_/X vssd1 vssd1 vccd1 vccd1 _3338_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout83_A _2475_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2393__B _2647_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2048__A2 _2731_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1753__A _2085_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3020_ _3045_/B _3096_/A vssd1 vssd1 vccd1 vccd1 _3054_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_92_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2584__A _2647_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2804_ _2790_/A _2790_/B _2802_/Y _2789_/S _2803_/X vssd1 vssd1 vccd1 vccd1 _2804_/Y
+ sky130_fd_sc_hd__a221oi_1
XFILLER_0_73_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2747__A0 _2867_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2735_ _2735_/A _2735_/B vssd1 vssd1 vccd1 vccd1 _2740_/B sky130_fd_sc_hd__or2_1
X_2666_ hold163/X _2361_/A _2667_/S vssd1 vssd1 vccd1 vccd1 _2666_/X sky130_fd_sc_hd__mux2_1
X_1617_ _2182_/A vssd1 vssd1 vccd1 vccd1 _2301_/A sky130_fd_sc_hd__inv_2
X_2597_ hold271/X _2099_/X _2597_/S vssd1 vssd1 vccd1 vccd1 _2597_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_5_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_31_wb_clk_i clkbuf_3_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3728_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_3218_ _3666_/CLK _3218_/D vssd1 vssd1 vccd1 vccd1 _3218_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_hold1033_A _3349_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3149_ _3622_/Q _2886_/A _3137_/C vssd1 vssd1 vccd1 vccd1 _3149_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_92_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1789__A1 _2245_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1838__A _1889_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold280 _2222_/X vssd1 vssd1 vccd1 vccd1 _3257_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold291 _3337_/Q vssd1 vssd1 vccd1 vccd1 hold291/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2269__A2 _2245_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_14_wb_clk_i_A clkbuf_3_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_55_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2520_ hold529/X _3198_/A0 _2520_/S vssd1 vssd1 vccd1 vccd1 _2520_/X sky130_fd_sc_hd__mux2_1
X_2451_ _2647_/A _2528_/B vssd1 vssd1 vccd1 vccd1 _2457_/S sky130_fd_sc_hd__and2_2
XFILLER_0_23_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_53_wb_clk_i_A clkbuf_leaf_5_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_2382_ _3195_/A0 hold735/X _2385_/S vssd1 vssd1 vccd1 vccd1 _2382_/X sky130_fd_sc_hd__mux2_1
Xinput4 io_in[13] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__buf_1
X_3003_ _2961_/B hold939/X _2961_/A vssd1 vssd1 vccd1 vccd1 _3003_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_36_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2480__C _2480_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout133_A _1760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3767_ _3768_/A vssd1 vssd1 vccd1 vccd1 _3767_/X sky130_fd_sc_hd__buf_1
X_2718_ _2718_/A _2718_/B _2738_/A vssd1 vssd1 vccd1 vccd1 _2718_/X sky130_fd_sc_hd__or3b_1
X_3698_ _3714_/CLK _3698_/D vssd1 vssd1 vccd1 vccd1 _3698_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2649_ _2355_/A hold337/X _2653_/S vssd1 vssd1 vccd1 vccd1 _2649_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_77_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1824__C _3045_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2959__A0 _2050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2671__B _2868_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_452 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2187__A1 _2648_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output27_A _3773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1951_ _3548_/Q _3560_/Q _3572_/Q _3237_/Q _2289_/B _2289_/C vssd1 vssd1 vccd1 vccd1
+ _1951_/X sky130_fd_sc_hd__mux4_1
XANTENNA__1848__S1 _2479_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1882_ hold53/A _3741_/Q _1988_/S vssd1 vssd1 vccd1 vccd1 _1883_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_83_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3621_ _3674_/CLK _3621_/D vssd1 vssd1 vccd1 vccd1 _3621_/Q sky130_fd_sc_hd__dfxtp_2
X_3552_ _3587_/CLK _3552_/D vssd1 vssd1 vccd1 vccd1 _3552_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2503_ _2643_/A1 hold481/X _2506_/S vssd1 vssd1 vccd1 vccd1 _2503_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_3_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3483_ _3735_/CLK _3483_/D vssd1 vssd1 vccd1 vccd1 _3483_/Q sky130_fd_sc_hd__dfxtp_1
X_2434_ hold629/X _3203_/A1 _2436_/S vssd1 vssd1 vccd1 vccd1 _2434_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2102__A _3348_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2365_ _2365_/A _2598_/A vssd1 vssd1 vccd1 vccd1 _2371_/S sky130_fd_sc_hd__nand2_2
XANTENNA__1784__S0 _2244_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2296_ hold41/X _2653_/A0 _2296_/S vssd1 vssd1 vccd1 vccd1 hold42/A sky130_fd_sc_hd__mux2_1
XFILLER_0_78_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3108__A _3108_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2012__A _2289_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1775__S0 _2000_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2877__C1 _2960_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1851__A _2085_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2682__A _3595_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2150_ _2149_/B _2149_/C _3705_/Q vssd1 vssd1 vccd1 vccd1 _2150_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_17_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2081_ _3628_/Q _2741_/B vssd1 vssd1 vccd1 vccd1 _2082_/D sky130_fd_sc_hd__or2_2
XANTENNA__1843__B1 _2428_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2983_ hold647/X _2983_/A1 _2987_/S vssd1 vssd1 vccd1 vccd1 _2983_/X sky130_fd_sc_hd__mux2_1
X_1934_ _3500_/Q _3512_/Q _3524_/Q _3536_/Q _1937_/S _2245_/B vssd1 vssd1 vccd1 vccd1
+ _1934_/X sky130_fd_sc_hd__mux4_1
XANTENNA__1936__A _2006_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1865_ _2228_/A _1829_/X _2195_/B vssd1 vssd1 vccd1 vccd1 _1865_/Y sky130_fd_sc_hd__o21ai_1
X_1796_ hold57/A _3303_/Q _2005_/S vssd1 vssd1 vccd1 vccd1 _1797_/B sky130_fd_sc_hd__mux2_1
X_3604_ _3661_/CLK _3604_/D vssd1 vssd1 vccd1 vccd1 _3604_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold802 _3001_/X vssd1 vssd1 vccd1 vccd1 _3675_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3535_ _3561_/CLK _3535_/D vssd1 vssd1 vccd1 vccd1 _3535_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold813 _3702_/Q vssd1 vssd1 vccd1 vccd1 _3092_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold835 _3242_/Q vssd1 vssd1 vccd1 vccd1 _1824_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold846 _3690_/Q vssd1 vssd1 vccd1 vccd1 hold846/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold824 _2498_/X vssd1 vssd1 vccd1 vccd1 _3448_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2020__B1 _2195_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold857 _1703_/X vssd1 vssd1 vccd1 vccd1 _3241_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold879 _3164_/X vssd1 vssd1 vccd1 vccd1 _3717_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold868 _3178_/X vssd1 vssd1 vccd1 vccd1 _3724_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3466_ _3735_/CLK _3466_/D vssd1 vssd1 vccd1 vccd1 _3466_/Q sky130_fd_sc_hd__dfxtp_1
X_2417_ hold649/X _2475_/A1 _2420_/S vssd1 vssd1 vccd1 vccd1 _2417_/X sky130_fd_sc_hd__mux2_1
X_3397_ _3732_/CLK _3397_/D vssd1 vssd1 vccd1 vccd1 _3397_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2348_ _3108_/A _2348_/B vssd1 vssd1 vccd1 vccd1 _3326_/D sky130_fd_sc_hd__or2_1
X_2279_ _1716_/X _2480_/C _2653_/A0 _2278_/X _3058_/A vssd1 vssd1 vccd1 vccd1 _2279_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_39_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2562__A1 _2363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2219__B_N _2480_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1748__S0 _2085_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1650_ _1650_/A _1701_/A vssd1 vssd1 vccd1 vccd1 _2159_/B sky130_fd_sc_hd__nor2_1
Xhold109 _3501_/Q vssd1 vssd1 vccd1 vccd1 hold109/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3320_ _3738_/CLK _3320_/D vssd1 vssd1 vccd1 vccd1 _3320_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2553__A1 _3196_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3251_ _3543_/CLK _3251_/D vssd1 vssd1 vccd1 vccd1 _3251_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2202_ _2660_/A0 hold495/X _2202_/S vssd1 vssd1 vccd1 vccd1 _2202_/X sky130_fd_sc_hd__mux2_1
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3182_ hold948/X _3158_/Y _3181_/X _3086_/A vssd1 vssd1 vccd1 vccd1 _3182_/X sky130_fd_sc_hd__o211a_1
XANTENNA__2856__A2 _2940_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2133_ _3177_/A _2137_/A vssd1 vssd1 vccd1 vccd1 _2135_/C sky130_fd_sc_hd__nor2_1
X_2064_ _2071_/A _3045_/B _2071_/D vssd1 vssd1 vccd1 vccd1 _2067_/S sky130_fd_sc_hd__nor3_1
XANTENNA__2069__B1 _2868_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_56_wb_clk_i clkbuf_leaf_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3649_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_2966_ hold389/X _2966_/A1 _2992_/S vssd1 vssd1 vccd1 vccd1 _2966_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2241__A0 _2651_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2897_ _3137_/A _3615_/Q _3614_/Q vssd1 vssd1 vccd1 vccd1 _2904_/B sky130_fd_sc_hd__and3_1
X_1917_ _2228_/A _1906_/X _1913_/X _1916_/Y vssd1 vssd1 vccd1 vccd1 _1917_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_71_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1848_ _1847_/X _1846_/X _1844_/X _1845_/X _2289_/A _2479_/B vssd1 vssd1 vccd1 vccd1
+ _1848_/X sky130_fd_sc_hd__mux4_1
Xhold610 _2111_/X vssd1 vssd1 vccd1 vccd1 _3217_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold621 _3657_/Q vssd1 vssd1 vccd1 vccd1 hold621/X sky130_fd_sc_hd__dlygate4sd3_1
X_1779_ hold29/A _3745_/Q _1937_/S vssd1 vssd1 vccd1 vccd1 _1779_/X sky130_fd_sc_hd__mux2_1
Xhold643 _3505_/Q vssd1 vssd1 vccd1 vccd1 hold643/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold632 _2634_/X vssd1 vssd1 vccd1 vccd1 _3564_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold654 _2403_/X vssd1 vssd1 vccd1 vccd1 _3372_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3518_ _3545_/CLK _3518_/D vssd1 vssd1 vccd1 vccd1 _3518_/Q sky130_fd_sc_hd__dfxtp_1
Xhold676 _2371_/X vssd1 vssd1 vccd1 vccd1 _3339_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold665 _3334_/Q vssd1 vssd1 vccd1 vccd1 hold665/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold687 _3447_/Q vssd1 vssd1 vccd1 vccd1 hold687/X sky130_fd_sc_hd__dlygate4sd3_1
X_3449_ _3636_/CLK _3449_/D vssd1 vssd1 vccd1 vccd1 _3449_/Q sky130_fd_sc_hd__dfxtp_1
Xhold698 _2205_/X vssd1 vssd1 vccd1 vccd1 _3245_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2960__A _2960_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2783__A1 _2797_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2854__B _2854_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2471__A0 _2363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2820_ _1711_/X _2819_/X _1691_/B vssd1 vssd1 vccd1 vccd1 _2822_/B sky130_fd_sc_hd__o21a_1
XANTENNA__2223__A0 _2357_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2751_ _2867_/B hold923/X _2812_/S vssd1 vssd1 vccd1 vccd1 _2752_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_81_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1702_ _2819_/A _2054_/A _1701_/X _2876_/A vssd1 vssd1 vccd1 vccd1 _1702_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_5_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2682_ _3595_/Q _2682_/B _2682_/C vssd1 vssd1 vccd1 vccd1 _2742_/C sky130_fd_sc_hd__nand3_2
XFILLER_0_53_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1633_ _3037_/C _2310_/B vssd1 vssd1 vccd1 vccd1 _3097_/B sky130_fd_sc_hd__or2_2
XANTENNA__2526__A1 _2361_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_422 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3303_ _3728_/CLK _3303_/D vssd1 vssd1 vccd1 vccd1 _3303_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3234_ _3436_/CLK hold4/X vssd1 vssd1 vccd1 vccd1 hold3/A sky130_fd_sc_hd__dfxtp_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2829__A2 _1696_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3165_ _3165_/A _3181_/B vssd1 vssd1 vccd1 vccd1 _3165_/X sky130_fd_sc_hd__or2_1
X_3096_ _3096_/A _3096_/B _3096_/C vssd1 vssd1 vccd1 vccd1 _3096_/X sky130_fd_sc_hd__and3_1
X_2116_ _2650_/A0 hold685/X _2119_/S vssd1 vssd1 vccd1 vccd1 _2116_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2256__S _2259_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2047_ _2031_/Y _2045_/X _2046_/X _2495_/A vssd1 vssd1 vccd1 vccd1 _3348_/D sky130_fd_sc_hd__o211a_1
XANTENNA__2462__A0 _3196_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2214__A0 _2656_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2949_ hold888/X _2949_/A2 _2948_/Y _2947_/X _2885_/B vssd1 vssd1 vccd1 vccd1 _2949_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_72_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold440 _2546_/X vssd1 vssd1 vccd1 vccd1 _3489_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold462 _2199_/X vssd1 vssd1 vccd1 vccd1 _3237_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold451 _3576_/Q vssd1 vssd1 vccd1 vccd1 hold451/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3190__A1 _2361_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold484 _2609_/X vssd1 vssd1 vccd1 vccd1 _3543_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold495 _3240_/Q vssd1 vssd1 vccd1 vccd1 hold495/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold473 _3668_/Q vssd1 vssd1 vccd1 vccd1 hold473/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout76_A _2097_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2955__A _2955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2205__A0 _2355_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2508__A1 _2353_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_1_wb_clk_i clkbuf_leaf_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3655_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_clkbuf_leaf_43_wb_clk_i_A clkbuf_3_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_50_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2803_ _2803_/A _2803_/B _2803_/C vssd1 vssd1 vccd1 vccd1 _2803_/X sky130_fd_sc_hd__and3_1
XANTENNA__2747__A1 hold918/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2105__A _2570_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2734_ _2742_/C _2734_/B _2734_/C vssd1 vssd1 vccd1 vccd1 _2735_/B sky130_fd_sc_hd__and3_1
X_2665_ hold387/X _3203_/A1 _2667_/S vssd1 vssd1 vccd1 vccd1 _2665_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1944__A _2185_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2596_ hold173/X _2361_/A _2597_/S vssd1 vssd1 vccd1 vccd1 _2596_/X sky130_fd_sc_hd__mux2_1
X_1616_ _2797_/A vssd1 vssd1 vccd1 vccd1 _1616_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_1_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3217_ _3739_/CLK _3217_/D vssd1 vssd1 vccd1 vccd1 _3217_/Q sky130_fd_sc_hd__dfxtp_1
X_3148_ _2161_/A _3131_/X hold976/X _3103_/A vssd1 vssd1 vccd1 vccd1 _3148_/X sky130_fd_sc_hd__o211a_1
XANTENNA__2683__B1 _3595_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3079_ _3124_/A _3078_/Y _3076_/Y _3118_/A vssd1 vssd1 vccd1 vccd1 _3080_/C sky130_fd_sc_hd__a211o_1
XFILLER_0_64_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold270 _3200_/X vssd1 vssd1 vccd1 vccd1 _3740_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2910__A1 _2876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold281 _3418_/Q vssd1 vssd1 vccd1 vccd1 hold281/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold292 _2369_/X vssd1 vssd1 vccd1 vccd1 _3337_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2269__A3 _2648_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2977__A1 _3595_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2450_ _3198_/A0 hold719/X _2450_/S vssd1 vssd1 vccd1 vccd1 _2450_/X sky130_fd_sc_hd__mux2_1
X_2381_ _2656_/A0 hold463/X _2385_/S vssd1 vssd1 vccd1 vccd1 _2381_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2362__C1 _3172_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput5 io_in[14] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__buf_1
X_3002_ _2854_/B _1767_/Y _2885_/A vssd1 vssd1 vccd1 vccd1 _3002_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_36_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout126_A _1849_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1928__C1 _1979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2717_ _2717_/A _2717_/B vssd1 vssd1 vccd1 vccd1 _2718_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_42_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3697_ _3714_/CLK _3697_/D vssd1 vssd1 vccd1 vccd1 _3697_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2648_ _2648_/A0 hold451/X _2653_/S vssd1 vssd1 vccd1 vccd1 _2648_/X sky130_fd_sc_hd__mux2_1
X_2579_ _2656_/A0 hold715/X _2583_/S vssd1 vssd1 vccd1 vccd1 _2579_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_77_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2656__A0 _2656_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2408__A0 _2655_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2895__B1 _2867_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1950_ _3282_/Q _3354_/Q _3366_/Q _3378_/Q _2289_/B _2289_/C vssd1 vssd1 vccd1 vccd1
+ _1950_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_7_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1881_ _3499_/Q _3511_/Q _3523_/Q _3535_/Q _1988_/S _2245_/B vssd1 vssd1 vccd1 vccd1
+ _1881_/X sky130_fd_sc_hd__mux4_1
X_3620_ _3672_/CLK _3620_/D vssd1 vssd1 vccd1 vccd1 _3620_/Q sky130_fd_sc_hd__dfxtp_1
X_3551_ _3575_/CLK hold72/X vssd1 vssd1 vccd1 vccd1 hold71/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1925__A2 _2731_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2502_ _3194_/A0 hold603/X _2506_/S vssd1 vssd1 vccd1 vccd1 _2502_/X sky130_fd_sc_hd__mux2_1
X_3482_ _3558_/CLK _3482_/D vssd1 vssd1 vccd1 vccd1 _3482_/Q sky130_fd_sc_hd__dfxtp_1
X_2433_ hold761/X _2357_/A _2436_/S vssd1 vssd1 vccd1 vccd1 _2433_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2102__B _2244_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2364_ hold995/X _2351_/Y _2363_/X _3172_/C1 vssd1 vssd1 vccd1 vccd1 _3333_/D sky130_fd_sc_hd__o211a_1
XANTENNA__1784__S1 _2185_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2295_ hold89/X _2652_/A0 _2296_/S vssd1 vssd1 vccd1 vccd1 hold90/A sky130_fd_sc_hd__mux2_1
XANTENNA__2638__A0 _2097_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1669__A _2876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1775__S1 _2219_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2080_ _2080_/A _2080_/B _2080_/C vssd1 vssd1 vccd1 vccd1 _2084_/A sky130_fd_sc_hd__and3_4
XFILLER_0_17_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2096__A1 _2651_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2982_ hold621/X _2982_/A1 _2987_/S vssd1 vssd1 vccd1 vccd1 _2982_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_56_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1933_ _1931_/X _1932_/X _1930_/X _1929_/X _2085_/A _2228_/C vssd1 vssd1 vccd1 vccd1
+ _1933_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_33_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1864_ _2479_/A _1836_/X _1843_/X _1863_/Y vssd1 vssd1 vccd1 vccd1 _1867_/B sky130_fd_sc_hd__a31o_1
XFILLER_0_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3603_ _3661_/CLK _3603_/D vssd1 vssd1 vccd1 vccd1 _3603_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold803 _3696_/Q vssd1 vssd1 vccd1 vccd1 hold803/X sky130_fd_sc_hd__dlygate4sd3_1
X_1795_ _3297_/Q _3447_/Q _3581_/Q _3405_/Q _2005_/S _1849_/S1 vssd1 vssd1 vccd1 vccd1
+ _1795_/X sky130_fd_sc_hd__mux4_1
X_3534_ _3558_/CLK _3534_/D vssd1 vssd1 vccd1 vccd1 _3534_/Q sky130_fd_sc_hd__dfxtp_1
Xhold814 _3129_/X vssd1 vssd1 vccd1 vccd1 _3702_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold825 _3697_/Q vssd1 vssd1 vccd1 vccd1 hold825/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold836 _1695_/Y vssd1 vssd1 vccd1 vccd1 hold836/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold858 _3708_/Q vssd1 vssd1 vccd1 vccd1 hold858/X sky130_fd_sc_hd__buf_1
Xhold847 _3071_/X vssd1 vssd1 vccd1 vccd1 _3690_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold869 _3720_/Q vssd1 vssd1 vccd1 vccd1 _3169_/A sky130_fd_sc_hd__dlygate4sd3_1
X_3465_ _3735_/CLK _3465_/D vssd1 vssd1 vccd1 vccd1 _3465_/Q sky130_fd_sc_hd__dfxtp_1
X_2416_ hold103/X _3194_/A0 _2420_/S vssd1 vssd1 vccd1 vccd1 _2416_/X sky130_fd_sc_hd__mux2_1
X_3396_ _3592_/CLK _3396_/D vssd1 vssd1 vccd1 vccd1 _3396_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1671__B _1979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2259__S _2259_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2347_ _2652_/A0 hold895/X _2349_/S vssd1 vssd1 vccd1 vccd1 _2348_/B sky130_fd_sc_hd__mux2_1
X_2278_ _2278_/A _2278_/B vssd1 vssd1 vccd1 vccd1 _2278_/X sky130_fd_sc_hd__or2_1
XANTENNA__2007__B _2244_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1748__S1 _2014_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2250__A1 _2651_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1772__A _1979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3250_ _3587_/CLK _3250_/D vssd1 vssd1 vccd1 vccd1 _3250_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2201_ _2659_/A0 hold535/X _2202_/S vssd1 vssd1 vccd1 vccd1 _2201_/X sky130_fd_sc_hd__mux2_1
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3181_ _3726_/Q _3181_/B vssd1 vssd1 vccd1 vccd1 _3181_/X sky130_fd_sc_hd__or2_1
X_2132_ _3726_/Q _3713_/Q _2132_/C _3714_/Q vssd1 vssd1 vccd1 vccd1 _2132_/X sky130_fd_sc_hd__or4b_1
X_2063_ _2050_/A _2955_/A _2076_/C hold973/X _1979_/A vssd1 vssd1 vccd1 vccd1 _2063_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_48_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2965_ hold571/X _2965_/A1 _2999_/S vssd1 vssd1 vccd1 vccd1 _2965_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_44_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2896_ _3615_/Q _3614_/Q _3137_/A vssd1 vssd1 vccd1 vccd1 _2896_/Y sky130_fd_sc_hd__a21oi_1
X_1916_ _2228_/A _1880_/X _2195_/B vssd1 vssd1 vccd1 vccd1 _1916_/Y sky130_fd_sc_hd__o21ai_1
X_1847_ hold47/A hold63/A hold49/A _3235_/Q _2289_/B _2289_/C vssd1 vssd1 vccd1 vccd1
+ _1847_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_44_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_25_wb_clk_i clkbuf_3_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3741_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold611 _3536_/Q vssd1 vssd1 vccd1 vccd1 hold611/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold600 _2638_/X vssd1 vssd1 vccd1 vccd1 _3568_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_71_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3517_ _3543_/CLK _3517_/D vssd1 vssd1 vccd1 vccd1 _3517_/Q sky130_fd_sc_hd__dfxtp_1
Xhold644 _2565_/X vssd1 vssd1 vccd1 vccd1 _3505_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1778_ _3503_/Q _3515_/Q _3527_/Q _3539_/Q _1988_/S _2245_/B vssd1 vssd1 vccd1 vccd1
+ _1778_/X sky130_fd_sc_hd__mux4_1
Xhold633 _3303_/Q vssd1 vssd1 vccd1 vccd1 hold633/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold622 _2982_/X vssd1 vssd1 vccd1 vccd1 _3657_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold655 _3381_/Q vssd1 vssd1 vccd1 vccd1 hold655/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold677 _3742_/Q vssd1 vssd1 vccd1 vccd1 hold677/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold666 _2366_/X vssd1 vssd1 vccd1 vccd1 _3334_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold688 _2494_/X vssd1 vssd1 vccd1 vccd1 _3447_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold699 _3272_/Q vssd1 vssd1 vccd1 vccd1 hold699/X sky130_fd_sc_hd__dlygate4sd3_1
X_3448_ _3636_/CLK _3448_/D vssd1 vssd1 vccd1 vccd1 _3448_/Q sky130_fd_sc_hd__dfxtp_1
X_3379_ _3585_/CLK _3379_/D vssd1 vssd1 vccd1 vccd1 _3379_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1857__A _2289_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_33_wb_clk_i_A clkbuf_3_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_85_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2750_ hold918/X _2730_/Y _2748_/X _2749_/X _2859_/A vssd1 vssd1 vccd1 vccd1 _2750_/X
+ sky130_fd_sc_hd__o221a_1
X_1701_ _1701_/A _3130_/A vssd1 vssd1 vccd1 vccd1 _1701_/X sky130_fd_sc_hd__or2_1
XFILLER_0_30_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2681_ _3596_/Q _2867_/B vssd1 vssd1 vccd1 vccd1 _2754_/A sky130_fd_sc_hd__xnor2_4
X_1632_ _3063_/B _3682_/Q vssd1 vssd1 vccd1 vccd1 _2310_/B sky130_fd_sc_hd__or2_2
XFILLER_0_1_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2598__A _2598_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3302_ _3344_/CLK _3302_/D vssd1 vssd1 vccd1 vccd1 _3302_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3233_ _3743_/CLK _3233_/D vssd1 vssd1 vccd1 vccd1 _3233_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3164_ _3705_/Q _3158_/Y hold878/X _3166_/C1 vssd1 vssd1 vccd1 vccd1 _3164_/X sky130_fd_sc_hd__o211a_1
X_3095_ _3108_/A _3095_/B vssd1 vssd1 vccd1 vccd1 _3692_/D sky130_fd_sc_hd__nor2_1
X_2115_ _2355_/A hold365/X _2119_/S vssd1 vssd1 vccd1 vccd1 _2115_/X sky130_fd_sc_hd__mux2_1
X_2046_ _2046_/A _2050_/B vssd1 vssd1 vccd1 vccd1 _2046_/X sky130_fd_sc_hd__or2_1
XFILLER_0_49_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1896__S0 _2000_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout156_A _3172_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2948_ _2948_/A _2948_/B vssd1 vssd1 vccd1 vccd1 _2948_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_17_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2879_ _3613_/Q _3630_/Q vssd1 vssd1 vccd1 vccd1 _2879_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_32_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold463 _3353_/Q vssd1 vssd1 vccd1 vccd1 hold463/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold430 _2576_/X vssd1 vssd1 vccd1 vccd1 _3515_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold441 _3445_/Q vssd1 vssd1 vccd1 vccd1 hold441/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold452 _2648_/X vssd1 vssd1 vccd1 vccd1 _3576_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold496 _2202_/X vssd1 vssd1 vccd1 vccd1 _3240_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2922__C1 _3103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold474 _2993_/X vssd1 vssd1 vccd1 vccd1 _3668_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold485 _3465_/Q vssd1 vssd1 vccd1 vccd1 hold485/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2453__A1 _3201_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2690__B _2867_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2245__D_N _1937_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1878__S0 _1981_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2802_ _2802_/A _2851_/B vssd1 vssd1 vccd1 vccd1 _2802_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_41_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2733_ hold908/X _2730_/Y _2732_/X _2729_/X _2859_/A vssd1 vssd1 vccd1 vccd1 _2733_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_26_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2664_ hold203/X _2357_/A _2667_/S vssd1 vssd1 vccd1 vccd1 _2664_/X sky130_fd_sc_hd__mux2_1
X_2595_ hold43/X _3203_/A1 _2597_/S vssd1 vssd1 vccd1 vccd1 hold44/A sky130_fd_sc_hd__mux2_1
X_1615_ _2034_/B vssd1 vssd1 vccd1 vccd1 _2669_/A sky130_fd_sc_hd__inv_2
XFILLER_0_1_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1802__S0 _2085_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2380__A0 _2089_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3216_ _3738_/CLK _3216_/D vssd1 vssd1 vccd1 vccd1 _3216_/Q sky130_fd_sc_hd__dfxtp_1
X_3147_ _2924_/A _2886_/A _3137_/C vssd1 vssd1 vccd1 vccd1 _3147_/X sky130_fd_sc_hd__a21o_1
X_3078_ _2305_/A _3077_/X _3037_/D vssd1 vssd1 vccd1 vccd1 _3078_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_49_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2435__A1 _2361_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2029_ _3103_/A _2029_/B vssd1 vssd1 vccd1 vccd1 _3609_/D sky130_fd_sc_hd__and2_1
XFILLER_0_92_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_40_wb_clk_i clkbuf_3_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3724_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_60_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3148__C1 _3103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold271 _3533_/Q vssd1 vssd1 vccd1 vccd1 hold271/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold260 _2599_/X vssd1 vssd1 vccd1 vccd1 _3534_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2371__A0 _3198_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold293 _3363_/Q vssd1 vssd1 vccd1 vccd1 hold293/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 _2459_/X vssd1 vssd1 vccd1 vccd1 _3418_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2426__A1 _2659_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2380_ _2089_/X hold747/X _2385_/S vssd1 vssd1 vccd1 vccd1 _2380_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2876__A _2876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2114__A0 _2648_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput6 io_in[15] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__buf_1
XANTENNA__2665__A1 _3203_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3001_ hold801/X _3000_/X _2961_/B _3166_/C1 vssd1 vssd1 vccd1 vccd1 _3001_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_86_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2417__A1 _2475_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1955__A _2006_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3696_ _3702_/CLK _3696_/D vssd1 vssd1 vccd1 vccd1 _3696_/Q sky130_fd_sc_hd__dfxtp_1
X_2716_ _3612_/Q _2716_/B vssd1 vssd1 vccd1 vccd1 _2738_/A sky130_fd_sc_hd__nand2_2
X_2647_ _2647_/A _2647_/B vssd1 vssd1 vccd1 vccd1 _2653_/S sky130_fd_sc_hd__nand2_4
XFILLER_0_65_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2578_ _2655_/A0 hold723/X _2583_/S vssd1 vssd1 vccd1 vccd1 _2578_/X sky130_fd_sc_hd__mux2_1
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1804__S _1937_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1880_ _1878_/X _1879_/X _1877_/X _1876_/X _2085_/A _2228_/C vssd1 vssd1 vccd1 vccd1
+ _1880_/X sky130_fd_sc_hd__mux4_1
X_3550_ _3561_/CLK hold8/X vssd1 vssd1 vccd1 vccd1 hold7/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__2583__A0 _2660_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2501_ _2655_/A0 hold597/X _2506_/S vssd1 vssd1 vccd1 vccd1 _2501_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_11_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3481_ _3735_/CLK hold68/X vssd1 vssd1 vccd1 vccd1 hold67/A sky130_fd_sc_hd__dfxtp_1
X_2432_ hold347/X _3201_/A1 _2436_/S vssd1 vssd1 vccd1 vccd1 _2432_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2335__A0 _3196_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2363_ _2363_/A _2363_/B vssd1 vssd1 vccd1 vccd1 _2363_/X sky130_fd_sc_hd__or2_1
X_2294_ hold73/X _2651_/A0 _2296_/S vssd1 vssd1 vccd1 vccd1 hold74/A sky130_fd_sc_hd__mux2_1
XFILLER_0_63_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2271__C1 _3058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1685__A _2885_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2574__A0 _3203_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3679_ _3727_/CLK _3679_/D vssd1 vssd1 vccd1 vccd1 _3679_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2877__A1 _2876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2565__A0 _2656_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2203__B _2570_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2981_ hold759/X _3599_/Q _2987_/S vssd1 vssd1 vccd1 vccd1 _2981_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_33_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1932_ _3432_/Q _3420_/Q _3408_/Q _3264_/Q _1760_/A _1760_/B vssd1 vssd1 vccd1 vccd1
+ _1932_/X sky130_fd_sc_hd__mux4_1
X_1863_ _2479_/A _1848_/X _2228_/B vssd1 vssd1 vccd1 vccd1 _1863_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_16_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3602_ _3661_/CLK _3602_/D vssd1 vssd1 vccd1 vccd1 _3602_/Q sky130_fd_sc_hd__dfxtp_1
X_1794_ _1793_/X _1792_/X _1790_/X _1791_/X _2289_/A _2479_/B vssd1 vssd1 vccd1 vccd1
+ _1794_/X sky130_fd_sc_hd__mux4_1
X_3533_ _3745_/CLK _3533_/D vssd1 vssd1 vccd1 vccd1 _3533_/Q sky130_fd_sc_hd__dfxtp_1
Xhold804 _3111_/X vssd1 vssd1 vccd1 vccd1 _3696_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold826 _3114_/X vssd1 vssd1 vccd1 vccd1 _3697_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold837 _1699_/Y vssd1 vssd1 vccd1 vccd1 _3242_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold815 _3635_/Q vssd1 vssd1 vccd1 vccd1 hold815/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2113__B _2619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3464_ _3496_/CLK _3464_/D vssd1 vssd1 vccd1 vccd1 _3464_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold859 _3144_/X vssd1 vssd1 vccd1 vccd1 _3708_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold848 _3616_/Q vssd1 vssd1 vccd1 vccd1 _3137_/A sky130_fd_sc_hd__buf_1
X_2415_ hold169/X _3193_/A0 _2420_/S vssd1 vssd1 vccd1 vccd1 _2415_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_58_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3395_ _3733_/CLK _3395_/D vssd1 vssd1 vccd1 vccd1 _3395_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2346_ _3108_/A _2346_/B vssd1 vssd1 vccd1 vccd1 _3325_/D sky130_fd_sc_hd__or2_1
X_2277_ _1716_/X _2245_/C _2652_/A0 _2276_/X _3058_/A vssd1 vssd1 vccd1 vccd1 _2277_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_74_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2547__A0 _2361_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_23_wb_clk_i_A clkbuf_3_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__1770__A1 _2854_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2200_ _2658_/A0 hold539/X _2202_/S vssd1 vssd1 vccd1 vccd1 _2200_/X sky130_fd_sc_hd__mux2_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3180_ hold838/X _3158_/Y _3179_/X _3058_/A vssd1 vssd1 vccd1 vccd1 _3180_/X sky130_fd_sc_hd__o211a_1
X_2131_ hold838/X _2126_/Y _2130_/X vssd1 vssd1 vccd1 vccd1 _2131_/X sky130_fd_sc_hd__a21bo_1
X_2062_ _2854_/A _2062_/B vssd1 vssd1 vccd1 vccd1 _2062_/X sky130_fd_sc_hd__or2_1
XANTENNA__2069__A2 _2731_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1816__A2 _1922_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2964_ hold595/X _2964_/A1 _2992_/S vssd1 vssd1 vccd1 vccd1 _2964_/X sky130_fd_sc_hd__mux2_1
X_1915_ _2479_/A _1887_/X _1894_/X _1914_/Y vssd1 vssd1 vccd1 vccd1 _1915_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_84_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2895_ hold595/X _1767_/Y _2867_/B _2819_/A vssd1 vssd1 vccd1 vccd1 _2895_/X sky130_fd_sc_hd__o22a_1
X_1846_ _3280_/Q _3352_/Q _3364_/Q _3376_/Q _2289_/B _2289_/C vssd1 vssd1 vccd1 vccd1
+ _1846_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold612 _2601_/X vssd1 vssd1 vccd1 vccd1 _3536_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold601 _3235_/Q vssd1 vssd1 vccd1 vccd1 hold601/X sky130_fd_sc_hd__dlygate4sd3_1
X_1777_ _1775_/X _1776_/X _1774_/X _1773_/X _2085_/A _2228_/C vssd1 vssd1 vccd1 vccd1
+ _1777_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_12_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3516_ _3739_/CLK _3516_/D vssd1 vssd1 vccd1 vccd1 _3516_/Q sky130_fd_sc_hd__dfxtp_1
Xhold634 _2288_/X vssd1 vssd1 vccd1 vccd1 _3303_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1963__A _2014_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold645 _3289_/Q vssd1 vssd1 vccd1 vccd1 hold645/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold623 _3316_/Q vssd1 vssd1 vccd1 vccd1 hold623/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold667 _3285_/Q vssd1 vssd1 vccd1 vccd1 hold667/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold656 _2413_/X vssd1 vssd1 vccd1 vccd1 _3381_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold678 _3202_/X vssd1 vssd1 vccd1 vccd1 _3742_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold689 _3267_/Q vssd1 vssd1 vccd1 vccd1 hold689/X sky130_fd_sc_hd__dlygate4sd3_1
X_3447_ _3447_/CLK _3447_/D vssd1 vssd1 vccd1 vccd1 _3447_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3378_ _3586_/CLK _3378_/D vssd1 vssd1 vccd1 vccd1 _3378_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2329_ _2308_/Y _2328_/X _2318_/B vssd1 vssd1 vccd1 vccd1 _2329_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_39_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2768__A0 _2867_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1991__A1 _1889_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3193__A0 _3193_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1700_ _2876_/A _1690_/B _1680_/X vssd1 vssd1 vccd1 vccd1 _1700_/Y sky130_fd_sc_hd__o21bai_1
X_2680_ _3596_/Q _2867_/B vssd1 vssd1 vccd1 vccd1 _2680_/X sky130_fd_sc_hd__or2_1
XANTENNA__2879__A _3613_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1631_ _2309_/A _3045_/A vssd1 vssd1 vccd1 vccd1 _3037_/C sky130_fd_sc_hd__or2_2
XFILLER_0_30_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3184__B1 _2961_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3301_ _3344_/CLK _3301_/D vssd1 vssd1 vccd1 vccd1 _3301_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3232_ _3322_/CLK _3232_/D vssd1 vssd1 vccd1 vccd1 _3232_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3163_ _3163_/A _3181_/B vssd1 vssd1 vccd1 vccd1 _3163_/X sky130_fd_sc_hd__or2_1
X_2114_ _2648_/A0 hold673/X _2119_/S vssd1 vssd1 vccd1 vccd1 _2114_/X sky130_fd_sc_hd__mux2_1
X_3094_ _1600_/Y _3093_/X _3094_/S vssd1 vssd1 vccd1 vccd1 _3094_/X sky130_fd_sc_hd__mux2_1
X_2045_ _2085_/A _2036_/Y _2044_/X _2083_/B vssd1 vssd1 vccd1 vccd1 _2045_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1896__S1 _2219_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout149_A _2859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2947_ _1712_/A _2999_/A1 hold349/X _1766_/Y vssd1 vssd1 vccd1 vccd1 _2947_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_17_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2878_ _2878_/A _2878_/B _2878_/C vssd1 vssd1 vccd1 vccd1 _3130_/B sky130_fd_sc_hd__or3_2
XFILLER_0_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1973__A1 input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold420 _2643_/X vssd1 vssd1 vccd1 vccd1 _3572_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1829_ _1827_/X _1828_/X _1826_/X _1825_/X _2085_/A _2228_/C vssd1 vssd1 vccd1 vccd1
+ _1829_/X sky130_fd_sc_hd__mux4_1
Xhold453 _3508_/Q vssd1 vssd1 vccd1 vccd1 hold453/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold431 _3545_/Q vssd1 vssd1 vccd1 vccd1 hold431/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold442 _2492_/X vssd1 vssd1 vccd1 vccd1 _3445_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold464 _2381_/X vssd1 vssd1 vccd1 vccd1 _3353_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold475 _3366_/Q vssd1 vssd1 vccd1 vccd1 hold475/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold486 _2518_/X vssd1 vssd1 vccd1 vccd1 _3465_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold497 _3642_/Q vssd1 vssd1 vccd1 vccd1 hold497/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2029__A _3103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1878__S1 _1981_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2801_ _2675_/X _2788_/B _2677_/B vssd1 vssd1 vccd1 vccd1 _2851_/B sky130_fd_sc_hd__o21a_1
X_2732_ _2797_/A hold407/X _2731_/X vssd1 vssd1 vccd1 vccd1 _2732_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_54_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2663_ hold153/X _3201_/A1 _2667_/S vssd1 vssd1 vccd1 vccd1 _2663_/X sky130_fd_sc_hd__mux2_1
X_2594_ hold191/X _2650_/A0 _2597_/S vssd1 vssd1 vccd1 vccd1 _2594_/X sky130_fd_sc_hd__mux2_1
X_1614_ _2717_/B vssd1 vssd1 vccd1 vccd1 _2741_/A sky130_fd_sc_hd__inv_2
XANTENNA__1802__S1 _2014_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3215_ _3737_/CLK _3215_/D vssd1 vssd1 vccd1 vccd1 _3215_/Q sky130_fd_sc_hd__dfxtp_1
X_3146_ hold914/X _3131_/X _3145_/X _3166_/C1 vssd1 vssd1 vccd1 vccd1 _3146_/X sky130_fd_sc_hd__o211a_1
X_3077_ _3687_/Q _3686_/Q _3007_/A vssd1 vssd1 vccd1 vccd1 _3077_/X sky130_fd_sc_hd__or3b_1
XFILLER_0_89_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2028_ _2050_/A _2027_/X _2028_/S vssd1 vssd1 vccd1 vccd1 _2029_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_49_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold261 _3560_/Q vssd1 vssd1 vccd1 vccd1 hold261/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold250 _2962_/X vssd1 vssd1 vccd1 vccd1 _3637_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold272 _2597_/X vssd1 vssd1 vccd1 vccd1 _3533_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold283 _3461_/Q vssd1 vssd1 vccd1 vccd1 hold283/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_3_1__f_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold294 _2392_/X vssd1 vssd1 vccd1 vccd1 _3363_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout81_A _2651_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1870__B _1922_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output62_A _3676_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput7 io_in[16] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__buf_1
X_3000_ _3689_/Q _3058_/B vssd1 vssd1 vccd1 vccd1 _3000_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_86_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1720__S0 _1981_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1928__A1 _2076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3695_ _3695_/CLK _3695_/D vssd1 vssd1 vccd1 vccd1 _3695_/Q sky130_fd_sc_hd__dfxtp_1
X_2715_ _3612_/Q _2716_/B vssd1 vssd1 vccd1 vccd1 _2718_/A sky130_fd_sc_hd__nor2_1
X_2646_ hold299/X _2660_/A0 _2646_/S vssd1 vssd1 vccd1 vccd1 _2646_/X sky130_fd_sc_hd__mux2_1
X_2577_ _2654_/A _2647_/A vssd1 vssd1 vccd1 vccd1 _2583_/S sky130_fd_sc_hd__nand2_4
XANTENNA__1971__A _2022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3129_ _3092_/A _3120_/A _3128_/X _3055_/A vssd1 vssd1 vccd1 vccd1 _3129_/X sky130_fd_sc_hd__o211a_1
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1919__A1 _2022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2592__A1 _2353_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1778__S0 _1988_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2895__A2 _1767_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3057__C1 _3108_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2280__B1 _2480_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2500_ _2619_/A _2500_/B vssd1 vssd1 vccd1 vccd1 _2506_/S sky130_fd_sc_hd__nand2_4
X_3480_ _3496_/CLK _3480_/D vssd1 vssd1 vccd1 vccd1 _3480_/Q sky130_fd_sc_hd__dfxtp_1
X_2431_ hold741/X _2353_/A _2436_/S vssd1 vssd1 vccd1 vccd1 _2431_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_11_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2362_ hold962/X _2351_/Y _2361_/X _3172_/C1 vssd1 vssd1 vccd1 vccd1 _3332_/D sky130_fd_sc_hd__o211a_1
X_2293_ hold51/X _2650_/A0 _2296_/S vssd1 vssd1 vccd1 vccd1 hold52/A sky130_fd_sc_hd__mux2_1
XFILLER_0_47_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_19_wb_clk_i clkbuf_3_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3575_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_fanout131_A _1849_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_13_wb_clk_i_A clkbuf_3_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_88_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3678_ _3727_/CLK _3678_/D vssd1 vssd1 vccd1 vccd1 _3678_/Q sky130_fd_sc_hd__dfxtp_1
X_2629_ hold261/X _2643_/A1 _2632_/S vssd1 vssd1 vccd1 vccd1 _2629_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2797__A _2797_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1932__S0 _1760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_52_wb_clk_i_A clkbuf_leaf_5_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_77_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1999__S0 _2000_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2500__A _2619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output25_A _3772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2980_ hold565/X _3598_/Q _2987_/S vssd1 vssd1 vccd1 vccd1 _2980_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_56_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1931_ _3494_/Q _3482_/Q _3464_/Q _3452_/Q _1760_/A _1760_/B vssd1 vssd1 vccd1 vccd1
+ _1931_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_56_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1862_ _2289_/A _1859_/Y _1861_/Y _2228_/C _1857_/Y vssd1 vssd1 vccd1 vccd1 _1862_/X
+ sky130_fd_sc_hd__a311o_1
Xinput10 io_in[19] vssd1 vssd1 vccd1 vccd1 input10/X sky130_fd_sc_hd__buf_1
X_3601_ _3661_/CLK _3601_/D vssd1 vssd1 vccd1 vccd1 _3601_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1793_ hold71/A _3563_/Q _3575_/Q _3240_/Q _2289_/B _2289_/C vssd1 vssd1 vccd1 vccd1
+ _1793_/X sky130_fd_sc_hd__mux4_1
X_3532_ _3732_/CLK _3532_/D vssd1 vssd1 vccd1 vccd1 _3532_/Q sky130_fd_sc_hd__dfxtp_1
Xhold805 _3670_/Q vssd1 vssd1 vccd1 vccd1 hold805/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold816 _2958_/X vssd1 vssd1 vccd1 vccd1 _3635_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold827 _3636_/Q vssd1 vssd1 vccd1 vccd1 hold827/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1725__S _1988_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold849 _2901_/X vssd1 vssd1 vccd1 vccd1 _3616_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold838 _3713_/Q vssd1 vssd1 vccd1 vccd1 hold838/X sky130_fd_sc_hd__clkbuf_2
X_3463_ _3735_/CLK _3463_/D vssd1 vssd1 vccd1 vccd1 _3463_/Q sky130_fd_sc_hd__dfxtp_1
X_2414_ _3192_/A _2612_/B vssd1 vssd1 vccd1 vccd1 _2420_/S sky130_fd_sc_hd__nor2_2
XFILLER_0_58_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3394_ _3728_/CLK _3394_/D vssd1 vssd1 vccd1 vccd1 _3394_/Q sky130_fd_sc_hd__dfxtp_1
X_2345_ _2651_/A0 hold883/X _2349_/S vssd1 vssd1 vccd1 vccd1 _2345_/X sky130_fd_sc_hd__mux2_1
X_2276_ _2276_/A _2278_/B vssd1 vssd1 vccd1 vccd1 _2276_/X sky130_fd_sc_hd__or2_1
XANTENNA__2492__A0 _2651_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2320__A _3055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2180__C1 _3055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2235__A0 _3197_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2868__C _2868_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3045__B _3045_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2171__C1 _3055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2130_ _3713_/Q _2126_/Y _2128_/Y _2129_/X _2132_/C vssd1 vssd1 vccd1 vccd1 _2130_/X
+ sky130_fd_sc_hd__o221a_1
X_2061_ _2046_/A _2955_/A _2076_/C hold983/X _1979_/A vssd1 vssd1 vccd1 vccd1 _2061_/X
+ sky130_fd_sc_hd__o311a_1
XANTENNA__2226__A0 _2653_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2963_ hold39/X _2963_/A1 _2999_/S vssd1 vssd1 vccd1 vccd1 hold40/A sky130_fd_sc_hd__mux2_1
XFILLER_0_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1914_ _2479_/A _1899_/X _2228_/B vssd1 vssd1 vccd1 vccd1 _1914_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_71_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2894_ _2892_/A _2944_/B hold989/X _2859_/A vssd1 vssd1 vccd1 vccd1 _3615_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_44_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2529__A1 _2353_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1845_ _3540_/Q _3250_/Q _3516_/Q _3504_/Q _2000_/S0 _2219_/C vssd1 vssd1 vccd1 vccd1
+ _1845_/X sky130_fd_sc_hd__mux4_1
Xhold602 _2197_/X vssd1 vssd1 vccd1 vccd1 _3235_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1776_ _3435_/Q _3423_/Q _3411_/Q _3267_/Q _1981_/S0 _1981_/S1 vssd1 vssd1 vccd1
+ vccd1 _1776_/X sky130_fd_sc_hd__mux4_1
Xhold635 _3355_/Q vssd1 vssd1 vccd1 vccd1 hold635/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold613 _3539_/Q vssd1 vssd1 vccd1 vccd1 hold613/X sky130_fd_sc_hd__dlygate4sd3_1
X_3515_ _3539_/CLK _3515_/D vssd1 vssd1 vccd1 vccd1 _3515_/Q sky130_fd_sc_hd__dfxtp_1
Xhold624 _2332_/X vssd1 vssd1 vccd1 vccd1 _3316_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold657 _3253_/Q vssd1 vssd1 vccd1 vccd1 hold657/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold668 _2259_/X vssd1 vssd1 vccd1 vccd1 _3285_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold646 _2264_/X vssd1 vssd1 vccd1 vccd1 _3289_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold679 _3287_/Q vssd1 vssd1 vccd1 vccd1 hold679/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3446_ _3447_/CLK _3446_/D vssd1 vssd1 vccd1 vccd1 _3446_/Q sky130_fd_sc_hd__dfxtp_1
X_3377_ _3583_/CLK _3377_/D vssd1 vssd1 vccd1 vccd1 _3377_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2328_ _2326_/X _2327_/X _3096_/A vssd1 vssd1 vccd1 vccd1 _2328_/X sky130_fd_sc_hd__o21a_1
X_2259_ hold667/X _2660_/A0 _2259_/S vssd1 vssd1 vccd1 vccd1 _2259_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_34_wb_clk_i clkbuf_3_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3344_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_67_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2217__A0 _2659_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2940__A1 _1712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2050__A _2050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2940__B2 _2940_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2208__A0 _2652_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1630_ _3035_/A _3027_/A _3677_/Q _3026_/B vssd1 vssd1 vccd1 vccd1 _1630_/X sky130_fd_sc_hd__or4_1
X_3300_ _3344_/CLK _3300_/D vssd1 vssd1 vccd1 vccd1 _3300_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3231_ _3322_/CLK _3231_/D vssd1 vssd1 vccd1 vccd1 _3231_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3162_ hold936/X _3158_/Y _3161_/X _3166_/C1 vssd1 vssd1 vccd1 vccd1 _3162_/X sky130_fd_sc_hd__o211a_1
X_2113_ _2237_/A _2619_/A vssd1 vssd1 vccd1 vccd1 _2119_/S sky130_fd_sc_hd__nand2_4
XFILLER_0_55_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3093_ wire109/X _2311_/B _3091_/X _3092_/Y vssd1 vssd1 vccd1 vccd1 _3093_/X sky130_fd_sc_hd__a31o_1
X_2044_ hold589/X _2731_/A2 _2867_/B _2034_/X vssd1 vssd1 vccd1 vccd1 _2044_/X sky130_fd_sc_hd__o22a_1
XANTENNA__2447__A0 _2475_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2946_ _3103_/A _2946_/B vssd1 vssd1 vccd1 vccd1 _3624_/D sky130_fd_sc_hd__and2_1
X_2877_ _2876_/A _2876_/B _2159_/B _2876_/X _2960_/A vssd1 vssd1 vccd1 vccd1 _2877_/X
+ sky130_fd_sc_hd__o311a_2
XFILLER_0_44_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1828_ _3430_/Q _3418_/Q _3406_/Q _3262_/Q _1760_/A _1760_/B vssd1 vssd1 vccd1 vccd1
+ _1828_/X sky130_fd_sc_hd__mux4_1
Xhold410 _2971_/X vssd1 vssd1 vccd1 vccd1 _3646_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold421 _3743_/Q vssd1 vssd1 vccd1 vccd1 hold421/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold454 _2568_/X vssd1 vssd1 vccd1 vccd1 _3508_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold432 _2611_/X vssd1 vssd1 vccd1 vccd1 _3545_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold443 _3521_/Q vssd1 vssd1 vccd1 vccd1 hold443/X sky130_fd_sc_hd__dlygate4sd3_1
X_1759_ _1755_/Y _1756_/X _1758_/X _2022_/A vssd1 vssd1 vccd1 vccd1 _1759_/Y sky130_fd_sc_hd__o211ai_1
Xhold465 _3541_/Q vssd1 vssd1 vccd1 vccd1 hold465/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold476 _2396_/X vssd1 vssd1 vccd1 vccd1 _3366_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold487 _3454_/Q vssd1 vssd1 vccd1 vccd1 hold487/X sky130_fd_sc_hd__dlygate4sd3_1
X_3429_ _3733_/CLK _3429_/D vssd1 vssd1 vccd1 vccd1 _3429_/Q sky130_fd_sc_hd__dfxtp_1
Xhold498 _2967_/X vssd1 vssd1 vccd1 vccd1 _3642_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2989__A1 _1760_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2610__A0 _2659_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2800_ _2803_/B _2803_/C _2789_/S vssd1 vssd1 vccd1 vccd1 _2800_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_81_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2601__A0 _3195_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2731_ _2082_/C _2731_/A2 _2854_/B vssd1 vssd1 vccd1 vccd1 _2731_/X sky130_fd_sc_hd__a21o_2
XFILLER_0_54_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2662_ hold237/X _2353_/A _2667_/S vssd1 vssd1 vccd1 vccd1 _2662_/X sky130_fd_sc_hd__mux2_1
X_2593_ hold111/X _3201_/A1 _2597_/S vssd1 vssd1 vccd1 vccd1 _2593_/X sky130_fd_sc_hd__mux2_1
X_1613_ _3626_/Q vssd1 vssd1 vccd1 vccd1 _2712_/A sky130_fd_sc_hd__inv_2
XANTENNA__1733__S _2244_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3214_ _3739_/CLK _3214_/D vssd1 vssd1 vccd1 vccd1 _3214_/Q sky130_fd_sc_hd__dfxtp_1
X_3145_ _2924_/B _2886_/A _3137_/C vssd1 vssd1 vccd1 vccd1 _3145_/X sky130_fd_sc_hd__a21o_1
X_3076_ _2310_/B _3075_/X _3048_/B vssd1 vssd1 vccd1 vccd1 _3076_/Y sky130_fd_sc_hd__o21ai_1
X_2027_ _2997_/A1 _1769_/Y _2026_/X _2854_/B vssd1 vssd1 vccd1 vccd1 _2027_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_82_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2929_ _2929_/A _2941_/C vssd1 vssd1 vccd1 vccd1 _2935_/B sky130_fd_sc_hd__and2_1
XFILLER_0_17_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold251 _3429_/Q vssd1 vssd1 vccd1 vccd1 hold251/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold262 _2629_/X vssd1 vssd1 vccd1 vccd1 _3560_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2356__C1 _3058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold240 _2994_/X vssd1 vssd1 vccd1 vccd1 _3669_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold273 _3478_/Q vssd1 vssd1 vccd1 vccd1 hold273/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold295 _3472_/Q vssd1 vssd1 vccd1 vccd1 hold295/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold284 _2513_/X vssd1 vssd1 vccd1 vccd1 _3461_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2659__A0 _2659_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout74_A _2099_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput8 io_in[17] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__buf_1
XFILLER_0_78_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1873__B2 _2854_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1720__S1 _1981_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3694_ _3714_/CLK _3694_/D vssd1 vssd1 vccd1 vccd1 _3694_/Q sky130_fd_sc_hd__dfxtp_1
X_2714_ _2803_/A _2714_/B vssd1 vssd1 vccd1 vccd1 _2716_/B sky130_fd_sc_hd__xnor2_1
X_2645_ hold151/X _2659_/A0 _2646_/S vssd1 vssd1 vccd1 vccd1 _2645_/X sky130_fd_sc_hd__mux2_1
X_2576_ _2363_/A hold429/X _2576_/S vssd1 vssd1 vccd1 vccd1 _2576_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_10_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1864__A1 _2479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3128_ hold811/X _3118_/A _3126_/A _3115_/X vssd1 vssd1 vccd1 vccd1 _3128_/X sky130_fd_sc_hd__a211o_1
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3059_ _3059_/A _3059_/B _3226_/Q _2153_/A vssd1 vssd1 vccd1 vccd1 _3096_/C sky130_fd_sc_hd__or4b_2
XANTENNA_clkbuf_leaf_42_wb_clk_i_A clkbuf_3_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_37_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2041__B2 _2854_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2041__A1 _1760_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2042__B _2076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1778__S1 _2245_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1855__A1 _2244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2280__A1 _2480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3048__B _3048_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2430_ _2619_/A _2528_/B vssd1 vssd1 vccd1 vccd1 _2436_/S sky130_fd_sc_hd__and2_2
X_2361_ _2361_/A _2363_/B vssd1 vssd1 vccd1 vccd1 _2361_/X sky130_fd_sc_hd__or2_1
XFILLER_0_47_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2292_ hold55/X _2355_/A _2296_/S vssd1 vssd1 vccd1 vccd1 hold56/A sky130_fd_sc_hd__mux2_1
XFILLER_0_37_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1941__S1 _2185_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2271__A1 _2022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout124_A _3348_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3677_ _3727_/CLK _3677_/D vssd1 vssd1 vccd1 vccd1 _3677_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_30_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2628_ hold579/X _2656_/A0 _2632_/S vssd1 vssd1 vccd1 vccd1 _2628_/X sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_9_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_2559_ hold235/X _2357_/A _2562_/S vssd1 vssd1 vccd1 vccd1 _2559_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1932__S1 _1760_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1831__S _1937_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1930_ _3384_/Q _3372_/Q _3360_/Q _3288_/Q _1981_/S0 _1981_/S1 vssd1 vssd1 vccd1
+ vccd1 _1930_/X sky130_fd_sc_hd__mux4_1
X_1861_ _2085_/C _1861_/B vssd1 vssd1 vccd1 vccd1 _1861_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_56_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput11 io_in[20] vssd1 vssd1 vccd1 vccd1 input11/X sky130_fd_sc_hd__buf_1
X_3600_ _3662_/CLK _3600_/D vssd1 vssd1 vccd1 vccd1 _3600_/Q sky130_fd_sc_hd__dfxtp_1
X_3531_ _3732_/CLK hold44/X vssd1 vssd1 vccd1 vccd1 hold43/A sky130_fd_sc_hd__dfxtp_1
X_1792_ _3285_/Q _3357_/Q _3369_/Q _3381_/Q _2000_/S0 _2219_/C vssd1 vssd1 vccd1 vccd1
+ _1792_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold817 _3698_/Q vssd1 vssd1 vccd1 vccd1 hold817/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold806 _2995_/X vssd1 vssd1 vccd1 vccd1 _3670_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold828 _2959_/X vssd1 vssd1 vccd1 vccd1 _3636_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold839 _3180_/X vssd1 vssd1 vccd1 vccd1 _3725_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3462_ _3496_/CLK _3462_/D vssd1 vssd1 vccd1 vccd1 _3462_/Q sky130_fd_sc_hd__dfxtp_1
X_2413_ _2660_/A0 hold655/X _2413_/S vssd1 vssd1 vccd1 vccd1 _2413_/X sky130_fd_sc_hd__mux2_1
X_3393_ _3587_/CLK _3393_/D vssd1 vssd1 vccd1 vccd1 _3393_/Q sky130_fd_sc_hd__dfxtp_1
X_2344_ _3108_/A _2344_/B vssd1 vssd1 vccd1 vccd1 _3324_/D sky130_fd_sc_hd__or2_1
X_2275_ _1716_/X _2245_/C _2651_/A0 _2274_/X _3058_/A vssd1 vssd1 vccd1 vccd1 _2275_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_90_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3729_ _3733_/CLK _3729_/D vssd1 vssd1 vccd1 vccd1 _3729_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2483__A1 _2355_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1746__B1 _2087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_4_wb_clk_i clkbuf_leaf_5_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3419_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__2868__D _2868_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2230__B _2598_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2060_ _2717_/B _2062_/B vssd1 vssd1 vccd1 vccd1 _2060_/X sky130_fd_sc_hd__or2_1
XFILLER_0_44_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1797__A _2085_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2962_ hold249/X _2962_/A1 _2992_/S vssd1 vssd1 vccd1 vccd1 _2962_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_29_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1913_ _2085_/A _1910_/Y _1912_/Y _2228_/C _1908_/Y vssd1 vssd1 vccd1 vccd1 _1913_/X
+ sky130_fd_sc_hd__a311o_1
X_2893_ _2876_/A _2891_/X _2892_/Y _2948_/B _2944_/B vssd1 vssd1 vccd1 vccd1 _2893_/Y
+ sky130_fd_sc_hd__o221ai_1
X_1844_ _3388_/Q _3582_/Q _3564_/Q _3552_/Q _2000_/S0 _2219_/C vssd1 vssd1 vccd1 vccd1
+ _1844_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_44_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1775_ _3497_/Q hold15/A _3467_/Q _3455_/Q _2000_/S0 _2219_/C vssd1 vssd1 vccd1 vccd1
+ _1775_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_4_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold603 _3451_/Q vssd1 vssd1 vccd1 vccd1 hold603/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold625 _3377_/Q vssd1 vssd1 vccd1 vccd1 hold625/X sky130_fd_sc_hd__dlygate4sd3_1
X_3514_ _3741_/CLK _3514_/D vssd1 vssd1 vccd1 vccd1 _3514_/Q sky130_fd_sc_hd__dfxtp_1
Xhold636 _2383_/X vssd1 vssd1 vccd1 vccd1 _3355_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold614 _2604_/X vssd1 vssd1 vccd1 vccd1 _3539_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold658 _2216_/X vssd1 vssd1 vccd1 vccd1 _3253_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold669 _3491_/Q vssd1 vssd1 vccd1 vccd1 hold669/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold647 _3658_/Q vssd1 vssd1 vccd1 vccd1 hold647/X sky130_fd_sc_hd__dlygate4sd3_1
X_3445_ _3725_/CLK _3445_/D vssd1 vssd1 vccd1 vccd1 _3445_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3376_ _3570_/CLK _3376_/D vssd1 vssd1 vccd1 vccd1 _3376_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2327_ _3706_/Q _3089_/B _2316_/Y _3714_/Q vssd1 vssd1 vccd1 vccd1 _2327_/X sky130_fd_sc_hd__a22o_1
X_2258_ hold147/X _2659_/A0 _2259_/S vssd1 vssd1 vccd1 vccd1 _2258_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3111__C1 _3055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1899__S0 _2289_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2189_ hold175/X _2357_/A _2192_/S vssd1 vssd1 vccd1 vccd1 _2189_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1976__B1 _2867_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3178__C1 _3058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2456__A1 _2361_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2000__S0 _2000_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2392__A0 _3198_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3230_ _3322_/CLK hold24/X vssd1 vssd1 vccd1 vccd1 hold23/A sky130_fd_sc_hd__dfxtp_1
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3161_ _3716_/Q _3181_/B vssd1 vssd1 vccd1 vccd1 _3161_/X sky130_fd_sc_hd__or2_1
X_2112_ _2084_/A _2084_/B _2244_/A _2085_/B _2014_/A vssd1 vssd1 vccd1 vccd1 _2619_/A
+ sky130_fd_sc_hd__o2111a_4
X_3092_ _3092_/A _3183_/B vssd1 vssd1 vccd1 vccd1 _3092_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_55_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2043_ _2031_/Y _2041_/X _2042_/X _1979_/A vssd1 vssd1 vccd1 vccd1 _2043_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_49_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2945_ _2944_/B _2943_/X _2944_/Y hold888/X vssd1 vssd1 vccd1 vccd1 _2946_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1958__B1 _2087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2876_ _2876_/A _2876_/B _2876_/C vssd1 vssd1 vccd1 vccd1 _2876_/X sky130_fd_sc_hd__or3_1
X_1827_ hold19/A _3480_/Q _3462_/Q _3450_/Q _1760_/A _1760_/B vssd1 vssd1 vccd1 vccd1
+ _1827_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold400 _2402_/X vssd1 vssd1 vccd1 vccd1 _3371_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold411 _3320_/Q vssd1 vssd1 vccd1 vccd1 hold411/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2383__A0 _2658_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold422 _3203_/X vssd1 vssd1 vccd1 vccd1 _3743_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold444 _2583_/X vssd1 vssd1 vccd1 vccd1 _3521_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold433 _3582_/Q vssd1 vssd1 vccd1 vccd1 hold433/X sky130_fd_sc_hd__dlygate4sd3_1
X_1758_ _2228_/A _1747_/X _1754_/X _1757_/Y vssd1 vssd1 vccd1 vccd1 _1758_/X sky130_fd_sc_hd__a31o_1
Xhold466 _2607_/X vssd1 vssd1 vccd1 vccd1 _3541_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold477 _3369_/Q vssd1 vssd1 vccd1 vccd1 hold477/X sky130_fd_sc_hd__dlygate4sd3_1
X_1689_ _2669_/A _2868_/B _1654_/B _2159_/D _2819_/A vssd1 vssd1 vccd1 vccd1 _1690_/B
+ sky130_fd_sc_hd__o2111a_1
XFILLER_0_40_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold455 _3579_/Q vssd1 vssd1 vccd1 vccd1 hold455/X sky130_fd_sc_hd__dlygate4sd3_1
X_3428_ _3733_/CLK _3428_/D vssd1 vssd1 vccd1 vccd1 _3428_/Q sky130_fd_sc_hd__dfxtp_1
Xhold499 _3264_/Q vssd1 vssd1 vccd1 vccd1 hold499/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold488 _2505_/X vssd1 vssd1 vccd1 vccd1 _3454_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3359_ _3387_/CLK _3359_/D vssd1 vssd1 vccd1 vccd1 _3359_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2438__A1 _2648_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2730_ _2082_/C _2731_/A2 _2854_/B vssd1 vssd1 vccd1 vccd1 _2730_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_0_26_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2661_ _3199_/A _3185_/B vssd1 vssd1 vccd1 vccd1 _2667_/S sky130_fd_sc_hd__nor2_2
X_1612_ _3322_/Q vssd1 vssd1 vccd1 vccd1 _3769_/A sky130_fd_sc_hd__inv_2
X_2592_ hold93/X _2353_/A _2597_/S vssd1 vssd1 vccd1 vccd1 hold94/A sky130_fd_sc_hd__mux2_1
XFILLER_0_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2117__A0 _2651_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3213_ _3737_/CLK _3213_/D vssd1 vssd1 vccd1 vccd1 _3213_/Q sky130_fd_sc_hd__dfxtp_1
X_3144_ hold858/X _3131_/X _3143_/X _3166_/C1 vssd1 vssd1 vccd1 vccd1 _3144_/X sky130_fd_sc_hd__o211a_1
X_3075_ _3097_/C _3075_/B _3075_/C vssd1 vssd1 vccd1 vccd1 _3075_/X sky130_fd_sc_hd__and3_1
XFILLER_0_77_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_32_wb_clk_i_A clkbuf_3_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_2026_ hold285/X _2731_/A2 _2867_/C _1713_/X vssd1 vssd1 vccd1 vccd1 _2026_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_92_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout154_A _3172_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2928_ _1712_/A _3608_/Q hold313/X _2940_/B2 vssd1 vssd1 vccd1 vccd1 _2928_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_72_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2859_ _2859_/A _2859_/B _2859_/C vssd1 vssd1 vccd1 vccd1 _3612_/D sky130_fd_sc_hd__and3_1
XFILLER_0_31_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold252 _2471_/X vssd1 vssd1 vccd1 vccd1 _3429_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold241 _3232_/Q vssd1 vssd1 vccd1 vccd1 hold241/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold230 _3194_/X vssd1 vssd1 vccd1 vccd1 _3735_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold274 _2533_/X vssd1 vssd1 vccd1 vccd1 _3478_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold296 _2526_/X vssd1 vssd1 vccd1 vccd1 _3472_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold285 _3672_/Q vssd1 vssd1 vccd1 vccd1 hold285/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold263 _3274_/Q vssd1 vssd1 vccd1 vccd1 hold263/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2108__A0 _3195_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2347__A0 _2652_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput9 io_in[18] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__buf_1
XFILLER_0_86_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2586__A0 _2656_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3693_ _3714_/CLK _3693_/D vssd1 vssd1 vccd1 vccd1 _3693_/Q sky130_fd_sc_hd__dfxtp_1
X_2713_ _2809_/A _2713_/B _2711_/Y vssd1 vssd1 vccd1 vccd1 _2713_/X sky130_fd_sc_hd__or3b_1
X_2644_ hold605/X _2658_/A0 _2646_/S vssd1 vssd1 vccd1 vccd1 _2644_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_72_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2575_ _2361_/A hold221/X _2576_/S vssd1 vssd1 vccd1 vccd1 _2575_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2889__A1 _2876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3127_ hold811/X _3120_/A _3126_/X _3055_/A vssd1 vssd1 vccd1 vccd1 _3127_/X sky130_fd_sc_hd__o211a_1
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3058_ _3058_/A _3058_/B vssd1 vssd1 vccd1 vccd1 _3689_/D sky130_fd_sc_hd__and2_1
X_2009_ _2244_/A _2004_/X _2087_/A vssd1 vssd1 vccd1 vccd1 _2009_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_92_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2042__C _3045_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2501__A0 _2655_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2280__A2 _2195_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2568__A0 _2659_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2514__A _2640_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2360_ hold956/X _2351_/Y _2359_/X _3172_/C1 vssd1 vssd1 vccd1 vccd1 _3331_/D sky130_fd_sc_hd__o211a_1
X_2291_ hold131/X _2648_/A0 _2296_/S vssd1 vssd1 vccd1 vccd1 _2291_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_47_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2099__A2 _2084_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_22 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2271__A2 _2245_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3745_ _3745_/CLK _3745_/D vssd1 vssd1 vccd1 vccd1 _3745_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2023__A2 _2022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1782__A1 _2006_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3676_ _3676_/CLK _3676_/D vssd1 vssd1 vccd1 vccd1 _3676_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA_fanout117_A _2480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_28_wb_clk_i clkbuf_3_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3733_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_2627_ hold63/X _2089_/X _2632_/S vssd1 vssd1 vccd1 vccd1 hold64/A sky130_fd_sc_hd__mux2_1
XFILLER_0_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2558_ hold141/X _3201_/A1 _2562_/S vssd1 vssd1 vccd1 vccd1 _2558_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_10_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2731__B1 _2854_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2489_ _2648_/A0 hold225/X _2494_/S vssd1 vssd1 vccd1 vccd1 _2489_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_77_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2798__B1 _2731_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2244__A _2244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1860_ _3229_/Q _3244_/Q _2085_/B vssd1 vssd1 vccd1 vccd1 _1861_/B sky130_fd_sc_hd__mux2_1
Xinput12 io_in[29] vssd1 vssd1 vccd1 vccd1 _3058_/B sky130_fd_sc_hd__buf_1
XFILLER_0_83_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3202__A1 _2357_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1791_ _3545_/Q _3255_/Q _3521_/Q _3509_/Q _2000_/S0 _2219_/C vssd1 vssd1 vccd1 vccd1
+ _1791_/X sky130_fd_sc_hd__mux4_1
X_3530_ _3592_/CLK _3530_/D vssd1 vssd1 vccd1 vccd1 _3530_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold818 _3117_/X vssd1 vssd1 vccd1 vccd1 _3698_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold807 _3694_/Q vssd1 vssd1 vccd1 vccd1 hold807/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1764__A1 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3461_ _3745_/CLK _3461_/D vssd1 vssd1 vccd1 vccd1 _3461_/Q sky130_fd_sc_hd__dfxtp_1
Xhold829 _3683_/Q vssd1 vssd1 vccd1 vccd1 _3063_/B sky130_fd_sc_hd__buf_2
X_2412_ _2659_/A0 hold355/X _2413_/S vssd1 vssd1 vccd1 vccd1 _2412_/X sky130_fd_sc_hd__mux2_1
X_3392_ _3586_/CLK _3392_/D vssd1 vssd1 vccd1 vccd1 _3392_/Q sky130_fd_sc_hd__dfxtp_1
X_2343_ _2650_/A0 hold880/X _2349_/S vssd1 vssd1 vccd1 vccd1 _2344_/B sky130_fd_sc_hd__mux2_1
X_2274_ _2274_/A _2278_/B vssd1 vssd1 vccd1 vccd1 _2274_/X sky130_fd_sc_hd__or2_1
XFILLER_0_90_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1989_ _2245_/B _1989_/B vssd1 vssd1 vccd1 vccd1 _1989_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_70_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3728_ _3728_/CLK hold32/X vssd1 vssd1 vccd1 vccd1 hold31/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3659_ _3661_/CLK _3659_/D vssd1 vssd1 vccd1 vccd1 _3659_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3196__A0 _3196_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1746__A1 _2244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2961_ _2961_/A _2961_/B vssd1 vssd1 vccd1 vccd1 _2961_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_8_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1912_ _2085_/C _1912_/B vssd1 vssd1 vccd1 vccd1 _1912_/Y sky130_fd_sc_hd__nand2_1
X_2892_ _2892_/A _2892_/B vssd1 vssd1 vccd1 vccd1 _2892_/Y sky130_fd_sc_hd__xnor2_1
X_1843_ _2185_/A _1840_/Y _1842_/Y _2428_/C _1838_/Y vssd1 vssd1 vccd1 vccd1 _1843_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_0_8_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1774_ _3387_/Q _3375_/Q _3363_/Q _3291_/Q _1981_/S0 _1981_/S1 vssd1 vssd1 vccd1
+ vccd1 _1774_/X sky130_fd_sc_hd__mux4_1
Xhold626 _2409_/X vssd1 vssd1 vccd1 vccd1 _3377_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3513_ _3741_/CLK _3513_/D vssd1 vssd1 vccd1 vccd1 _3513_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2421__B _2612_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold604 _2502_/X vssd1 vssd1 vccd1 vccd1 _3451_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold615 _3423_/Q vssd1 vssd1 vccd1 vccd1 hold615/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold648 _2983_/X vssd1 vssd1 vccd1 vccd1 _3658_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold637 _3409_/Q vssd1 vssd1 vccd1 vccd1 hold637/X sky130_fd_sc_hd__dlygate4sd3_1
X_3444_ _3581_/CLK _3444_/D vssd1 vssd1 vccd1 vccd1 _3444_/Q sky130_fd_sc_hd__dfxtp_1
Xhold659 _3301_/Q vssd1 vssd1 vccd1 vccd1 hold659/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1752__S _1937_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3375_ _3387_/CLK _3375_/D vssd1 vssd1 vccd1 vccd1 _3375_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2326_ _3710_/Q _3226_/Q _3089_/A _3227_/Q vssd1 vssd1 vccd1 vccd1 _2326_/X sky130_fd_sc_hd__o211a_1
X_2257_ hold135/X _2658_/A0 _2259_/S vssd1 vssd1 vccd1 vccd1 _2257_/X sky130_fd_sc_hd__mux2_1
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1899__S1 _2479_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2188_ hold23/X _2355_/A _2192_/S vssd1 vssd1 vccd1 vccd1 hold24/A sky130_fd_sc_hd__mux2_1
XFILLER_0_79_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_43_wb_clk_i clkbuf_3_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3692_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__1728__A1 _1889_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2331__B _2647_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout97_A _2987_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2000__S1 _2219_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1967__A1 _2479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3160_ hold898/X _3158_/Y hold964/X _3086_/A vssd1 vssd1 vccd1 vccd1 _3160_/X sky130_fd_sc_hd__o211a_1
X_2111_ _2660_/A0 hold609/X _2111_/S vssd1 vssd1 vccd1 vccd1 _2111_/X sky130_fd_sc_hd__mux2_1
X_3091_ _2300_/A _3089_/X _3090_/Y _3048_/B vssd1 vssd1 vccd1 vccd1 _3091_/X sky130_fd_sc_hd__a31o_1
Xhold1 hold1/A vssd1 vssd1 vccd1 vccd1 hold1/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2042_ _2071_/A _2076_/A _3045_/B _2042_/D vssd1 vssd1 vccd1 vccd1 _2042_/X sky130_fd_sc_hd__or4_1
XANTENNA_clkbuf_leaf_22_wb_clk_i_A clkbuf_3_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_49_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2944_ _2942_/Y _2944_/B vssd1 vssd1 vccd1 vccd1 _2944_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__1958__A1 _2244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2875_ _2823_/Y _2873_/X _2875_/B1 _2859_/A vssd1 vssd1 vccd1 vccd1 _2875_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_29_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1826_ _3382_/Q _3370_/Q _3358_/Q _3286_/Q _1981_/S0 _1981_/S1 vssd1 vssd1 vccd1
+ vccd1 _1826_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_40_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold401 _3212_/Q vssd1 vssd1 vccd1 vccd1 hold401/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold445 _3510_/Q vssd1 vssd1 vccd1 vccd1 hold445/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold434 _2655_/X vssd1 vssd1 vccd1 vccd1 _3582_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1757_ _2480_/A _1721_/X _2195_/B vssd1 vssd1 vccd1 vccd1 _1757_/Y sky130_fd_sc_hd__o21ai_1
Xhold423 _3633_/Q vssd1 vssd1 vccd1 vccd1 _1870_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold412 _2336_/X vssd1 vssd1 vccd1 vccd1 _3320_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold478 _2399_/X vssd1 vssd1 vccd1 vccd1 _3369_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1688_ _2819_/A _2159_/D vssd1 vssd1 vccd1 vccd1 _2878_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_40_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold456 _2651_/X vssd1 vssd1 vccd1 vccd1 _3579_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold467 _3223_/Q vssd1 vssd1 vccd1 vccd1 hold467/X sky130_fd_sc_hd__dlygate4sd3_1
X_3427_ _3732_/CLK _3427_/D vssd1 vssd1 vccd1 vccd1 _3427_/Q sky130_fd_sc_hd__dfxtp_1
Xhold489 _3664_/Q vssd1 vssd1 vccd1 vccd1 hold489/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3358_ _3654_/CLK _3358_/D vssd1 vssd1 vccd1 vccd1 _3358_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2309_ _2309_/A _3045_/A vssd1 vssd1 vccd1 vccd1 _3007_/A sky130_fd_sc_hd__nand2_2
XANTENNA__1894__B1 _2428_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3289_ _3654_/CLK _3289_/D vssd1 vssd1 vccd1 vccd1 _3289_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2342__A _3108_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3157__B _3157_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2374__A1 _2355_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold990 _3228_/Q vssd1 vssd1 vccd1 vccd1 _2182_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_25_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1980__S0 _1981_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2834__C1 _2859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2660_ _2660_/A0 hold301/X _2660_/S vssd1 vssd1 vccd1 vccd1 _2660_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1611_ _3323_/Q vssd1 vssd1 vccd1 vccd1 _3770_/A sky130_fd_sc_hd__inv_2
X_2591_ _2640_/A _3185_/B vssd1 vssd1 vccd1 vccd1 _2597_/S sky130_fd_sc_hd__nor2_4
XFILLER_0_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3212_ _3737_/CLK _3212_/D vssd1 vssd1 vccd1 vccd1 _3212_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3143_ _2914_/A _2886_/A _3137_/C vssd1 vssd1 vccd1 vccd1 _3143_/X sky130_fd_sc_hd__a21o_1
X_3074_ _3688_/Q _3687_/Q _3097_/A _3037_/C vssd1 vssd1 vccd1 vccd1 _3075_/C sky130_fd_sc_hd__or4b_1
XFILLER_0_77_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2025_ hold827/X _1922_/B _2023_/X _2024_/X vssd1 vssd1 vccd1 vccd1 _2867_/C sky130_fd_sc_hd__o22a_4
XFILLER_0_49_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout147_A _2961_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2927_ _2924_/A _2944_/B hold993/X _3103_/A vssd1 vssd1 vccd1 vccd1 _3621_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_45_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1800__B1 _2087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2858_ hold996/X _2858_/B vssd1 vssd1 vccd1 vccd1 _2859_/C sky130_fd_sc_hd__nand2b_1
X_1809_ _2087_/A _1785_/Y _1789_/Y _1783_/Y _2479_/A vssd1 vssd1 vccd1 vccd1 _1809_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_60_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2789_ _2709_/C _2788_/Y _2789_/S vssd1 vssd1 vccd1 vccd1 _2790_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_32_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold220 _2554_/X vssd1 vssd1 vccd1 vccd1 _3496_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold231 _3426_/Q vssd1 vssd1 vccd1 vccd1 hold231/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold253 _3439_/Q vssd1 vssd1 vccd1 vccd1 hold253/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold242 _2190_/X vssd1 vssd1 vccd1 vccd1 _3232_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold286 _2997_/X vssd1 vssd1 vccd1 vccd1 _3672_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold264 _2247_/X vssd1 vssd1 vccd1 vccd1 _3274_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold275 _3453_/Q vssd1 vssd1 vccd1 vccd1 hold275/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold297 _3644_/Q vssd1 vssd1 vccd1 vccd1 hold297/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2044__B1 _2867_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2595__A1 _3203_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1850__S _1954_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2283__A0 _2648_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2035__B1 _2701_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2712_ _2712_/A _3627_/Q _3628_/Q vssd1 vssd1 vccd1 vccd1 _2713_/B sky130_fd_sc_hd__or3_1
X_3692_ _3692_/CLK _3692_/D vssd1 vssd1 vccd1 vccd1 _3692_/Q sky130_fd_sc_hd__dfxtp_1
X_2643_ hold419/X _2643_/A1 _2646_/S vssd1 vssd1 vccd1 vccd1 _2643_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_14_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2574_ _3203_/A1 hold223/X _2576_/S vssd1 vssd1 vccd1 vccd1 _2574_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_77_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2510__A1 _2357_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3126_ _3126_/A _3126_/B vssd1 vssd1 vccd1 vccd1 _3126_/X sky130_fd_sc_hd__or2_1
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3057_ _3065_/A _3055_/C _3056_/X _3108_/A vssd1 vssd1 vccd1 vccd1 _3057_/Y sky130_fd_sc_hd__a211oi_1
X_2008_ _3772_/A _2005_/S _2006_/A _2007_/Y vssd1 vssd1 vccd1 vccd1 _2008_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_77_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2026__B1 _2867_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1935__S _1937_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold908_A _3594_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2265__A0 _3197_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2017__B1 _2087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2280__A3 _2087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2290_ _2290_/A _2612_/B vssd1 vssd1 vccd1 vccd1 _2296_/S sky130_fd_sc_hd__nor2_2
XFILLER_0_2_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2271__A3 _2355_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2008__B1 _2006_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2559__A1 _2357_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3744_ _3744_/CLK _3744_/D vssd1 vssd1 vccd1 vccd1 _3744_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3675_ _3676_/CLK _3675_/D vssd1 vssd1 vccd1 vccd1 _3675_/Q sky130_fd_sc_hd__dfxtp_1
X_2626_ _2640_/B _3199_/A vssd1 vssd1 vccd1 vccd1 _2632_/S sky130_fd_sc_hd__nor2_2
XFILLER_0_2_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2557_ hold183/X _2353_/A _2562_/S vssd1 vssd1 vccd1 vccd1 _2557_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2488_ _2570_/A _2647_/B vssd1 vssd1 vccd1 vccd1 _2494_/S sky130_fd_sc_hd__nand2_4
X_3109_ hold785/X _3037_/D _3183_/B vssd1 vssd1 vccd1 vccd1 _3110_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_65_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2798__A1 _2797_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2350__A _3108_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2228__C _2228_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2238__A0 _2648_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2244__B _2244_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput13 io_in[3] vssd1 vssd1 vccd1 vccd1 _2074_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_83_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1790_ _3393_/Q _3587_/Q _3569_/Q _3557_/Q _2000_/S0 _2219_/C vssd1 vssd1 vccd1 vccd1
+ _1790_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_12_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold808 _3102_/Y vssd1 vssd1 vccd1 vccd1 _3103_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold819 _3650_/Q vssd1 vssd1 vccd1 vccd1 _1627_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3460_ _3745_/CLK hold12/X vssd1 vssd1 vccd1 vccd1 hold11/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2411_ _2658_/A0 hold709/X _2413_/S vssd1 vssd1 vccd1 vccd1 _2411_/X sky130_fd_sc_hd__mux2_1
X_3391_ _3585_/CLK _3391_/D vssd1 vssd1 vccd1 vccd1 _3391_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2342_ _3108_/A _2342_/B vssd1 vssd1 vccd1 vccd1 _3323_/D sky130_fd_sc_hd__or2_1
XANTENNA__1921__C1 _1922_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1604__A _2876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2273_ _2022_/A _2245_/C _2650_/A0 _2272_/X _3058_/A vssd1 vssd1 vccd1 vccd1 _3294_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_74_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2229__B1 _2480_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1988_ hold77/A _3489_/Q _1988_/S vssd1 vssd1 vccd1 vccd1 _1989_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_7_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3727_ _3727_/CLK _3727_/D vssd1 vssd1 vccd1 vccd1 _3727_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2401__A0 _3193_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3658_ _3661_/CLK _3658_/D vssd1 vssd1 vccd1 vccd1 _3658_/Q sky130_fd_sc_hd__dfxtp_1
X_2609_ _2658_/A0 hold483/X _2611_/S vssd1 vssd1 vccd1 vccd1 _2609_/X sky130_fd_sc_hd__mux2_1
X_3589_ _3745_/CLK _3589_/D vssd1 vssd1 vccd1 vccd1 _3589_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2180__A2 _3157_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2468__A0 _2650_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2064__B _3045_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2943__A1 _2885_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_12_wb_clk_i_A clkbuf_3_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__2459__A0 _3193_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1682__A1 _2960_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output23_A _3771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2960_ _2960_/A _3137_/B vssd1 vssd1 vccd1 vccd1 _2961_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_84_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2891_ hold39/X _2940_/B2 _2687_/B _2819_/A vssd1 vssd1 vccd1 vccd1 _2891_/X sky130_fd_sc_hd__o2bb2a_1
X_1911_ hold23/A _3245_/Q _2085_/B vssd1 vssd1 vccd1 vccd1 _1912_/B sky130_fd_sc_hd__mux2_1
X_1842_ _2006_/A _1842_/B vssd1 vssd1 vccd1 vccd1 _1842_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_44_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3187__A1 _3201_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1773_ _3739_/Q _3217_/Q _3321_/Q _3339_/Q _1981_/S0 _2219_/C vssd1 vssd1 vccd1 vccd1
+ _1773_/X sky130_fd_sc_hd__mux4_1
XANTENNA__2934__A1 _1712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold605 _3573_/Q vssd1 vssd1 vccd1 vccd1 hold605/X sky130_fd_sc_hd__dlygate4sd3_1
X_3512_ _3539_/CLK _3512_/D vssd1 vssd1 vccd1 vccd1 _3512_/Q sky130_fd_sc_hd__dfxtp_1
Xhold627 _3506_/Q vssd1 vssd1 vccd1 vccd1 hold627/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2934__B2 _2940_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold616 _2464_/X vssd1 vssd1 vccd1 vccd1 _3423_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold649 _3384_/Q vssd1 vssd1 vccd1 vccd1 hold649/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold638 _2448_/X vssd1 vssd1 vccd1 vccd1 _3409_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3443_ _3724_/CLK _3443_/D vssd1 vssd1 vccd1 vccd1 _3443_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_51_wb_clk_i_A clkbuf_3_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3374_ _3654_/CLK _3374_/D vssd1 vssd1 vccd1 vccd1 _3374_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2325_ hold840/X _2318_/B _2324_/Y _3108_/A vssd1 vssd1 vccd1 vccd1 _2325_/X sky130_fd_sc_hd__a211o_1
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2256_ hold413/X _3195_/A0 _2259_/S vssd1 vssd1 vccd1 vccd1 _2256_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_79_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2187_ hold145/X _2648_/A0 _2192_/S vssd1 vssd1 vccd1 vccd1 _2187_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2622__A0 _3195_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1976__A2 _2731_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2612__B _2612_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1943__S _2244_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_12_wb_clk_i clkbuf_3_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3587_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__3102__A1 _3045_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2916__A1 _2885_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3090_ hold927/X _2313_/X _3089_/B hold898/X vssd1 vssd1 vccd1 vccd1 _3090_/Y sky130_fd_sc_hd__a22oi_1
Xhold2 hold2/A vssd1 vssd1 vccd1 vccd1 hold2/X sky130_fd_sc_hd__dlygate4sd3_1
X_2110_ _3197_/A0 hold763/X _2111_/S vssd1 vssd1 vccd1 vccd1 _2110_/X sky130_fd_sc_hd__mux2_1
X_2041_ _1760_/B _2036_/Y _2040_/X _2854_/B vssd1 vssd1 vccd1 vccd1 _2041_/X sky130_fd_sc_hd__o22a_1
XANTENNA__2604__A0 _2363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2943_ _2885_/B _2940_/X _2949_/A2 _2942_/Y vssd1 vssd1 vccd1 vccd1 _2943_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_29_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2874_ _2874_/A _2874_/B vssd1 vssd1 vccd1 vccd1 _2874_/X sky130_fd_sc_hd__or2_1
X_1825_ _3734_/Q _3212_/Q _3316_/Q _3334_/Q _1981_/S0 _1981_/S1 vssd1 vssd1 vccd1
+ vccd1 _1825_/X sky130_fd_sc_hd__mux4_1
X_1756_ _2479_/A _1728_/X _1735_/X _2195_/B vssd1 vssd1 vccd1 vccd1 _1756_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_4_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold402 _2106_/X vssd1 vssd1 vccd1 vccd1 _3212_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold413 _3282_/Q vssd1 vssd1 vccd1 vccd1 hold413/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold424 _2956_/X vssd1 vssd1 vccd1 vccd1 _3633_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold435 _3666_/Q vssd1 vssd1 vccd1 vccd1 hold435/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold446 _2571_/X vssd1 vssd1 vccd1 vccd1 _3510_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold457 _3248_/Q vssd1 vssd1 vccd1 vccd1 hold457/X sky130_fd_sc_hd__dlygate4sd3_1
X_1687_ _2797_/A _2960_/A _2854_/B _1979_/A vssd1 vssd1 vccd1 vccd1 _3312_/D sky130_fd_sc_hd__o211a_1
Xhold468 _2119_/X vssd1 vssd1 vccd1 vccd1 _3223_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3426_ _3592_/CLK _3426_/D vssd1 vssd1 vccd1 vccd1 _3426_/Q sky130_fd_sc_hd__dfxtp_1
Xhold479 _3290_/Q vssd1 vssd1 vccd1 vccd1 hold479/X sky130_fd_sc_hd__dlygate4sd3_1
X_3357_ _3583_/CLK _3357_/D vssd1 vssd1 vccd1 vccd1 _3357_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1894__A1 _1889_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2308_ _3053_/B _3097_/C _2308_/C vssd1 vssd1 vccd1 vccd1 _2308_/Y sky130_fd_sc_hd__nor3_1
X_3288_ _3387_/CLK _3288_/D vssd1 vssd1 vccd1 vccd1 _3288_/Q sky130_fd_sc_hd__dfxtp_1
X_2239_ _2355_/A hold551/X _2243_/S vssd1 vssd1 vccd1 vccd1 _2239_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1741__S1 _2014_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold991 _2184_/X vssd1 vssd1 vccd1 vccd1 _3228_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold980 _3402_/Q vssd1 vssd1 vccd1 vccd1 hold980/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_hold938_A _3676_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1980__S1 _1981_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1610_ _3324_/Q vssd1 vssd1 vccd1 vccd1 _3771_/A sky130_fd_sc_hd__inv_2
X_2590_ _2363_/A hold757/X _2590_/S vssd1 vssd1 vccd1 vccd1 _2590_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3211_ _3308_/CLK hold26/X vssd1 vssd1 vccd1 vccd1 hold25/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3142_ hold927/X _3131_/X hold960/X _3166_/C1 vssd1 vssd1 vccd1 vccd1 _3142_/X sky130_fd_sc_hd__o211a_1
X_3073_ _2166_/X _3072_/Y _3157_/B vssd1 vssd1 vccd1 vccd1 _3080_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_49_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2024_ input3/X _1920_/B _1677_/X vssd1 vssd1 vccd1 vccd1 _2024_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_15_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2926_ hold992/X _2923_/Y _2941_/C _2925_/Y _2944_/B vssd1 vssd1 vccd1 vccd1 _2926_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_0_72_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1800__A1 _2244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2857_ _2876_/B _2871_/A _2853_/Y _2856_/X vssd1 vssd1 vccd1 vccd1 _2859_/B sky130_fd_sc_hd__a31o_1
XFILLER_0_17_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1808_ _3348_/Q _1805_/Y _1807_/Y _2428_/C _1803_/Y vssd1 vssd1 vccd1 vccd1 _1808_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_0_60_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold210 _2631_/X vssd1 vssd1 vccd1 vccd1 _3562_/D sky130_fd_sc_hd__dlygate4sd3_1
X_2788_ _2788_/A _2788_/B vssd1 vssd1 vccd1 vccd1 _2788_/Y sky130_fd_sc_hd__xnor2_1
Xhold243 _3502_/Q vssd1 vssd1 vccd1 vccd1 hold243/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold221 _3514_/Q vssd1 vssd1 vccd1 vccd1 hold221/X sky130_fd_sc_hd__dlygate4sd3_1
X_1739_ hold7/A _3562_/Q _3574_/Q _3239_/Q _2289_/B _2289_/C vssd1 vssd1 vccd1 vccd1
+ _1739_/X sky130_fd_sc_hd__mux4_1
Xhold232 _2468_/X vssd1 vssd1 vccd1 vccd1 _3426_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold254 _2485_/X vssd1 vssd1 vccd1 vccd1 _3439_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold287 _3458_/Q vssd1 vssd1 vccd1 vccd1 hold287/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold265 _3483_/Q vssd1 vssd1 vccd1 vccd1 hold265/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold276 _2504_/X vssd1 vssd1 vccd1 vccd1 _3453_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold298 _2969_/X vssd1 vssd1 vccd1 vccd1 _3644_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3409_ _3665_/CLK _3409_/D vssd1 vssd1 vccd1 vccd1 _3409_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2292__A1 _2355_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2353__A _2353_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2528__A _2570_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1953__S1 _2014_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2711_ _1606_/Y _2868_/D _2803_/C vssd1 vssd1 vccd1 vccd1 _2711_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_14_106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3691_ _3692_/CLK _3691_/D vssd1 vssd1 vccd1 vccd1 _3691_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2642_ hold619/X _2091_/X _2646_/S vssd1 vssd1 vccd1 vccd1 _2642_/X sky130_fd_sc_hd__mux2_1
X_2573_ _2357_/A hold547/X _2576_/S vssd1 vssd1 vccd1 vccd1 _2573_/X sky130_fd_sc_hd__mux2_1
X_3125_ hold809/X _3183_/B _3118_/X _3124_/Y vssd1 vssd1 vccd1 vccd1 _3126_/B sky130_fd_sc_hd__o22a_1
X_3056_ _3096_/A _3038_/Y _3054_/B _3183_/B _2305_/A vssd1 vssd1 vccd1 vccd1 _3056_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_89_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2007_ _3331_/Q _2244_/B vssd1 vssd1 vccd1 vccd1 _2007_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_77_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2909_ _2914_/B _2914_/C vssd1 vssd1 vccd1 vccd1 _2909_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1880__S0 _2085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout72_A _2099_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2348__A _3108_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2017__A1 _2289_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3150__C1 _3103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output53_A _3310_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2256__A1 _3195_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2008__A1 _3772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3743_ _3743_/CLK _3743_/D vssd1 vssd1 vccd1 vccd1 _3743_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3674_ _3674_/CLK _3674_/D vssd1 vssd1 vccd1 vccd1 _3674_/Q sky130_fd_sc_hd__dfxtp_1
X_2625_ _2660_/A0 hold561/X _2625_/S vssd1 vssd1 vccd1 vccd1 _2625_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_23_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2556_ _3192_/B _3199_/B vssd1 vssd1 vccd1 vccd1 _2562_/S sky130_fd_sc_hd__nor2_2
XFILLER_0_10_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2487_ hold29/X _2363_/A _2487_/S vssd1 vssd1 vccd1 vccd1 hold30/A sky130_fd_sc_hd__mux2_1
XANTENNA__2731__A2 _2731_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3108_ _3108_/A _3108_/B vssd1 vssd1 vccd1 vccd1 _3695_/D sky130_fd_sc_hd__nor2_1
X_3039_ _3040_/A _3038_/Y _3054_/A vssd1 vssd1 vccd1 vccd1 _3039_/X sky130_fd_sc_hd__o21a_1
XANTENNA__2247__A1 _2648_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_37_wb_clk_i clkbuf_3_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3308_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2486__A1 _2361_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2228__D _2480_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput14 io_in[4] vssd1 vssd1 vccd1 vccd1 _2076_/A sky130_fd_sc_hd__buf_4
XANTENNA__1844__S0 _2000_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold809 _3700_/Q vssd1 vssd1 vccd1 vccd1 hold809/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2410_ _2643_/A1 hold585/X _2413_/S vssd1 vssd1 vccd1 vccd1 _2410_/X sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_41_wb_clk_i_A clkbuf_3_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__2260__B _2619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3390_ _3586_/CLK hold84/X vssd1 vssd1 vccd1 vccd1 hold83/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2341_ _2355_/A hold891/X _2349_/S vssd1 vssd1 vccd1 vccd1 _2341_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_58_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2272_ _2272_/A _2278_/B vssd1 vssd1 vccd1 vccd1 _2272_/X sky130_fd_sc_hd__or2_1
XANTENNA__3123__C1 _3055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2477__A1 _3197_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2716__A _3612_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2229__A1 _2289_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1620__A _3058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_423 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1987_ _2006_/A _1987_/B vssd1 vssd1 vccd1 vccd1 _1987_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_74_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2451__A _2647_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout122_A _3349_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3726_ _3727_/CLK _3726_/D vssd1 vssd1 vccd1 vccd1 _3726_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3657_ _3662_/CLK _3657_/D vssd1 vssd1 vccd1 vccd1 _3657_/Q sky130_fd_sc_hd__dfxtp_1
X_2608_ _3195_/A0 hold505/X _2611_/S vssd1 vssd1 vccd1 vccd1 _2608_/X sky130_fd_sc_hd__mux2_1
X_3588_ _3728_/CLK _3588_/D vssd1 vssd1 vccd1 vccd1 _3588_/Q sky130_fd_sc_hd__dfxtp_1
X_2539_ hold265/X _2658_/A0 _2541_/S vssd1 vssd1 vccd1 vccd1 _2539_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3114__C1 _3055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2361__A _2361_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1826__S0 _1981_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2003__S0 _2289_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_8_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_84_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2631__A1 _2659_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2890_ _2892_/B _2883_/Y _2889_/Y _3103_/A vssd1 vssd1 vccd1 vccd1 _2890_/X sky130_fd_sc_hd__o211a_1
X_1910_ _2014_/A _1910_/B vssd1 vssd1 vccd1 vccd1 _1910_/Y sky130_fd_sc_hd__nand2_1
X_1841_ _3456_/Q _3588_/Q _2244_/B vssd1 vssd1 vccd1 vccd1 _1842_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_44_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2395__A0 _2656_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1772_ _1979_/A _1772_/B vssd1 vssd1 vccd1 vccd1 _3610_/D sky130_fd_sc_hd__and2_1
XFILLER_0_52_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold606 _2644_/X vssd1 vssd1 vccd1 vccd1 _3573_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3511_ _3741_/CLK _3511_/D vssd1 vssd1 vccd1 vccd1 _3511_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold617 _3634_/Q vssd1 vssd1 vccd1 vccd1 _1922_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold639 _3365_/Q vssd1 vssd1 vccd1 vccd1 hold639/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold628 _2566_/X vssd1 vssd1 vccd1 vccd1 _3506_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3442_ _3724_/CLK _3442_/D vssd1 vssd1 vccd1 vccd1 _3442_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3373_ _3654_/CLK _3373_/D vssd1 vssd1 vccd1 vccd1 _3373_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2324_ _2311_/B _2323_/Y _2318_/B vssd1 vssd1 vccd1 vccd1 _2324_/Y sky130_fd_sc_hd__a21oi_1
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2255_ hold129/X _2656_/A0 _2259_/S vssd1 vssd1 vccd1 vccd1 _2255_/X sky130_fd_sc_hd__mux2_1
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2186_ _2290_/A _3192_/B vssd1 vssd1 vccd1 vccd1 _2192_/S sky130_fd_sc_hd__nor2_2
XFILLER_0_79_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3709_ _3718_/CLK _3709_/D vssd1 vssd1 vccd1 vccd1 _3709_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_52_wb_clk_i clkbuf_leaf_5_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3666_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_78_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2613__A1 _3193_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3 hold3/A vssd1 vssd1 vccd1 vccd1 hold3/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2040_ hold489/X _2731_/A2 _2867_/A _2034_/X vssd1 vssd1 vccd1 vccd1 _2040_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_84_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2942_ hold888/X _2941_/X _2948_/B vssd1 vssd1 vccd1 vccd1 _2942_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_72_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2873_ _2797_/A _2872_/X _2862_/X vssd1 vssd1 vccd1 vccd1 _2873_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_4_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1824_ _1824_/A _1824_/B _3045_/B _2042_/D vssd1 vssd1 vccd1 vccd1 _2028_/S sky130_fd_sc_hd__or4_4
XANTENNA__2368__A0 _3195_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1755_ _2479_/A _1755_/B vssd1 vssd1 vccd1 vccd1 _1755_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_13_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xmax_cap100 _2083_/Y vssd1 vssd1 vccd1 vccd1 _2099_/B1 sky130_fd_sc_hd__buf_4
XFILLER_0_40_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold425 _3503_/Q vssd1 vssd1 vccd1 vccd1 hold425/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold414 _2256_/X vssd1 vssd1 vccd1 vccd1 _3282_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold436 _2991_/X vssd1 vssd1 vccd1 vccd1 _3666_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold403 _3259_/Q vssd1 vssd1 vccd1 vccd1 hold403/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold469 _3368_/Q vssd1 vssd1 vccd1 vccd1 hold469/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold458 _2208_/X vssd1 vssd1 vccd1 vccd1 _3248_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1686_ _1684_/X _1685_/Y _2961_/A vssd1 vssd1 vccd1 vccd1 _3310_/D sky130_fd_sc_hd__a21o_1
Xhold447 _3647_/Q vssd1 vssd1 vccd1 vccd1 hold447/X sky130_fd_sc_hd__dlygate4sd3_1
X_3425_ _3733_/CLK _3425_/D vssd1 vssd1 vccd1 vccd1 _3425_/Q sky130_fd_sc_hd__dfxtp_1
X_3356_ _3583_/CLK _3356_/D vssd1 vssd1 vccd1 vccd1 _3356_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2307_ _3014_/A _3045_/A _2310_/B vssd1 vssd1 vccd1 vccd1 _2308_/C sky130_fd_sc_hd__or3_1
X_3287_ _3387_/CLK _3287_/D vssd1 vssd1 vccd1 vccd1 _3287_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2238_ _2648_/A0 hold591/X _2243_/S vssd1 vssd1 vccd1 vccd1 _2238_/X sky130_fd_sc_hd__mux2_1
X_2169_ _2301_/C _2169_/B vssd1 vssd1 vccd1 vccd1 _3158_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_45_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1954__S _1954_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold981 _3330_/Q vssd1 vssd1 vccd1 vccd1 hold981/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold970 _3094_/X vssd1 vssd1 vccd1 vccd1 _3095_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold992 _3310_/Q vssd1 vssd1 vccd1 vccd1 hold992/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__2086__A _2087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2047__C1 _2495_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3210_ _3666_/CLK _3210_/D vssd1 vssd1 vccd1 vccd1 _3210_/Q sky130_fd_sc_hd__dfxtp_1
X_3141_ _2914_/B _2886_/A _3137_/C vssd1 vssd1 vccd1 vccd1 _3141_/X sky130_fd_sc_hd__a21o_1
X_3072_ _3059_/A _3081_/B _2181_/Y vssd1 vssd1 vccd1 vccd1 _3072_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_82_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2023_ input9/X _2022_/A _1762_/X _2022_/Y vssd1 vssd1 vccd1 vccd1 _2023_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_89_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2589__A0 _2361_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2925_ _2924_/A _2919_/X _2935_/A vssd1 vssd1 vccd1 vccd1 _2925_/Y sky130_fd_sc_hd__o21ai_1
X_2856_ hold793/X _2940_/B2 _2858_/B _2855_/X vssd1 vssd1 vccd1 vccd1 _2856_/X sky130_fd_sc_hd__a211o_1
X_1807_ _2085_/C _1807_/B vssd1 vssd1 vccd1 vccd1 _1807_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__3002__A1 _2854_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold211 _3464_/Q vssd1 vssd1 vccd1 vccd1 hold211/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold200 _2968_/X vssd1 vssd1 vccd1 vccd1 _3643_/D sky130_fd_sc_hd__dlygate4sd3_1
X_2787_ _2690_/X _2771_/B _2691_/X vssd1 vssd1 vccd1 vccd1 _2788_/B sky130_fd_sc_hd__o21a_1
Xhold233 _3425_/Q vssd1 vssd1 vccd1 vccd1 hold233/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold222 _2575_/X vssd1 vssd1 vccd1 vccd1 _3514_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1738_ _3284_/Q _3356_/Q _3368_/Q _3380_/Q _2000_/S0 _2219_/C vssd1 vssd1 vccd1 vccd1
+ _1738_/X sky130_fd_sc_hd__mux4_1
Xhold244 _2561_/X vssd1 vssd1 vccd1 vccd1 _3502_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold277 _3391_/Q vssd1 vssd1 vccd1 vccd1 hold277/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold266 _2539_/X vssd1 vssd1 vccd1 vccd1 _3483_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1669_ _2876_/A _1685_/B vssd1 vssd1 vccd1 vccd1 _2822_/A sky130_fd_sc_hd__nor2_1
Xhold255 _3462_/Q vssd1 vssd1 vccd1 vccd1 hold255/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold288 _2510_/X vssd1 vssd1 vccd1 vccd1 _3458_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold299 _3575_/Q vssd1 vssd1 vccd1 vccd1 hold299/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3408_ _3665_/CLK _3408_/D vssd1 vssd1 vccd1 vccd1 _3408_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3339_ _3739_/CLK _3339_/D vssd1 vssd1 vccd1 vccd1 _3339_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1803__A _2085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2277__C1 _3058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2044__A2 _2731_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2504__A0 _3196_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2035__A2 _2731_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2710_ _2710_/A _2809_/A vssd1 vssd1 vccd1 vccd1 _2710_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_14_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3690_ _3727_/CLK _3690_/D vssd1 vssd1 vccd1 vccd1 _3690_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2641_ hold49/X _3193_/A0 _2646_/S vssd1 vssd1 vccd1 vccd1 hold50/A sky130_fd_sc_hd__mux2_1
XFILLER_0_2_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2572_ _3201_/A1 hold179/X _2576_/S vssd1 vssd1 vccd1 vccd1 _2572_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_50_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1623__A _2195_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3124_ _3124_/A _3124_/B vssd1 vssd1 vccd1 vccd1 _3124_/Y sky130_fd_sc_hd__nor2_1
X_3055_ _3055_/A _3055_/B _3055_/C vssd1 vssd1 vccd1 vccd1 _3055_/X sky130_fd_sc_hd__and3_1
X_2006_ _2006_/A _2006_/B vssd1 vssd1 vccd1 vccd1 _2006_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_77_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout152_A _3172_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2026__A2 _2731_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2908_ _1712_/A _2868_/C _2940_/B2 hold389/X vssd1 vssd1 vccd1 vccd1 _2908_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_0_45_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2839_ _2871_/A _2839_/B vssd1 vssd1 vccd1 vccd1 _2839_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__1880__S1 _2228_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_31_wb_clk_i_A clkbuf_3_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_7_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3496_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__1700__A1 _2876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3205__A1 _2363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3742_ _3743_/CLK _3742_/D vssd1 vssd1 vccd1 vccd1 _3742_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3673_ _3674_/CLK _3673_/D vssd1 vssd1 vccd1 vccd1 _3673_/Q sky130_fd_sc_hd__dfxtp_1
X_2624_ _2097_/X hold581/X _2625_/S vssd1 vssd1 vccd1 vccd1 _2624_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_30_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2192__A1 _2653_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2555_ hold321/X _3198_/A0 _2555_/S vssd1 vssd1 vccd1 vccd1 _2555_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_10_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2486_ hold61/X _2361_/A _2487_/S vssd1 vssd1 vccd1 vccd1 hold62/A sky130_fd_sc_hd__mux2_1
X_3107_ hold785/X _3126_/A _3106_/X vssd1 vssd1 vccd1 vccd1 _3107_/Y sky130_fd_sc_hd__a21oi_1
X_3038_ _3687_/Q _3038_/B vssd1 vssd1 vccd1 vccd1 _3038_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_65_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1962__S _2085_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2359__A _2359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput15 io_in[5] vssd1 vssd1 vccd1 vccd1 _2046_/A sky130_fd_sc_hd__buf_2
XFILLER_0_64_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1844__S1 _2219_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2340_ hold783/X _2349_/S _2339_/X vssd1 vssd1 vccd1 vccd1 _2340_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_20_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2271_ _2022_/A _2245_/C _2355_/A _2270_/X _3058_/A vssd1 vssd1 vccd1 vccd1 _3293_/D
+ sky130_fd_sc_hd__o311a_1
XANTENNA__2229__A2 _1954_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1986_ _3439_/Q _3743_/Q _1988_/S vssd1 vssd1 vccd1 vccd1 _1987_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_7_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3725_ _3725_/CLK _3725_/D vssd1 vssd1 vccd1 vccd1 _3725_/Q sky130_fd_sc_hd__dfxtp_1
X_3656_ _3662_/CLK _3656_/D vssd1 vssd1 vccd1 vccd1 _3656_/Q sky130_fd_sc_hd__dfxtp_1
X_2607_ _2656_/A0 hold465/X _2611_/S vssd1 vssd1 vccd1 vccd1 _2607_/X sky130_fd_sc_hd__mux2_1
X_3587_ _3587_/CLK _3587_/D vssd1 vssd1 vccd1 vccd1 _3587_/Q sky130_fd_sc_hd__dfxtp_1
X_2538_ hold213/X _2643_/A1 _2541_/S vssd1 vssd1 vccd1 vccd1 _2538_/X sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_3_6__f_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2469_ _3203_/A1 hold587/X _2471_/S vssd1 vssd1 vccd1 vccd1 _2469_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2626__B _3199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3050__C1 _3108_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1826__S1 _1981_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3192__B _3192_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2003__S1 _2228_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1840_ _2185_/C _1840_/B vssd1 vssd1 vccd1 vccd1 _1840_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3510_ _3539_/CLK _3510_/D vssd1 vssd1 vccd1 vccd1 _3510_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1771_ _2074_/A _1770_/X _1819_/A vssd1 vssd1 vccd1 vccd1 _1772_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold607 _3660_/Q vssd1 vssd1 vccd1 vccd1 hold607/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold618 _2957_/X vssd1 vssd1 vccd1 vccd1 _3634_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold629 _3397_/Q vssd1 vssd1 vccd1 vccd1 hold629/X sky130_fd_sc_hd__dlygate4sd3_1
X_3441_ _3745_/CLK hold30/X vssd1 vssd1 vccd1 vccd1 hold29/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3372_ _3419_/CLK _3372_/D vssd1 vssd1 vccd1 vccd1 _3372_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2323_ _3096_/A _2323_/B vssd1 vssd1 vccd1 vccd1 _2323_/Y sky130_fd_sc_hd__nand2_1
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2254_ hold185/X _2089_/X _2259_/S vssd1 vssd1 vccd1 vccd1 _2254_/X sky130_fd_sc_hd__mux2_1
X_2185_ _2185_/A _2244_/B _2185_/C _2480_/C vssd1 vssd1 vccd1 vccd1 _3192_/B sky130_fd_sc_hd__or4_4
XANTENNA__2855__C1 _1696_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1969_ _2228_/A _1933_/X _2195_/B vssd1 vssd1 vccd1 vccd1 _1969_/Y sky130_fd_sc_hd__o21ai_1
X_3708_ _3718_/CLK _3708_/D vssd1 vssd1 vccd1 vccd1 _3708_/Q sky130_fd_sc_hd__dfxtp_1
X_3639_ _3676_/CLK _3639_/D vssd1 vssd1 vccd1 vccd1 _3639_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_21_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3558_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_53_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2377__A1 _2652_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1716__A _1760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4 hold4/A vssd1 vssd1 vccd1 vccd1 hold4/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1983__S0 _1760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2981__S _2987_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2941_ _2941_/A _2941_/B _2941_/C vssd1 vssd1 vccd1 vccd1 _2941_/X sky130_fd_sc_hd__and3_1
XFILLER_0_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2872_ _2816_/B _2839_/B _2843_/B _2863_/X _2871_/Y vssd1 vssd1 vccd1 vccd1 _2872_/X
+ sky130_fd_sc_hd__a41o_1
X_1823_ _2496_/C _2955_/A vssd1 vssd1 vccd1 vccd1 _2042_/D sky130_fd_sc_hd__or2_1
XFILLER_0_44_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1754_ _2289_/A _1751_/Y _1753_/Y _2228_/C _1749_/Y vssd1 vssd1 vccd1 vccd1 _1754_/X
+ sky130_fd_sc_hd__a311o_1
Xmax_cap101 _2083_/Y vssd1 vssd1 vccd1 vccd1 _2084_/B sky130_fd_sc_hd__buf_4
Xhold426 _2562_/X vssd1 vssd1 vccd1 vccd1 _3503_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold404 _2224_/X vssd1 vssd1 vccd1 vccd1 _3259_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold415 _3317_/Q vssd1 vssd1 vccd1 vccd1 hold415/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold459 _3250_/Q vssd1 vssd1 vccd1 vccd1 hold459/X sky130_fd_sc_hd__dlygate4sd3_1
X_3424_ _3592_/CLK _3424_/D vssd1 vssd1 vccd1 vccd1 _3424_/Q sky130_fd_sc_hd__dfxtp_1
X_1685_ _2885_/B _1685_/B vssd1 vssd1 vccd1 vccd1 _1685_/Y sky130_fd_sc_hd__nand2_1
Xhold448 _2972_/X vssd1 vssd1 vccd1 vccd1 _3647_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold437 _3298_/Q vssd1 vssd1 vccd1 vccd1 hold437/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3355_ _3585_/CLK _3355_/D vssd1 vssd1 vccd1 vccd1 _3355_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2306_ _3065_/A _3053_/A vssd1 vssd1 vccd1 vccd1 _3097_/C sky130_fd_sc_hd__nand2_1
X_3286_ _3654_/CLK _3286_/D vssd1 vssd1 vccd1 vccd1 _3286_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2540__A1 _3197_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2237_ _2237_/A _2598_/A vssd1 vssd1 vccd1 vccd1 _2243_/S sky130_fd_sc_hd__nand2_2
XFILLER_0_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2168_ _3059_/A _2160_/X _2166_/X _2167_/X _3055_/A vssd1 vssd1 vccd1 vccd1 _2168_/X
+ sky130_fd_sc_hd__o221a_1
X_2099_ hold934/X _2084_/A _2099_/B1 hold925/X vssd1 vssd1 vccd1 vccd1 _2099_/X sky130_fd_sc_hd__a22o_4
XFILLER_0_75_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout95_A _2089_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold982 _3628_/Q vssd1 vssd1 vccd1 vccd1 _2717_/B sky130_fd_sc_hd__clkbuf_2
Xhold960 _3141_/X vssd1 vssd1 vccd1 vccd1 hold960/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold971 _3404_/Q vssd1 vssd1 vccd1 vccd1 hold971/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold993 _2926_/Y vssd1 vssd1 vccd1 vccd1 hold993/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2531__A1 _2357_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1717__S0 _1981_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2976__S _2987_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2522__A1 _2353_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3140_ hold966/X _3131_/X _3139_/X _3166_/C1 vssd1 vssd1 vccd1 vccd1 _3140_/X sky130_fd_sc_hd__o211a_1
X_3071_ hold846/X _3069_/Y _3070_/X _3062_/X _3108_/A vssd1 vssd1 vccd1 vccd1 _3071_/X
+ sky130_fd_sc_hd__a221o_1
X_2022_ _2022_/A _2022_/B _2022_/C vssd1 vssd1 vccd1 vccd1 _2022_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__2286__A0 _2651_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2924_ _2924_/A _2924_/B _2924_/C vssd1 vssd1 vccd1 vccd1 _2941_/C sky130_fd_sc_hd__and3_1
X_2855_ hold908/X _1650_/A _1654_/B _1696_/Y vssd1 vssd1 vccd1 vccd1 _2855_/X sky130_fd_sc_hd__o211a_1
X_1806_ hold3/A _3249_/Q _1937_/S vssd1 vssd1 vccd1 vccd1 _1807_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_31_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2786_ _2786_/A vssd1 vssd1 vccd1 vccd1 _2786_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3002__A2 _1767_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold201 _3493_/Q vssd1 vssd1 vccd1 vccd1 hold201/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold223 _3513_/Q vssd1 vssd1 vccd1 vccd1 hold223/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold234 _2467_/X vssd1 vssd1 vccd1 vccd1 _3425_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1737_ _3544_/Q _3254_/Q _3520_/Q _3508_/Q _2000_/S0 _2219_/C vssd1 vssd1 vccd1 vccd1
+ _1737_/X sky130_fd_sc_hd__mux4_1
Xhold212 _2517_/X vssd1 vssd1 vccd1 vccd1 _3464_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold245 _3476_/Q vssd1 vssd1 vccd1 vccd1 hold245/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold278 _2425_/X vssd1 vssd1 vccd1 vccd1 _3391_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold267 _3424_/Q vssd1 vssd1 vccd1 vccd1 hold267/X sky130_fd_sc_hd__dlygate4sd3_1
X_1668_ _1667_/A _1698_/A _1667_/Y _1824_/A vssd1 vssd1 vccd1 vccd1 _1668_/X sky130_fd_sc_hd__a22o_1
Xhold256 _2515_/X vssd1 vssd1 vccd1 vccd1 _3462_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold289 _3479_/Q vssd1 vssd1 vccd1 vccd1 hold289/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3407_ _3419_/CLK _3407_/D vssd1 vssd1 vccd1 vccd1 _3407_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2513__A1 _2363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1599_ _1599_/A vssd1 vssd1 vccd1 vccd1 _1704_/B sky130_fd_sc_hd__inv_2
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3338_ _3738_/CLK _3338_/D vssd1 vssd1 vccd1 vccd1 _3338_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3269_ _3270_/CLK _3269_/D vssd1 vssd1 vccd1 vccd1 _3269_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2201__A0 _2659_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_21_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_31_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold790 _2390_/X vssd1 vssd1 vccd1 vccd1 _3361_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2640_ _2640_/A _2640_/B vssd1 vssd1 vccd1 vccd1 _2646_/S sky130_fd_sc_hd__nor2_2
XANTENNA__2991__A1 _2228_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2571_ _2353_/A hold445/X _2576_/S vssd1 vssd1 vccd1 vccd1 _2571_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_22_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1929__S0 _1981_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1703__C1 _2961_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3123_ hold809/X _3120_/A _3122_/X _3055_/A vssd1 vssd1 vccd1 vccd1 _3123_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_89_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3054_ _3054_/A _3054_/B vssd1 vssd1 vccd1 vccd1 _3055_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_77_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2005_ _3343_/Q _3301_/Q _2005_/S vssd1 vssd1 vccd1 vccd1 _2006_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_92_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2907_ _2904_/A _2944_/B _2906_/Y _3166_/C1 vssd1 vssd1 vccd1 vccd1 _2907_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_42_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2838_ hold950/X _2824_/X _2836_/X _2837_/X _2859_/A vssd1 vssd1 vccd1 vccd1 _2838_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_13_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2769_ _2769_/A vssd1 vssd1 vccd1 vccd1 _2769_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2498__A0 _2074_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1708__B _3048_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1724__A _2006_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2489__A0 _2648_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3741_ _3741_/CLK _3741_/D vssd1 vssd1 vccd1 vccd1 _3741_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2413__A0 _2660_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3672_ _3672_/CLK _3672_/D vssd1 vssd1 vccd1 vccd1 _3672_/Q sky130_fd_sc_hd__dfxtp_1
X_2623_ _2658_/A0 hold711/X _2625_/S vssd1 vssd1 vccd1 vccd1 _2623_/X sky130_fd_sc_hd__mux2_1
X_2554_ hold219/X _2659_/A0 _2555_/S vssd1 vssd1 vccd1 vccd1 _2554_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_50_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2485_ hold253/X _3203_/A1 _2487_/S vssd1 vssd1 vccd1 vccd1 _2485_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_10_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3106_ _3013_/Y _3118_/B _3120_/A _3183_/B vssd1 vssd1 vccd1 vccd1 _3106_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_37_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2465__A _2598_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3037_ _3065_/A _3097_/A _3037_/C _3037_/D vssd1 vssd1 vccd1 vccd1 _3038_/B sky130_fd_sc_hd__or4_1
XFILLER_0_77_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2652__A0 _2652_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2404__A0 _3196_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_46_wb_clk_i clkbuf_3_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3714_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_5_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2168__C1 _3055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1710__C _3045_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput16 io_in[6] vssd1 vssd1 vccd1 vccd1 _2050_/A sky130_fd_sc_hd__buf_2
XFILLER_0_24_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2270_ _2270_/A _2278_/B vssd1 vssd1 vccd1 vccd1 _2270_/X sky130_fd_sc_hd__or2_1
XANTENNA__2984__S _2987_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2882__B1 _2876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2229__A3 _2014_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2634__A0 _2655_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1985_ _3501_/Q _3513_/Q _3525_/Q _3537_/Q _1988_/S _2185_/C vssd1 vssd1 vccd1 vccd1
+ _1985_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_7_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3724_ _3724_/CLK _3724_/D vssd1 vssd1 vccd1 vccd1 _3724_/Q sky130_fd_sc_hd__dfxtp_1
X_3655_ _3655_/CLK _3655_/D vssd1 vssd1 vccd1 vccd1 _3655_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2606_ _2655_/A0 hold671/X _2611_/S vssd1 vssd1 vccd1 vccd1 _2606_/X sky130_fd_sc_hd__mux2_1
X_3586_ _3586_/CLK _3586_/D vssd1 vssd1 vccd1 vccd1 _3586_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2537_ hold67/X _3194_/A0 _2541_/S vssd1 vssd1 vccd1 vccd1 hold68/A sky130_fd_sc_hd__mux2_1
X_2468_ _2650_/A0 hold231/X _2471_/S vssd1 vssd1 vccd1 vccd1 _2468_/X sky130_fd_sc_hd__mux2_1
X_2399_ _2660_/A0 hold477/X _2399_/S vssd1 vssd1 vccd1 vccd1 _2399_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2195__A _2479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2625__A0 _2660_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2928__B2 _2940_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2928__A1 _1712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2092__A1 _2091_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3041__B1 _3055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1770_ _2854_/B _1768_/X _1769_/Y _2998_/A1 vssd1 vssd1 vccd1 vccd1 _1770_/X sky130_fd_sc_hd__o22a_1
XANTENNA__2979__S _2987_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold608 _2985_/X vssd1 vssd1 vccd1 vccd1 _3660_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold619 _3571_/Q vssd1 vssd1 vccd1 vccd1 hold619/X sky130_fd_sc_hd__dlygate4sd3_1
X_3440_ _3744_/CLK hold62/X vssd1 vssd1 vccd1 vccd1 hold61/A sky130_fd_sc_hd__dfxtp_1
X_3371_ _3419_/CLK _3371_/D vssd1 vssd1 vccd1 vccd1 _3371_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2322_ _3705_/Q _3089_/B _2321_/X _2303_/A vssd1 vssd1 vccd1 vccd1 _2323_/B sky130_fd_sc_hd__a211o_1
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2253_ _3192_/B _2640_/B vssd1 vssd1 vccd1 vccd1 _2259_/S sky130_fd_sc_hd__nor2_4
XANTENNA__1912__A _2085_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2184_ _2182_/A _3157_/B _2166_/X _2183_/X _3055_/A vssd1 vssd1 vccd1 vccd1 _2184_/X
+ sky130_fd_sc_hd__o221a_1
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
XANTENNA__2607__A0 _2656_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1968_ _2479_/A _1940_/X _1947_/X _1967_/Y vssd1 vssd1 vccd1 vccd1 _1971_/B sky130_fd_sc_hd__a31o_1
X_1899_ _1898_/X _1897_/X _1895_/X _1896_/X _2289_/A _2479_/B vssd1 vssd1 vccd1 vccd1
+ _1899_/X sky130_fd_sc_hd__mux4_1
X_3707_ _3718_/CLK _3707_/D vssd1 vssd1 vccd1 vccd1 _3707_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3638_ _3668_/CLK hold40/X vssd1 vssd1 vccd1 vccd1 hold39/A sky130_fd_sc_hd__dfxtp_1
X_3569_ _3587_/CLK _3569_/D vssd1 vssd1 vccd1 vccd1 _3569_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1992__S1 _2185_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2372__B _2612_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1716__B _1760_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1732__A _2185_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1983__S1 _1760_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold5 hold5/A vssd1 vssd1 vccd1 vccd1 hold5/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2837__B1 _2940_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output21_A _3770_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2940_ _1712_/A _2998_/A1 hold447/X _2940_/B2 vssd1 vssd1 vccd1 vccd1 _2940_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_29_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2065__B2 _2868_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2871_ _2871_/A _2871_/B vssd1 vssd1 vccd1 vccd1 _2871_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_29_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1822_ _2153_/A _2301_/C _1821_/X vssd1 vssd1 vccd1 vccd1 _2955_/A sky130_fd_sc_hd__or3b_4
XFILLER_0_44_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1753_ _2085_/C _1753_/B vssd1 vssd1 vccd1 vccd1 _1753_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_4_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold427 _3507_/Q vssd1 vssd1 vccd1 vccd1 hold427/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1684_ _2797_/A _1683_/Y _1685_/B _2080_/A vssd1 vssd1 vccd1 vccd1 _1684_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_20_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold405 _3291_/Q vssd1 vssd1 vccd1 vccd1 hold405/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold416 _2333_/X vssd1 vssd1 vccd1 vccd1 _3317_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3423_ _3665_/CLK _3423_/D vssd1 vssd1 vccd1 vccd1 _3423_/Q sky130_fd_sc_hd__dfxtp_1
Xhold449 _3443_/Q vssd1 vssd1 vccd1 vccd1 hold449/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold438 _2283_/X vssd1 vssd1 vccd1 vccd1 _3298_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3354_ _3585_/CLK _3354_/D vssd1 vssd1 vccd1 vccd1 _3354_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3285_ _3583_/CLK _3285_/D vssd1 vssd1 vccd1 vccd1 _3285_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2305_ _2305_/A _3053_/A _3097_/B vssd1 vssd1 vccd1 vccd1 _2311_/C sky130_fd_sc_hd__or3_1
XANTENNA__1642__A _2885_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2236_ _3198_/A0 hold689/X _2236_/S vssd1 vssd1 vccd1 vccd1 _2236_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2167_ _3045_/B _2167_/B _2167_/C vssd1 vssd1 vccd1 vccd1 _2167_/X sky130_fd_sc_hd__or3_1
XFILLER_0_45_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2098_ hold311/X _3197_/A0 _2100_/S vssd1 vssd1 vccd1 vccd1 _2098_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_48_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_11_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_90_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold950 _3603_/Q vssd1 vssd1 vccd1 vccd1 hold950/X sky130_fd_sc_hd__buf_1
Xhold961 _3142_/X vssd1 vssd1 vccd1 vccd1 _3707_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold972 _3629_/Q vssd1 vssd1 vccd1 vccd1 _2854_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold994 _3329_/Q vssd1 vssd1 vccd1 vccd1 hold994/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold983 _2060_/X vssd1 vssd1 vccd1 vccd1 hold983/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout88_A _2091_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1717__S1 _1981_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2295__A1 _2652_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2086__C _2480_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_50_wb_clk_i_A clkbuf_3_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_39_423 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3180__C1 _3058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3070_ _3228_/Q _3048_/B _3096_/C _3068_/Y vssd1 vssd1 vccd1 vccd1 _3070_/X sky130_fd_sc_hd__o31a_1
X_2021_ _2228_/A _2010_/X _2017_/X _2020_/Y vssd1 vssd1 vccd1 vccd1 _2022_/C sky130_fd_sc_hd__a31o_1
XFILLER_0_57_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2923_ _1712_/A _3607_/Q hold297/X _2940_/B2 vssd1 vssd1 vccd1 vccd1 _2923_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_0_17_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2854_ _2854_/A _2854_/B _2825_/A _2822_/B vssd1 vssd1 vccd1 vccd1 _2858_/B sky130_fd_sc_hd__or4bb_1
X_1805_ _2245_/B _1805_/B vssd1 vssd1 vccd1 vccd1 _1805_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_60_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2785_ _2868_/C _2861_/B _2812_/S vssd1 vssd1 vccd1 vccd1 _2786_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_32_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1736_ _3392_/Q _3586_/Q _3568_/Q _3556_/Q _2000_/S0 _2219_/C vssd1 vssd1 vccd1 vccd1
+ _1736_/X sky130_fd_sc_hd__mux4_1
Xhold202 _2551_/X vssd1 vssd1 vccd1 vccd1 _3493_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold224 _2574_/X vssd1 vssd1 vccd1 vccd1 _3513_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold235 _3500_/Q vssd1 vssd1 vccd1 vccd1 hold235/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold213 _3482_/Q vssd1 vssd1 vccd1 vccd1 hold213/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold246 _2531_/X vssd1 vssd1 vccd1 vccd1 _3476_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold257 _3252_/Q vssd1 vssd1 vccd1 vccd1 hold257/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold268 _2466_/X vssd1 vssd1 vccd1 vccd1 _3424_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1667_ _1667_/A _2846_/B _2876_/C vssd1 vssd1 vccd1 vccd1 _1667_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_13_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3406_ _3665_/CLK _3406_/D vssd1 vssd1 vccd1 vccd1 _3406_/Q sky130_fd_sc_hd__dfxtp_1
Xhold279 _3257_/Q vssd1 vssd1 vccd1 vccd1 hold279/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3337_ _3738_/CLK _3337_/D vssd1 vssd1 vccd1 vccd1 _3337_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3268_ _3270_/CLK _3268_/D vssd1 vssd1 vccd1 vccd1 _3268_/Q sky130_fd_sc_hd__dfxtp_1
X_3199_ _3199_/A _3199_/B vssd1 vssd1 vccd1 vccd1 _3205_/S sky130_fd_sc_hd__nor2_2
X_2219_ _2000_/S0 _2480_/C _2219_/C _3348_/Q vssd1 vssd1 vccd1 vccd1 _2647_/A sky130_fd_sc_hd__and4bb_4
XANTENNA__2277__A1 _1716_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1788__B1 _3348_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold791 _3526_/Q vssd1 vssd1 vccd1 vccd1 hold791/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold780 _2620_/X vssd1 vssd1 vccd1 vccd1 _3552_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_6_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2440__A1 _2650_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2570_ _2570_/A _2598_/B vssd1 vssd1 vccd1 vccd1 _2576_/S sky130_fd_sc_hd__nand2_4
XANTENNA__2987__S _2987_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1929__S1 _1981_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3122_ _3699_/Q _3118_/A _3126_/A _3115_/X vssd1 vssd1 vccd1 vccd1 _3122_/X sky130_fd_sc_hd__a211o_1
XANTENNA__2259__A1 _2660_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3053_ _3053_/A _3053_/B _3053_/C vssd1 vssd1 vccd1 vccd1 _3054_/B sky130_fd_sc_hd__and3_1
X_2004_ _3295_/Q _3445_/Q _3579_/Q _3403_/Q _1954_/S _2014_/A vssd1 vssd1 vccd1 vccd1
+ _2004_/X sky130_fd_sc_hd__mux4_1
XANTENNA__1920__A input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2431__A1 _2353_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2906_ _2876_/A _2902_/Y _2905_/X _2883_/Y vssd1 vssd1 vccd1 vccd1 _2906_/Y sky130_fd_sc_hd__o211ai_1
XANTENNA_fanout138_A _1954_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2837_ _2861_/B _1696_/Y _2940_/B2 hold607/X _2825_/Y vssd1 vssd1 vccd1 vccd1 _2837_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_60_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2768_ _2867_/C hold893/X _2812_/S vssd1 vssd1 vccd1 vccd1 _2769_/A sky130_fd_sc_hd__mux2_1
X_2699_ _2698_/B _2698_/C _2802_/A vssd1 vssd1 vccd1 vccd1 _2803_/C sky130_fd_sc_hd__o21ai_2
X_1719_ _3496_/Q hold95/A _3466_/Q _3454_/Q _1981_/S0 _1981_/S1 vssd1 vssd1 vccd1
+ vccd1 _1719_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_6_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2661__A _3199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2422__A1 _2655_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1856__S0 _2085_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2110__A0 _3197_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3740_ _3743_/CLK _3740_/D vssd1 vssd1 vccd1 vccd1 _3740_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3671_ _3672_/CLK _3671_/D vssd1 vssd1 vccd1 vccd1 _3671_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2290__B _2612_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2622_ _3195_/A0 hold731/X _2625_/S vssd1 vssd1 vccd1 vccd1 _2622_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_10_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2553_ hold13/X _3196_/A0 _2555_/S vssd1 vssd1 vccd1 vccd1 hold14/A sky130_fd_sc_hd__mux2_1
XFILLER_0_10_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2484_ hold69/X _2357_/A _2487_/S vssd1 vssd1 vccd1 vccd1 hold70/A sky130_fd_sc_hd__mux2_1
XFILLER_0_10_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3105_ _3677_/Q _3004_/Y _3023_/B vssd1 vssd1 vccd1 vccd1 _3126_/A sky130_fd_sc_hd__o21ai_4
X_3036_ _3086_/A _3036_/B _3036_/C vssd1 vssd1 vccd1 vccd1 _3036_/X sky130_fd_sc_hd__and3_1
XFILLER_0_77_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2481__A _2612_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3117__C1 _3055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_15_wb_clk_i clkbuf_3_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3583_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_68_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1829__S0 _2085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput17 io_in[9] vssd1 vssd1 vccd1 vccd1 _1626_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_91_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output51_A _3612_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2398__A0 _2659_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1984_ _1982_/X _1983_/X _1981_/X _1980_/X _2085_/A _2228_/C vssd1 vssd1 vccd1 vccd1
+ _1984_/X sky130_fd_sc_hd__mux4_1
X_3723_ _3723_/CLK _3723_/D vssd1 vssd1 vccd1 vccd1 _3723_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3654_ _3654_/CLK _3654_/D vssd1 vssd1 vccd1 vccd1 _3654_/Q sky130_fd_sc_hd__dfxtp_1
X_2605_ _3192_/B _2633_/B vssd1 vssd1 vccd1 vccd1 _2611_/S sky130_fd_sc_hd__or2_4
XFILLER_0_30_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3585_ _3585_/CLK _3585_/D vssd1 vssd1 vccd1 vccd1 _3585_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2536_ hold159/X _2655_/A0 _2541_/S vssd1 vssd1 vccd1 vccd1 _2536_/X sky130_fd_sc_hd__mux2_1
X_2467_ _3201_/A1 hold233/X _2471_/S vssd1 vssd1 vccd1 vccd1 _2467_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2398_ _2659_/A0 hold469/X _2399_/S vssd1 vssd1 vccd1 vccd1 _2398_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2873__A1 _2797_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2195__B _2195_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3019_ _3037_/C _3018_/X _3118_/B vssd1 vssd1 vccd1 vccd1 _3019_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__2389__A0 _2475_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3770__A _3770_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout150 _2495_/A vssd1 vssd1 vccd1 vccd1 _2859_/A sky130_fd_sc_hd__buf_4
XANTENNA__2864__A1 _3594_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2386__A _2640_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2616__A1 _2359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2077__C1 _2495_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold609 _3217_/Q vssd1 vssd1 vccd1 vccd1 hold609/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3370_ _3654_/CLK _3370_/D vssd1 vssd1 vccd1 vccd1 _3370_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2321_ _3709_/Q _2313_/X _2316_/Y hold838/X vssd1 vssd1 vccd1 vccd1 _2321_/X sky130_fd_sc_hd__a22o_1
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2252_ hold65/X _2653_/A0 _2252_/S vssd1 vssd1 vccd1 vccd1 hold66/A sky130_fd_sc_hd__mux2_1
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_52 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2855__A1 hold908/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2183_ _2173_/Y _2181_/Y _2182_/X _2169_/B vssd1 vssd1 vccd1 vccd1 _2183_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_62_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1967_ _2479_/A _1952_/X _2228_/B vssd1 vssd1 vccd1 vccd1 _1967_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout120_A _3349_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3706_ _3718_/CLK _3706_/D vssd1 vssd1 vccd1 vccd1 _3706_/Q sky130_fd_sc_hd__dfxtp_1
X_1898_ _3547_/Q _3559_/Q _3571_/Q _3236_/Q _2289_/B _2289_/C vssd1 vssd1 vccd1 vccd1
+ _1898_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_43_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3637_ _3637_/CLK _3637_/D vssd1 vssd1 vccd1 vccd1 _3637_/Q sky130_fd_sc_hd__dfxtp_1
X_3568_ _3587_/CLK _3568_/D vssd1 vssd1 vccd1 vccd1 _3568_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2543__A0 _2353_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2519_ hold101/X _3197_/A0 _2520_/S vssd1 vssd1 vccd1 vccd1 _2519_/X sky130_fd_sc_hd__mux2_1
X_3499_ _3539_/CLK _3499_/D vssd1 vssd1 vccd1 vccd1 _3499_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2059__C1 _1979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_40_wb_clk_i_A clkbuf_3_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_19_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_30_wb_clk_i clkbuf_3_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3592_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold6 hold6/A vssd1 vssd1 vccd1 vccd1 hold6/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_71_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2563__B _2598_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2065__A2 _2731_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2870_ _2864_/X _2865_/Y _2869_/X hold860/X vssd1 vssd1 vccd1 vccd1 _2871_/B sky130_fd_sc_hd__o22a_1
XFILLER_0_72_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1821_ _2182_/A _3059_/B _2316_/A vssd1 vssd1 vccd1 vccd1 _1821_/X sky130_fd_sc_hd__and3_2
XFILLER_0_44_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1752_ _3233_/Q _3248_/Q _1937_/S vssd1 vssd1 vccd1 vccd1 _1753_/B sky130_fd_sc_hd__mux2_1
X_1683_ _1667_/Y _1683_/B vssd1 vssd1 vccd1 vccd1 _1683_/Y sky130_fd_sc_hd__nand2b_1
Xhold417 _3667_/Q vssd1 vssd1 vccd1 vccd1 hold417/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold406 _2266_/X vssd1 vssd1 vccd1 vccd1 _3291_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold439 _3489_/Q vssd1 vssd1 vccd1 vccd1 hold439/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold428 _2567_/X vssd1 vssd1 vccd1 vccd1 _3507_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3422_ _3665_/CLK _3422_/D vssd1 vssd1 vccd1 vccd1 _3422_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3353_ _3583_/CLK _3353_/D vssd1 vssd1 vccd1 vccd1 _3353_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3284_ _3583_/CLK _3284_/D vssd1 vssd1 vccd1 vccd1 _3284_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2304_ _3688_/Q _3687_/Q _3097_/A _3097_/B vssd1 vssd1 vccd1 vccd1 _2304_/X sky130_fd_sc_hd__or4_1
XFILLER_0_29_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2828__A1 hold918/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1642__B _2797_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2235_ _3197_/A0 hold339/X _2236_/S vssd1 vssd1 vccd1 vccd1 _2235_/X sky130_fd_sc_hd__mux2_1
X_2166_ _2164_/X _2165_/X _2166_/C _2166_/D vssd1 vssd1 vccd1 vccd1 _2166_/X sky130_fd_sc_hd__and4bb_2
X_2097_ _2861_/B _2084_/A _2099_/B1 hold852/X vssd1 vssd1 vccd1 vccd1 _2097_/X sky130_fd_sc_hd__a22o_2
XFILLER_0_48_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2999_ hold375/X _2999_/A1 _2999_/S vssd1 vssd1 vccd1 vccd1 _2999_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_9_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold940 _3003_/Y vssd1 vssd1 vccd1 vccd1 _3676_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_7_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold962 _3332_/Q vssd1 vssd1 vccd1 vccd1 hold962/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold951 _2838_/X vssd1 vssd1 vccd1 vccd1 _3603_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold973 _2062_/X vssd1 vssd1 vccd1 vccd1 hold973/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold995 _3333_/Q vssd1 vssd1 vccd1 vccd1 hold995/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold984 _2061_/X vssd1 vssd1 vccd1 vccd1 _3628_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1743__A _2085_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2020_ _2228_/A _1984_/X _2195_/B vssd1 vssd1 vccd1 vccd1 _2020_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_89_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2922_ _2924_/B _2883_/Y _2921_/Y _3103_/A vssd1 vssd1 vccd1 vccd1 _2922_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_57_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2853_ _2718_/B _2849_/Y _2852_/X vssd1 vssd1 vccd1 vccd1 _2853_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_31_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1804_ _3261_/Q _3273_/Q _1937_/S vssd1 vssd1 vccd1 vccd1 _1805_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_60_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2784_ hold893/X _2730_/Y _2782_/Y _2783_/X _2859_/A vssd1 vssd1 vccd1 vccd1 _2784_/X
+ sky130_fd_sc_hd__o221a_1
X_1735_ _1889_/A _1732_/Y _1734_/Y _2428_/C _1730_/Y vssd1 vssd1 vccd1 vccd1 _1735_/X
+ sky130_fd_sc_hd__a311o_1
Xhold203 _3590_/Q vssd1 vssd1 vccd1 vccd1 hold203/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold214 _2538_/X vssd1 vssd1 vccd1 vccd1 _3482_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold225 _3442_/Q vssd1 vssd1 vccd1 vccd1 hold225/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold247 _3566_/Q vssd1 vssd1 vccd1 vccd1 hold247/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold258 _2215_/X vssd1 vssd1 vccd1 vccd1 _3252_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold236 _2559_/X vssd1 vssd1 vccd1 vccd1 _3500_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold269 _3740_/Q vssd1 vssd1 vccd1 vccd1 hold269/X sky130_fd_sc_hd__dlygate4sd3_1
X_1666_ _2868_/B _1673_/C vssd1 vssd1 vccd1 vccd1 _2876_/C sky130_fd_sc_hd__or2_1
XFILLER_0_21_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3405_ _3725_/CLK _3405_/D vssd1 vssd1 vccd1 vccd1 _3405_/Q sky130_fd_sc_hd__dfxtp_1
X_3336_ _3739_/CLK _3336_/D vssd1 vssd1 vccd1 vccd1 _3336_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3267_ _3419_/CLK _3267_/D vssd1 vssd1 vccd1 vccd1 _3267_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2218_ _2660_/A0 hold567/X _2218_/S vssd1 vssd1 vccd1 vccd1 _2218_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2277__A2 _2245_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3198_ _3198_/A0 hold523/X _3198_/S vssd1 vssd1 vccd1 vccd1 _3198_/X sky130_fd_sc_hd__mux2_1
X_2149_ _3705_/Q _2149_/B _2149_/C vssd1 vssd1 vccd1 vccd1 _2149_/Y sky130_fd_sc_hd__nor3_1
XANTENNA__1788__A1 _2006_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold770 _2587_/X vssd1 vssd1 vccd1 vccd1 _3524_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold781 _3407_/Q vssd1 vssd1 vccd1 vccd1 hold781/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold792 _2589_/X vssd1 vssd1 vccd1 vccd1 _3526_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2728__A0 _2701_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1703__B2 _2960_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3121_ hold821/X _3120_/A _3120_/Y _3055_/A vssd1 vssd1 vccd1 vccd1 _3121_/X sky130_fd_sc_hd__o211a_1
X_3052_ _3053_/B _3048_/X _3053_/A vssd1 vssd1 vccd1 vccd1 _3052_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_89_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2003_ _2002_/X _2001_/X _1999_/X _2000_/X _2289_/A _2228_/C vssd1 vssd1 vccd1 vccd1
+ _2003_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2905_ _2948_/B _2914_/C _2904_/X vssd1 vssd1 vccd1 vccd1 _2905_/X sky130_fd_sc_hd__or3b_1
X_2836_ hold893/X _2871_/A _2835_/Y _2876_/B vssd1 vssd1 vccd1 vccd1 _2836_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_60_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2767_ hold923/X _2730_/Y _2765_/Y _2766_/X _2859_/A vssd1 vssd1 vccd1 vccd1 _2767_/X
+ sky130_fd_sc_hd__o221a_1
X_2698_ _2802_/A _2698_/B _2698_/C vssd1 vssd1 vccd1 vccd1 _2803_/B sky130_fd_sc_hd__or3_1
X_1718_ _3386_/Q _3374_/Q _3362_/Q _3290_/Q _1981_/S0 _1981_/S1 vssd1 vssd1 vccd1
+ vccd1 _1718_/X sky130_fd_sc_hd__mux4_1
XANTENNA__2479__A _2479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1649_ _3630_/Q _1663_/B _1713_/B vssd1 vssd1 vccd1 vccd1 _1701_/A sky130_fd_sc_hd__nor3_1
XANTENNA_hold1050_A _3613_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3319_ _3738_/CLK _3319_/D vssd1 vssd1 vccd1 vccd1 _3319_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3103__A _3103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2958__A0 _2046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1856__S1 _2014_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3773__A _3773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1697__B1 _1696_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2894__C1 _2859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1792__S0 _2000_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3071__C1 _3108_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3670_ _3670_/CLK _3670_/D vssd1 vssd1 vccd1 vccd1 _3670_/Q sky130_fd_sc_hd__dfxtp_1
X_2621_ _2656_/A0 hold703/X _2625_/S vssd1 vssd1 vccd1 vccd1 _2621_/X sky130_fd_sc_hd__mux2_1
X_2552_ hold119/X _2643_/A1 _2555_/S vssd1 vssd1 vccd1 vccd1 _2552_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_23_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2483_ hold53/X _2355_/A _2487_/S vssd1 vssd1 vccd1 vccd1 hold54/A sky130_fd_sc_hd__mux2_1
X_3104_ _3677_/Q _3004_/Y _3023_/B vssd1 vssd1 vccd1 vccd1 _3120_/A sky130_fd_sc_hd__o21a_2
X_3035_ _3035_/A _3035_/B vssd1 vssd1 vccd1 vccd1 _3036_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout150_A _2495_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_279 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2819_ _2819_/A _2876_/C vssd1 vssd1 vccd1 vccd1 _2819_/X sky130_fd_sc_hd__and2_1
XANTENNA__1915__A1 _2479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1774__S0 _1981_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_55_wb_clk_i clkbuf_leaf_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3670_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__3768__A _3768_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1829__S1 _2228_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput18 rst_n vssd1 vssd1 vccd1 vccd1 input18/X sky130_fd_sc_hd__buf_2
XANTENNA_hold996_A _3612_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1906__A1 _2244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1751__A _2245_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1983_ _3433_/Q _3421_/Q _3409_/Q _3265_/Q _1760_/A _1760_/B vssd1 vssd1 vccd1 vccd1
+ _1983_/X sky130_fd_sc_hd__mux4_1
X_3722_ _3723_/CLK _3722_/D vssd1 vssd1 vccd1 vccd1 _3722_/Q sky130_fd_sc_hd__dfxtp_1
X_3653_ _3655_/CLK _3653_/D vssd1 vssd1 vccd1 vccd1 _3653_/Q sky130_fd_sc_hd__dfxtp_1
X_2604_ _2363_/A hold613/X _2604_/S vssd1 vssd1 vccd1 vccd1 _2604_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_70_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3584_ _3586_/CLK _3584_/D vssd1 vssd1 vccd1 vccd1 _3584_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2535_ _2549_/A _3199_/A vssd1 vssd1 vccd1 vccd1 _2541_/S sky130_fd_sc_hd__nor2_4
X_2466_ _2648_/A0 hold267/X _2471_/S vssd1 vssd1 vccd1 vccd1 _2466_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_48_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2397_ _2658_/A0 hold545/X _2399_/S vssd1 vssd1 vccd1 vccd1 _2397_/X sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_30_wb_clk_i_A clkbuf_3_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__2195__C _2479_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3018_ _3124_/A _3063_/B _3682_/Q vssd1 vssd1 vccd1 vccd1 _3018_/X sky130_fd_sc_hd__or3b_1
XFILLER_0_78_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2561__A1 _2361_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout140 _1988_/S vssd1 vssd1 vccd1 vccd1 _1937_/S sky130_fd_sc_hd__clkbuf_8
Xfanout151 input18/X vssd1 vssd1 vccd1 vccd1 _2495_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_84_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2320_ _3055_/A _2320_/B _2320_/C vssd1 vssd1 vccd1 vccd1 _2320_/X sky130_fd_sc_hd__and3_1
XFILLER_0_20_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2251_ hold1/X _2652_/A0 _2252_/S vssd1 vssd1 vccd1 vccd1 hold2/A sky130_fd_sc_hd__mux2_1
XANTENNA__1738__S0 _2000_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2182_ _2182_/A _2182_/B vssd1 vssd1 vccd1 vccd1 _2182_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_0_wb_clk_i clkbuf_leaf_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3661_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_1966_ _2085_/A _1963_/Y _1965_/Y _2087_/A _1961_/Y vssd1 vssd1 vccd1 vccd1 _1966_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_0_83_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3705_ _3718_/CLK _3705_/D vssd1 vssd1 vccd1 vccd1 _3705_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2240__A0 _2357_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1897_ _3281_/Q _3353_/Q _3365_/Q _3377_/Q _2000_/S0 _2219_/C vssd1 vssd1 vccd1 vccd1
+ _1897_/X sky130_fd_sc_hd__mux4_1
X_3636_ _3636_/CLK _3636_/D vssd1 vssd1 vccd1 vccd1 _3636_/Q sky130_fd_sc_hd__dfxtp_1
X_3567_ _3583_/CLK _3567_/D vssd1 vssd1 vccd1 vccd1 _3567_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2518_ hold485/X _3196_/A0 _2520_/S vssd1 vssd1 vccd1 vccd1 _2518_/X sky130_fd_sc_hd__mux2_1
X_3498_ _3743_/CLK _3498_/D vssd1 vssd1 vccd1 vccd1 _3498_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1729__S0 _2244_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3099__A2 _3048_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2449_ _3197_/A0 hold549/X _2450_/S vssd1 vssd1 vccd1 vccd1 _2449_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_66_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2231__A0 _3193_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2534__A1 _2363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold7 hold7/A vssd1 vssd1 vccd1 vccd1 hold7/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2837__A2 _1696_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2470__A0 _2652_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1820_ _2076_/A _1819_/A _1819_/Y _1979_/A vssd1 vssd1 vccd1 vccd1 _1820_/X sky130_fd_sc_hd__o211a_1
XANTENNA__2222__A0 _2355_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1751_ _2245_/B _1751_/B vssd1 vssd1 vccd1 vccd1 _1751_/Y sky130_fd_sc_hd__nand2_1
X_1682_ _2960_/A _1642_/X _1668_/X _1681_/X _1824_/A vssd1 vssd1 vccd1 vccd1 _1682_/X
+ sky130_fd_sc_hd__a32o_1
Xhold407 _3651_/Q vssd1 vssd1 vccd1 vccd1 hold407/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold418 _2992_/X vssd1 vssd1 vccd1 vccd1 _3667_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold429 _3515_/Q vssd1 vssd1 vccd1 vccd1 hold429/X sky130_fd_sc_hd__dlygate4sd3_1
X_3421_ _3665_/CLK _3421_/D vssd1 vssd1 vccd1 vccd1 _3421_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2525__A1 _3203_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3352_ _3575_/CLK _3352_/D vssd1 vssd1 vccd1 vccd1 _3352_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2303_ _2303_/A _3089_/A _2316_/B vssd1 vssd1 vccd1 vccd1 _2303_/X sky130_fd_sc_hd__or3b_2
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3283_ _3585_/CLK _3283_/D vssd1 vssd1 vccd1 vccd1 _3283_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1642__C _1979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2234_ _3196_/A0 hold513/X _2236_/S vssd1 vssd1 vccd1 vccd1 _2234_/X sky130_fd_sc_hd__mux2_1
X_2165_ _2131_/X _2132_/X _2153_/Y vssd1 vssd1 vccd1 vccd1 _2165_/X sky130_fd_sc_hd__a21bo_1
X_2096_ hold85/X _2651_/A0 _2100_/S vssd1 vssd1 vccd1 vccd1 hold86/A sky130_fd_sc_hd__mux2_1
XFILLER_0_45_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2461__A0 _2475_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2213__A0 _2655_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2998_ hold767/X _2998_/A1 _2999_/S vssd1 vssd1 vccd1 vccd1 _2998_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_16_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1949_ _3542_/Q _3252_/Q _3518_/Q _3506_/Q _2000_/S0 _2219_/C vssd1 vssd1 vccd1 vccd1
+ _1949_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_43_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3619_ _3672_/CLK _3619_/D vssd1 vssd1 vccd1 vccd1 _3619_/Q sky130_fd_sc_hd__dfxtp_1
Xhold930 _3033_/Y vssd1 vssd1 vccd1 vccd1 _3035_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold952 hold952/A vssd1 vssd1 vccd1 vccd1 _2892_/A sky130_fd_sc_hd__buf_1
Xhold963 _3715_/Q vssd1 vssd1 vccd1 vccd1 _3159_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold941 _3400_/Q vssd1 vssd1 vccd1 vccd1 hold941/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold985 _3328_/Q vssd1 vssd1 vccd1 vccd1 hold985/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold996 _3612_/Q vssd1 vssd1 vccd1 vccd1 hold996/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold974 _2063_/X vssd1 vssd1 vccd1 vccd1 _3629_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_66_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2204__A0 _2648_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2921_ _2876_/A _2918_/Y _2919_/X _2920_/Y _2944_/B vssd1 vssd1 vccd1 vccd1 _2921_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_0_15_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2852_ _2058_/A _2741_/A _2673_/B _2851_/Y _2850_/Y vssd1 vssd1 vccd1 vccd1 _2852_/X
+ sky130_fd_sc_hd__o41a_1
XANTENNA__1918__B _2022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2783_ _2797_/A hold569/X _2731_/X vssd1 vssd1 vccd1 vccd1 _2783_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_31_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1803_ _2085_/A _1803_/B vssd1 vssd1 vccd1 vccd1 _1803_/Y sky130_fd_sc_hd__nor2_1
X_1734_ _2006_/A _1734_/B vssd1 vssd1 vccd1 vccd1 _1734_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_13_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold215 _3593_/Q vssd1 vssd1 vccd1 vccd1 hold215/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold204 _2664_/X vssd1 vssd1 vccd1 vccd1 _3590_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold226 _2489_/X vssd1 vssd1 vccd1 vccd1 _3442_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold248 _2636_/X vssd1 vssd1 vccd1 vccd1 _3566_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold259 _3534_/Q vssd1 vssd1 vccd1 vccd1 hold259/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold237 _3588_/Q vssd1 vssd1 vccd1 vccd1 hold237/X sky130_fd_sc_hd__dlygate4sd3_1
X_1665_ _2669_/B _2741_/B _1673_/C vssd1 vssd1 vccd1 vccd1 _2846_/B sky130_fd_sc_hd__or3_2
X_3404_ _3725_/CLK _3404_/D vssd1 vssd1 vccd1 vccd1 _3404_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3335_ _3738_/CLK _3335_/D vssd1 vssd1 vccd1 vccd1 _3335_/Q sky130_fd_sc_hd__dfxtp_1
X_3266_ _3419_/CLK _3266_/D vssd1 vssd1 vccd1 vccd1 _3266_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2217_ _2659_/A0 hold555/X _2218_/S vssd1 vssd1 vccd1 vccd1 _2217_/X sky130_fd_sc_hd__mux2_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2765__A _2797_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2277__A3 _2652_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3197_ _3197_/A0 hold691/X _3198_/S vssd1 vssd1 vccd1 vccd1 _3197_/X sky130_fd_sc_hd__mux2_1
X_2148_ _3716_/Q _3715_/Q _3717_/Q vssd1 vssd1 vccd1 vccd1 _2149_/C sky130_fd_sc_hd__a21oi_1
X_2079_ _2669_/A _2079_/B vssd1 vssd1 vccd1 vccd1 _2080_/C sky130_fd_sc_hd__and2_1
XFILLER_0_72_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold760 _2981_/X vssd1 vssd1 vccd1 vccd1 _3656_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout93_A _2089_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold782 _2446_/X vssd1 vssd1 vccd1 vccd1 _3407_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold771 _3271_/Q vssd1 vssd1 vccd1 vccd1 hold771/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold793 _3649_/Q vssd1 vssd1 vccd1 vccd1 hold793/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2976__A1 _3594_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2728__A1 hold908/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3120_ _3120_/A _3120_/B vssd1 vssd1 vccd1 vccd1 _3120_/Y sky130_fd_sc_hd__nand2_1
X_3051_ _3053_/B _3048_/X _3050_/X vssd1 vssd1 vccd1 vccd1 _3051_/X sky130_fd_sc_hd__o21ba_1
X_2002_ _3549_/Q hold27/A _3573_/Q _3238_/Q _2289_/B _2289_/C vssd1 vssd1 vccd1 vccd1
+ _2002_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_26_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2904_ _2904_/A _2904_/B vssd1 vssd1 vccd1 vccd1 _2904_/X sky130_fd_sc_hd__or2_1
XFILLER_0_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2835_ _2871_/A _2863_/C vssd1 vssd1 vccd1 vccd1 _2835_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_60_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2766_ _2797_/A hold707/X _2731_/X vssd1 vssd1 vccd1 vccd1 _2766_/X sky130_fd_sc_hd__a21o_1
X_2697_ _2696_/A _2696_/B _2788_/A vssd1 vssd1 vccd1 vccd1 _2698_/C sky130_fd_sc_hd__a21boi_1
X_1717_ _3738_/Q _3216_/Q _3320_/Q _3338_/Q _1981_/S0 _1981_/S1 vssd1 vssd1 vccd1
+ vccd1 _1717_/X sky130_fd_sc_hd__mux4_1
XANTENNA__2479__B _2479_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1648_ _3626_/Q _3627_/Q _2669_/B vssd1 vssd1 vccd1 vccd1 _1713_/B sky130_fd_sc_hd__or3_2
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3318_ _3738_/CLK _3318_/D vssd1 vssd1 vccd1 vccd1 _3318_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3249_ _3436_/CLK _3249_/D vssd1 vssd1 vccd1 vccd1 _3249_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2495__A _2495_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2655__A0 _2655_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold590 _2990_/X vssd1 vssd1 vccd1 vccd1 _3665_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1792__S1 _2219_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1749__A _2085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2949__B2 _2885_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2620_ _2655_/A0 hold779/X _2625_/S vssd1 vssd1 vccd1 vccd1 _2620_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_88_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2551_ hold201/X _3194_/A0 _2555_/S vssd1 vssd1 vccd1 vccd1 _2551_/X sky130_fd_sc_hd__mux2_1
X_2482_ hold381/X _2353_/A _2487_/S vssd1 vssd1 vccd1 vccd1 _2482_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_2_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3103_ _3103_/A _3103_/B vssd1 vssd1 vccd1 vccd1 _3694_/D sky130_fd_sc_hd__nand2_1
XFILLER_0_37_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2637__A0 _2658_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_20_wb_clk_i_A clkbuf_3_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_3034_ _3086_/A _3034_/B _3035_/B vssd1 vssd1 vccd1 vccd1 _3034_/X sky130_fd_sc_hd__and3_1
XFILLER_0_37_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2254__S _2259_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout143_A _3346_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2818_ hold860/X _2080_/C _2871_/A _2082_/C vssd1 vssd1 vccd1 vccd1 _2825_/A sky130_fd_sc_hd__a211o_1
X_2749_ _2797_/A hold583/X _2731_/X vssd1 vssd1 vccd1 vccd1 _2749_/X sky130_fd_sc_hd__a21o_1
XANTENNA__2325__C1 _3108_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1774__S1 _1981_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2672__B _2868_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_24_wb_clk_i clkbuf_3_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3539_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_clkbuf_3_3__f_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1982_ hold13/A _3483_/Q _3465_/Q _3453_/Q _1760_/A _1760_/B vssd1 vssd1 vccd1 vccd1
+ _1982_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_23_98 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3721_ _3721_/CLK _3721_/D vssd1 vssd1 vccd1 vccd1 _3721_/Q sky130_fd_sc_hd__dfxtp_1
X_3652_ _3662_/CLK _3652_/D vssd1 vssd1 vccd1 vccd1 _3652_/Q sky130_fd_sc_hd__dfxtp_1
X_2603_ _2361_/A hold557/X _2604_/S vssd1 vssd1 vccd1 vccd1 _2603_/X sky130_fd_sc_hd__mux2_1
X_3583_ _3583_/CLK _3583_/D vssd1 vssd1 vccd1 vccd1 _3583_/Q sky130_fd_sc_hd__dfxtp_1
X_2534_ hold289/X _2363_/A _2534_/S vssd1 vssd1 vccd1 vccd1 _2534_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_70_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1942__A _2244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2465_ _2598_/A _2528_/B vssd1 vssd1 vccd1 vccd1 _2471_/S sky130_fd_sc_hd__nand2_4
X_2396_ _2643_/A1 hold475/X _2399_/S vssd1 vssd1 vccd1 vccd1 _2396_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2195__D _2480_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3017_ _3124_/A _3045_/D _3063_/A _3016_/X vssd1 vssd1 vccd1 vccd1 _3118_/B sky130_fd_sc_hd__o31a_1
XFILLER_0_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2010__A1 _2244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout130 _2185_/C vssd1 vssd1 vccd1 vccd1 _2245_/B sky130_fd_sc_hd__clkbuf_8
Xfanout141 _1988_/S vssd1 vssd1 vccd1 vccd1 _2244_/B sky130_fd_sc_hd__clkbuf_8
Xfanout152 _3172_/C1 vssd1 vssd1 vccd1 vccd1 _3103_/A sky130_fd_sc_hd__buf_4
XFILLER_0_69_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2250_ hold21/X _2651_/A0 _2252_/S vssd1 vssd1 vccd1 vccd1 hold22/A sky130_fd_sc_hd__mux2_1
XANTENNA__1738__S1 _2219_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2577__B _2647_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2181_ _2182_/A _2182_/B vssd1 vssd1 vccd1 vccd1 _2181_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_75_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1815__A1 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1965_ _2085_/C _1965_/B vssd1 vssd1 vccd1 vccd1 _1965_/Y sky130_fd_sc_hd__nand2_1
X_3704_ _3718_/CLK _3704_/D vssd1 vssd1 vccd1 vccd1 _3704_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1896_ _3541_/Q _3251_/Q _3517_/Q _3505_/Q _2000_/S0 _2219_/C vssd1 vssd1 vccd1 vccd1
+ _1896_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_43_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3635_ _3636_/CLK _3635_/D vssd1 vssd1 vccd1 vccd1 _3635_/Q sky130_fd_sc_hd__dfxtp_1
X_3566_ _3586_/CLK _3566_/D vssd1 vssd1 vccd1 vccd1 _3566_/Q sky130_fd_sc_hd__dfxtp_1
X_3497_ _3735_/CLK _3497_/D vssd1 vssd1 vccd1 vccd1 _3497_/Q sky130_fd_sc_hd__dfxtp_1
X_2517_ hold211/X _2643_/A1 _2520_/S vssd1 vssd1 vccd1 vccd1 _2517_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_59_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2448_ _3196_/A0 hold637/X _2450_/S vssd1 vssd1 vccd1 vccd1 _2448_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_52_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1729__S1 _2185_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2379_ _2570_/A _2407_/A vssd1 vssd1 vccd1 vccd1 _2385_/S sky130_fd_sc_hd__nand2_4
XANTENNA__2059__A1 _2076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2767__C1 _2859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1990__B1 _2428_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold8 hold8/A vssd1 vssd1 vccd1 vccd1 hold8/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1750_ _3260_/Q _3272_/Q _1937_/S vssd1 vssd1 vccd1 vccd1 _1751_/B sky130_fd_sc_hd__mux2_1
X_1681_ _1979_/A _1680_/X _2080_/B vssd1 vssd1 vccd1 vccd1 _1681_/X sky130_fd_sc_hd__a21o_1
Xhold408 _2976_/X vssd1 vssd1 vccd1 vccd1 _3651_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold419 _3572_/Q vssd1 vssd1 vccd1 vccd1 hold419/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3420_ _3496_/CLK _3420_/D vssd1 vssd1 vccd1 vccd1 _3420_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3351_ _3668_/CLK _3351_/D vssd1 vssd1 vccd1 vccd1 _3351_/Q sky130_fd_sc_hd__dfxtp_1
X_2302_ _2302_/A _3228_/Q _3227_/Q vssd1 vssd1 vccd1 vccd1 _2316_/B sky130_fd_sc_hd__or3b_1
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3282_ _3575_/CLK _3282_/D vssd1 vssd1 vccd1 vccd1 _3282_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2233_ _2475_/A1 hold499/X _2236_/S vssd1 vssd1 vccd1 vccd1 _2233_/X sky130_fd_sc_hd__mux2_1
X_2164_ _2164_/A _2164_/B _2164_/C _2164_/D vssd1 vssd1 vccd1 vccd1 _2164_/X sky130_fd_sc_hd__or4_1
X_2095_ hold893/X _2084_/A _2099_/B1 hold950/X vssd1 vssd1 vccd1 vccd1 _2359_/A sky130_fd_sc_hd__a22o_4
XFILLER_0_0_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1895__S0 _2000_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2997_ hold285/X _2997_/A1 _2999_/S vssd1 vssd1 vccd1 vccd1 _2997_/X sky130_fd_sc_hd__mux2_1
X_1948_ hold83/A _3584_/Q _3566_/Q _3554_/Q _2289_/B _2289_/C vssd1 vssd1 vccd1 vccd1
+ _1948_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_9_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1879_ _3431_/Q _3419_/Q _3407_/Q _3263_/Q _1981_/S0 _1981_/S1 vssd1 vssd1 vccd1
+ vccd1 _1879_/X sky130_fd_sc_hd__mux4_1
X_3618_ _3672_/CLK _3618_/D vssd1 vssd1 vccd1 vccd1 _3618_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold920 _3679_/Q vssd1 vssd1 vccd1 vccd1 _3030_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold931 _3034_/X vssd1 vssd1 vccd1 vccd1 _3680_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold953 _3135_/X vssd1 vssd1 vccd1 vccd1 hold953/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold964 _3159_/X vssd1 vssd1 vccd1 vccd1 hold964/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3174__C1 _3058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold942 _2438_/X vssd1 vssd1 vccd1 vccd1 _3400_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3549_ _3561_/CLK _3549_/D vssd1 vssd1 vccd1 vccd1 _3549_/Q sky130_fd_sc_hd__dfxtp_1
Xhold997 _2880_/X vssd1 vssd1 vccd1 vccd1 hold997/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold975 _3621_/Q vssd1 vssd1 vccd1 vccd1 _2924_/A sky130_fd_sc_hd__buf_1
Xhold986 _3682_/Q vssd1 vssd1 vccd1 vccd1 _3040_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__2452__A1 _2648_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2961__A _2961_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2680__B _2867_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2920_ _2924_/B _2924_/C _2935_/A vssd1 vssd1 vccd1 vccd1 _2920_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__2443__A1 _2653_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1877__S0 _1981_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2851_ _2851_/A _2851_/B vssd1 vssd1 vccd1 vccd1 _2851_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_31_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2782_ _2797_/A _2782_/B vssd1 vssd1 vccd1 vccd1 _2782_/Y sky130_fd_sc_hd__nor2_1
X_1802_ hold41/A hold65/A hold25/A _3223_/Q _2085_/B _2014_/A vssd1 vssd1 vccd1 vccd1
+ _1803_/B sky130_fd_sc_hd__mux4_1
X_1733_ hold11/A _3592_/Q _2244_/B vssd1 vssd1 vccd1 vccd1 _1734_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_31_98 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold216 _2667_/X vssd1 vssd1 vccd1 vccd1 _3593_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold205 _3431_/Q vssd1 vssd1 vccd1 vccd1 hold205/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold227 _3522_/Q vssd1 vssd1 vccd1 vccd1 hold227/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold238 _2662_/X vssd1 vssd1 vccd1 vccd1 _3588_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1664_ _2669_/B _2741_/B _1673_/C vssd1 vssd1 vccd1 vccd1 _3130_/A sky130_fd_sc_hd__nor3_4
XANTENNA__3156__C1 _3103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold249 _3637_/Q vssd1 vssd1 vccd1 vccd1 hold249/X sky130_fd_sc_hd__dlygate4sd3_1
X_3403_ _3725_/CLK _3403_/D vssd1 vssd1 vccd1 vccd1 _3403_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3334_ _3737_/CLK _3334_/D vssd1 vssd1 vccd1 vccd1 _3334_/Q sky130_fd_sc_hd__dfxtp_1
X_3265_ _3665_/CLK _3265_/D vssd1 vssd1 vccd1 vccd1 _3265_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2216_ _2658_/A0 hold657/X _2218_/S vssd1 vssd1 vccd1 vccd1 _2216_/X sky130_fd_sc_hd__mux2_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3196_ _3196_/A0 hold187/X _3198_/S vssd1 vssd1 vccd1 vccd1 _3196_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2257__S _2259_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2147_ _3706_/Q _2147_/B vssd1 vssd1 vccd1 vccd1 _2147_/Y sky130_fd_sc_hd__xnor2_1
X_2078_ _2669_/B _2742_/B vssd1 vssd1 vccd1 vccd1 _2079_/B sky130_fd_sc_hd__nor2_1
XANTENNA__2434__A1 _3203_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2198__A0 _2656_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_49_wb_clk_i clkbuf_3_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3672_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold761 _3396_/Q vssd1 vssd1 vccd1 vccd1 hold761/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold772 _2241_/X vssd1 vssd1 vccd1 vccd1 _3271_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold750 _2207_/X vssd1 vssd1 vccd1 vccd1 _3247_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout86_A _2650_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold794 _2974_/X vssd1 vssd1 vccd1 vccd1 _3649_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold783 _3322_/Q vssd1 vssd1 vccd1 vccd1 hold783/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2370__A0 _3197_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2675__B _2868_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2425__A1 _2658_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3050_ _3054_/A _3038_/Y _3048_/X _3053_/B _3108_/A vssd1 vssd1 vccd1 vccd1 _3050_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_leaf_10_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_2001_ _3283_/Q _3355_/Q _3367_/Q _3379_/Q _2289_/B _2289_/C vssd1 vssd1 vccd1 vccd1
+ _2001_/X sky130_fd_sc_hd__mux4_1
XANTENNA__2664__A1 _2357_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2903_ _2904_/A _2904_/B vssd1 vssd1 vccd1 vccd1 _2914_/C sky130_fd_sc_hd__and2_1
X_2834_ hold850/X _2824_/X _2832_/X _2833_/X _2859_/A vssd1 vssd1 vccd1 vccd1 _2834_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_5_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2765_ _2797_/A _2765_/B vssd1 vssd1 vccd1 vccd1 _2765_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_41_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3129__C1 _3055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2696_ _2696_/A _2696_/B vssd1 vssd1 vccd1 vccd1 _2700_/B sky130_fd_sc_hd__nand2_1
X_1716_ _1760_/A _1760_/B _2087_/B _1762_/B vssd1 vssd1 vccd1 vccd1 _1716_/X sky130_fd_sc_hd__or4_4
X_1647_ _2868_/B _1653_/C vssd1 vssd1 vccd1 vccd1 _1650_/A sky130_fd_sc_hd__nor2_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3317_ _3738_/CLK _3317_/D vssd1 vssd1 vccd1 vccd1 _3317_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3248_ _3436_/CLK _3248_/D vssd1 vssd1 vccd1 vccd1 _3248_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3179_ _3725_/Q _3181_/B vssd1 vssd1 vccd1 vccd1 _3179_/X sky130_fd_sc_hd__or2_1
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2678__A_N _2867_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2016__A _2085_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold580 _2628_/X vssd1 vssd1 vccd1 vccd1 _3559_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2343__A0 _2650_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold591 _3268_/Q vssd1 vssd1 vccd1 vccd1 hold591/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2646__A1 _2660_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2582__A0 _2659_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2550_ hold19/X _2655_/A0 _2555_/S vssd1 vssd1 vccd1 vccd1 hold20/A sky130_fd_sc_hd__mux2_1
X_2481_ _2612_/B _3199_/B vssd1 vssd1 vccd1 vccd1 _2487_/S sky130_fd_sc_hd__nor2_2
XFILLER_0_50_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2334__A0 _3195_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3102_ _3045_/B _2304_/X hold807/X vssd1 vssd1 vccd1 vccd1 _3102_/Y sky130_fd_sc_hd__o21ai_1
X_3033_ _3033_/A _3033_/B vssd1 vssd1 vccd1 vccd1 _3033_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_37_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout136_A _3346_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2817_ hold908/X _2871_/A _2816_/Y _2876_/B vssd1 vssd1 vccd1 vccd1 _2817_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_5_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2573__A0 _2357_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2748_ _3630_/Q _2746_/Y _2747_/X _2811_/A _2876_/B vssd1 vssd1 vccd1 vccd1 _2748_/X
+ sky130_fd_sc_hd__o221a_1
X_2679_ _3596_/Q _2867_/B vssd1 vssd1 vccd1 vccd1 _2759_/A sky130_fd_sc_hd__and2_1
XTAP_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2628__A1 _2656_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2564__A0 _2655_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2095__A2 _2084_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3044__A1 _3045_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1981_ _3385_/Q _3373_/Q _3361_/Q _3289_/Q _1981_/S0 _1981_/S1 vssd1 vssd1 vccd1
+ vccd1 _1981_/X sky130_fd_sc_hd__mux4_2
X_3720_ _3721_/CLK _3720_/D vssd1 vssd1 vccd1 vccd1 _3720_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3651_ _3662_/CLK _3651_/D vssd1 vssd1 vccd1 vccd1 _3651_/Q sky130_fd_sc_hd__dfxtp_1
X_2602_ _3203_/A1 hold533/X _2604_/S vssd1 vssd1 vccd1 vccd1 _2602_/X sky130_fd_sc_hd__mux2_1
X_3582_ _3735_/CLK _3582_/D vssd1 vssd1 vccd1 vccd1 _3582_/Q sky130_fd_sc_hd__dfxtp_1
X_2533_ hold273/X _2652_/A0 _2534_/S vssd1 vssd1 vccd1 vccd1 _2533_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_2_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2464_ _3198_/A0 hold615/X _2464_/S vssd1 vssd1 vccd1 vccd1 _2464_/X sky130_fd_sc_hd__mux2_1
X_2395_ _2656_/A0 hold639/X _2399_/S vssd1 vssd1 vccd1 vccd1 _2395_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3016_ _3124_/A _3015_/X _3013_/Y vssd1 vssd1 vccd1 vccd1 _3016_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_19_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2546__A0 _3203_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout120 _3349_/Q vssd1 vssd1 vccd1 vccd1 _2479_/B sky130_fd_sc_hd__clkbuf_4
Xfanout131 _1849_/S1 vssd1 vssd1 vccd1 vccd1 _2185_/C sky130_fd_sc_hd__clkbuf_8
Xfanout142 _1988_/S vssd1 vssd1 vccd1 vccd1 _1996_/S sky130_fd_sc_hd__clkbuf_4
Xfanout153 _3172_/C1 vssd1 vssd1 vccd1 vccd1 _3166_/C1 sky130_fd_sc_hd__buf_4
XFILLER_0_69_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1809__C1 _2479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2785__A0 _2868_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2180_ _3059_/B _3157_/B _2166_/X _2179_/X _3055_/A vssd1 vssd1 vccd1 vccd1 _2180_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_87_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1964_ _3231_/Q _3246_/Q _2085_/B vssd1 vssd1 vccd1 vccd1 _1965_/B sky130_fd_sc_hd__mux2_1
X_3703_ _3718_/CLK _3703_/D vssd1 vssd1 vccd1 vccd1 _3703_/Q sky130_fd_sc_hd__dfxtp_1
X_1895_ _3389_/Q _3583_/Q _3565_/Q _3553_/Q _2000_/S0 _2219_/C vssd1 vssd1 vccd1 vccd1
+ _1895_/X sky130_fd_sc_hd__mux4_1
X_3634_ _3668_/CLK _3634_/D vssd1 vssd1 vccd1 vccd1 _3634_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3565_ _3583_/CLK _3565_/D vssd1 vssd1 vccd1 vccd1 _3565_/Q sky130_fd_sc_hd__dfxtp_1
X_3496_ _3496_/CLK _3496_/D vssd1 vssd1 vccd1 vccd1 _3496_/Q sky130_fd_sc_hd__dfxtp_1
X_2516_ hold149/X _3194_/A0 _2520_/S vssd1 vssd1 vccd1 vccd1 _2516_/X sky130_fd_sc_hd__mux2_1
X_2447_ _2475_/A1 hold717/X _2450_/S vssd1 vssd1 vccd1 vccd1 _2447_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2378_ hold57/X _2653_/A0 _2378_/S vssd1 vssd1 vccd1 vccd1 hold58/A sky130_fd_sc_hd__mux2_1
XANTENNA__2059__A2 _2955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1990__A1 _1889_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold9 hold9/A vssd1 vssd1 vccd1 vccd1 hold9/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_71_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2860__C _3595_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold409 _3646_/Q vssd1 vssd1 vccd1 vccd1 hold409/X sky130_fd_sc_hd__dlygate4sd3_1
X_1680_ _1642_/X _1654_/B _2878_/B _1685_/B vssd1 vssd1 vccd1 vccd1 _1680_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_52_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3350_ _3668_/CLK _3350_/D vssd1 vssd1 vccd1 vccd1 _3350_/Q sky130_fd_sc_hd__dfxtp_1
X_2301_ _2301_/A _3225_/Q _2301_/C vssd1 vssd1 vccd1 vccd1 _3089_/A sky130_fd_sc_hd__and3_1
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3281_ _3583_/CLK _3281_/D vssd1 vssd1 vccd1 vccd1 _3281_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2232_ _3194_/A0 hold377/X _2236_/S vssd1 vssd1 vccd1 vccd1 _2232_/X sky130_fd_sc_hd__mux2_1
X_2163_ _2163_/A _2163_/B _2163_/C _2152_/X vssd1 vssd1 vccd1 vccd1 _2164_/D sky130_fd_sc_hd__or4b_1
X_2094_ hold91/X _2650_/A0 _2100_/S vssd1 vssd1 vccd1 vccd1 hold92/A sky130_fd_sc_hd__mux2_1
XANTENNA__1895__S1 _2219_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2749__B1 _2731_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2996_ hold385/X _2996_/A1 _2999_/S vssd1 vssd1 vccd1 vccd1 _2996_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_16_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1947_ _2185_/A _1944_/Y _1946_/Y _2428_/C _1942_/Y vssd1 vssd1 vccd1 vccd1 _1947_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_0_16_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1878_ _3493_/Q hold67/A _3463_/Q _3451_/Q _1981_/S0 _1981_/S1 vssd1 vssd1 vccd1
+ vccd1 _1878_/X sky130_fd_sc_hd__mux4_1
Xhold910 _3686_/Q vssd1 vssd1 vccd1 vccd1 _3053_/B sky130_fd_sc_hd__buf_2
X_3617_ _3718_/CLK _3617_/D vssd1 vssd1 vccd1 vccd1 _3617_/Q sky130_fd_sc_hd__dfxtp_1
Xhold921 _3029_/X vssd1 vssd1 vccd1 vccd1 _3031_/C sky130_fd_sc_hd__dlygate4sd3_1
X_3548_ _3575_/CLK _3548_/D vssd1 vssd1 vccd1 vccd1 _3548_/Q sky130_fd_sc_hd__dfxtp_1
Xhold943 _3601_/Q vssd1 vssd1 vccd1 vccd1 hold943/X sky130_fd_sc_hd__buf_1
Xhold932 hold932/A vssd1 vssd1 vccd1 vccd1 _2080_/A sky130_fd_sc_hd__clkbuf_2
Xhold954 _3136_/X vssd1 vssd1 vccd1 vccd1 _3704_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold998 _2882_/Y vssd1 vssd1 vccd1 vccd1 hold998/X sky130_fd_sc_hd__buf_1
Xhold987 _3041_/Y vssd1 vssd1 vccd1 vccd1 _3682_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold976 _3147_/X vssd1 vssd1 vccd1 vccd1 hold976/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold965 _3160_/X vssd1 vssd1 vccd1 vccd1 _3715_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3479_ _3732_/CLK _3479_/D vssd1 vssd1 vccd1 vccd1 _3479_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2912__B1 _2868_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2850_ _2809_/A _2711_/Y _2809_/B vssd1 vssd1 vccd1 vccd1 _2850_/Y sky130_fd_sc_hd__o21bai_1
XANTENNA__1877__S1 _1981_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1801_ _2244_/A _1797_/Y _1799_/X _1800_/Y vssd1 vssd1 vccd1 vccd1 _1801_/X sky130_fd_sc_hd__a31o_1
X_2781_ _2769_/Y _2863_/C _2811_/A vssd1 vssd1 vccd1 vccd1 _2782_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_25_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1732_ _2185_/C _1732_/B vssd1 vssd1 vccd1 vccd1 _1732_/Y sky130_fd_sc_hd__nand2_1
X_1663_ _3630_/Q _1663_/B vssd1 vssd1 vccd1 vccd1 _1673_/C sky130_fd_sc_hd__nand2_2
Xhold217 _3387_/Q vssd1 vssd1 vccd1 vccd1 hold217/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold206 _2474_/X vssd1 vssd1 vccd1 vccd1 _3431_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold228 _2585_/X vssd1 vssd1 vccd1 vccd1 _3522_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold239 _3669_/Q vssd1 vssd1 vccd1 vccd1 hold239/X sky130_fd_sc_hd__dlygate4sd3_1
X_3402_ _3725_/CLK _3402_/D vssd1 vssd1 vccd1 vccd1 _3402_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3333_ _3728_/CLK _3333_/D vssd1 vssd1 vccd1 vccd1 _3333_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3264_ _3496_/CLK _3264_/D vssd1 vssd1 vccd1 vccd1 _3264_/Q sky130_fd_sc_hd__dfxtp_1
X_2215_ _3195_/A0 hold257/X _2218_/S vssd1 vssd1 vccd1 vccd1 _2215_/X sky130_fd_sc_hd__mux2_1
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3195_ _3195_/A0 hold527/X _3198_/S vssd1 vssd1 vccd1 vccd1 _3195_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2146_ _2146_/A _2146_/B vssd1 vssd1 vccd1 vccd1 _2147_/B sky130_fd_sc_hd__or2_1
XFILLER_0_72_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2077_ _1663_/B _2073_/Y _2076_/X _2495_/A vssd1 vssd1 vccd1 vccd1 _2077_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_8_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2979_ hold569/X _2979_/A1 _2987_/S vssd1 vssd1 vccd1 vccd1 _2979_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_29_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold740 _2198_/X vssd1 vssd1 vccd1 vccd1 _3236_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold762 _2433_/X vssd1 vssd1 vccd1 vccd1 _3396_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold773 _3364_/Q vssd1 vssd1 vccd1 vccd1 hold773/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold751 _3358_/Q vssd1 vssd1 vccd1 vccd1 hold751/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold795 _3565_/Q vssd1 vssd1 vccd1 vccd1 hold795/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold784 _2340_/X vssd1 vssd1 vccd1 vccd1 _3322_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_18_wb_clk_i clkbuf_3_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3561_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_fanout79_A _3196_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2691__B _2867_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2830__C1 _2859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2189__A1 _2357_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2212__A _2570_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2000_ _3543_/Q _3253_/Q _3519_/Q _3507_/Q _2000_/S0 _2219_/C vssd1 vssd1 vccd1 vccd1
+ _2000_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_26_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2891__A2_N _2940_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1872__B1 _2701_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_6_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_2902_ hold571/X _2940_/B2 _2867_/C _1712_/A vssd1 vssd1 vccd1 vccd1 _2902_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_0_18_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2833_ _3597_/Q _1696_/Y _2940_/B2 hold327/X _2825_/Y vssd1 vssd1 vccd1 vccd1 _2833_/X
+ sky130_fd_sc_hd__a221o_1
X_2764_ _2752_/Y _2863_/B _2811_/A vssd1 vssd1 vccd1 vccd1 _2765_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_41_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1715_ _2085_/A _2228_/C vssd1 vssd1 vccd1 vccd1 _1762_/B sky130_fd_sc_hd__nand2_2
X_2695_ _2735_/A _2703_/C _2771_/A _2754_/A vssd1 vssd1 vccd1 vccd1 _2696_/B sky130_fd_sc_hd__o211ai_2
X_1646_ _1653_/C vssd1 vssd1 vccd1 vccd1 _1646_/Y sky130_fd_sc_hd__inv_2
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1961__A _2085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3316_ _3737_/CLK _3316_/D vssd1 vssd1 vccd1 vccd1 _3316_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3247_ _3322_/CLK _3247_/D vssd1 vssd1 vccd1 vccd1 _3247_/Q sky130_fd_sc_hd__dfxtp_1
X_3178_ _3712_/Q _3158_/Y hold867/X _3058_/A vssd1 vssd1 vccd1 vccd1 _3178_/X sky130_fd_sc_hd__o211a_1
X_2129_ _3726_/Q _3714_/Q vssd1 vssd1 vccd1 vccd1 _2129_/X sky130_fd_sc_hd__and2_1
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2040__B1 _2867_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold581 _3556_/Q vssd1 vssd1 vccd1 vccd1 hold581/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold570 _2979_/X vssd1 vssd1 vccd1 vccd1 _3654_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1777__S0 _2085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold592 _2238_/X vssd1 vssd1 vccd1 vccd1 _3268_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1854__B1 _2087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2480_ _2480_/A _3351_/Q _2480_/C _2428_/C vssd1 vssd1 vccd1 vccd1 _3199_/B sky130_fd_sc_hd__or4b_4
XFILLER_0_23_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3101_ _3103_/A _3101_/B vssd1 vssd1 vccd1 vccd1 _3693_/D sky130_fd_sc_hd__nand2_1
XFILLER_0_37_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3032_ _3033_/A _3033_/B vssd1 vssd1 vccd1 vccd1 _3034_/B sky130_fd_sc_hd__or2_1
X_2816_ _2871_/A _2816_/B vssd1 vssd1 vccd1 vccd1 _2816_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_26_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout129_A _1849_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2747_ _2867_/A hold918/X _2812_/S vssd1 vssd1 vccd1 vccd1 _2747_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_5_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2678_ _2867_/C _3597_/Q vssd1 vssd1 vccd1 vccd1 _2678_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_78_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1629_ _3681_/Q _3678_/Q _3677_/Q _3026_/B vssd1 vssd1 vccd1 vccd1 _1629_/Y sky130_fd_sc_hd__nor4_1
XFILLER_0_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1931__S0 _1760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2261__A0 _3193_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_33_wb_clk_i clkbuf_3_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3581_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_90_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1980_ _3737_/Q _3215_/Q _3319_/Q _3337_/Q _1981_/S0 _1981_/S1 vssd1 vssd1 vccd1
+ vccd1 _1980_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_55_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3650_ _3662_/CLK _3650_/D vssd1 vssd1 vccd1 vccd1 _3650_/Q sky130_fd_sc_hd__dfxtp_1
X_2601_ _3195_/A0 hold611/X _2604_/S vssd1 vssd1 vccd1 vccd1 _2601_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_70_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3581_ _3581_/CLK _3581_/D vssd1 vssd1 vccd1 vccd1 _3581_/Q sky130_fd_sc_hd__dfxtp_1
X_2532_ hold521/X _3203_/A1 _2534_/S vssd1 vssd1 vccd1 vccd1 _2532_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2555__A1 _3198_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2463_ _3197_/A0 hold799/X _2464_/S vssd1 vssd1 vccd1 vccd1 _2463_/X sky130_fd_sc_hd__mux2_1
X_2394_ _2655_/A0 hold773/X _2399_/S vssd1 vssd1 vccd1 vccd1 _2394_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_3_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3015_ _2310_/B _3007_/A _3014_/X vssd1 vssd1 vccd1 vccd1 _3015_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_3_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2491__A0 _2650_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2243__A0 _2653_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout110 _2006_/A vssd1 vssd1 vccd1 vccd1 _2085_/C sky130_fd_sc_hd__buf_4
XFILLER_0_10_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout121 _3349_/Q vssd1 vssd1 vccd1 vccd1 _2087_/A sky130_fd_sc_hd__clkbuf_8
Xfanout143 _3346_/Q vssd1 vssd1 vccd1 vccd1 _1988_/S sky130_fd_sc_hd__buf_4
Xfanout154 _3172_/C1 vssd1 vssd1 vccd1 vccd1 _3055_/A sky130_fd_sc_hd__buf_4
Xfanout132 hold1038/X vssd1 vssd1 vccd1 vccd1 _1849_/S1 sky130_fd_sc_hd__buf_4
XFILLER_0_69_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2234__A0 _3196_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2225__A0 _2652_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1963_ _2014_/A _1963_/B vssd1 vssd1 vccd1 vccd1 _1963_/Y sky130_fd_sc_hd__nand2_1
X_1894_ _1889_/A _1891_/Y _1893_/Y _2428_/C _1889_/Y vssd1 vssd1 vccd1 vccd1 _1894_/X
+ sky130_fd_sc_hd__a311o_1
X_3702_ _3702_/CLK _3702_/D vssd1 vssd1 vccd1 vccd1 _3702_/Q sky130_fd_sc_hd__dfxtp_1
X_3633_ _3668_/CLK _3633_/D vssd1 vssd1 vccd1 vccd1 _3633_/Q sky130_fd_sc_hd__dfxtp_1
X_3564_ _3587_/CLK _3564_/D vssd1 vssd1 vccd1 vccd1 _3564_/Q sky130_fd_sc_hd__dfxtp_1
X_2515_ hold255/X _2655_/A0 _2520_/S vssd1 vssd1 vccd1 vccd1 _2515_/X sky130_fd_sc_hd__mux2_1
X_3495_ _3496_/CLK hold14/X vssd1 vssd1 vccd1 vccd1 hold13/A sky130_fd_sc_hd__dfxtp_1
X_2446_ _3194_/A0 hold781/X _2450_/S vssd1 vssd1 vccd1 vccd1 _2446_/X sky130_fd_sc_hd__mux2_1
X_2377_ hold87/X _2652_/A0 _2378_/S vssd1 vssd1 vccd1 vccd1 hold88/A sky130_fd_sc_hd__mux2_1
XFILLER_0_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2464__A0 _3198_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2216__A0 _2658_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2519__A1 _3197_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2207__A0 _2651_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3280_ _3570_/CLK _3280_/D vssd1 vssd1 vccd1 vccd1 _3280_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2930__B2 _2885_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2300_ _2300_/A vssd1 vssd1 vccd1 vccd1 _2303_/A sky130_fd_sc_hd__inv_2
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2231_ _3193_/A0 hold517/X _2236_/S vssd1 vssd1 vccd1 vccd1 _2231_/X sky130_fd_sc_hd__mux2_1
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2162_ _3715_/Q _3703_/Q _2147_/Y _2149_/Y _2150_/X vssd1 vssd1 vccd1 vccd1 _2163_/C
+ sky130_fd_sc_hd__a2111o_1
X_2093_ hold923/X _2084_/A _2099_/B1 hold850/X vssd1 vssd1 vccd1 vccd1 _2093_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_45_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2749__A1 _2797_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2995_ hold805/X _3607_/Q _2999_/S vssd1 vssd1 vccd1 vccd1 _2995_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_16_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1946_ _2006_/A _1946_/B vssd1 vssd1 vccd1 vccd1 _1946_/Y sky130_fd_sc_hd__nand2_1
X_1877_ _3383_/Q _3371_/Q _3359_/Q _3287_/Q _1981_/S0 _1981_/S1 vssd1 vssd1 vccd1
+ vccd1 _1877_/X sky130_fd_sc_hd__mux4_1
Xhold911 _3051_/X vssd1 vssd1 vccd1 vccd1 _3686_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3616_ _3676_/CLK _3616_/D vssd1 vssd1 vccd1 vccd1 _3616_/Q sky130_fd_sc_hd__dfxtp_1
Xhold922 _3031_/X vssd1 vssd1 vccd1 vccd1 _3679_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold900 _3327_/Q vssd1 vssd1 vccd1 vccd1 hold900/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1972__A2 _2022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3547_ _3561_/CLK _3547_/D vssd1 vssd1 vccd1 vccd1 _3547_/Q sky130_fd_sc_hd__dfxtp_1
Xhold944 _2830_/X vssd1 vssd1 vccd1 vccd1 _3601_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold933 _1693_/X vssd1 vssd1 vccd1 vccd1 _3311_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold955 _3405_/Q vssd1 vssd1 vccd1 vccd1 hold955/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold988 _3312_/Q vssd1 vssd1 vccd1 vccd1 hold988/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2921__A1 _2876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold977 _3148_/X vssd1 vssd1 vccd1 vccd1 _3710_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold966 _3706_/Q vssd1 vssd1 vccd1 vccd1 hold966/X sky130_fd_sc_hd__dlygate4sd3_1
X_3478_ _3732_/CLK _3478_/D vssd1 vssd1 vccd1 vccd1 _3478_/Q sky130_fd_sc_hd__dfxtp_1
Xhold999 _2911_/X vssd1 vssd1 vccd1 vccd1 _3618_/D sky130_fd_sc_hd__dlygate4sd3_1
X_2429_ _3185_/B vssd1 vssd1 vccd1 vccd1 _2528_/B sky130_fd_sc_hd__inv_2
XANTENNA__2988__A1 _1760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2437__B1 _2598_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2912__B2 _1712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1800_ _2244_/A _1795_/X _2087_/A vssd1 vssd1 vccd1 vccd1 _1800_/Y sky130_fd_sc_hd__o21ai_1
X_2780_ _2718_/B _2774_/Y _2790_/A _2777_/Y _2779_/X vssd1 vssd1 vccd1 vccd1 _2863_/C
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_31_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2600__A0 _3201_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1731_ _3532_/Q _3398_/Q _1996_/S vssd1 vssd1 vccd1 vccd1 _1732_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_13_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold207 _3233_/Q vssd1 vssd1 vccd1 vccd1 hold207/X sky130_fd_sc_hd__dlygate4sd3_1
X_1662_ _1678_/A _1662_/B vssd1 vssd1 vccd1 vccd1 _1698_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_53_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3401_ _3725_/CLK _3401_/D vssd1 vssd1 vccd1 vccd1 _3401_/Q sky130_fd_sc_hd__dfxtp_1
Xhold218 _2420_/X vssd1 vssd1 vccd1 vccd1 _3387_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold229 _3735_/Q vssd1 vssd1 vccd1 vccd1 hold229/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2364__C1 _3172_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3332_ _3447_/CLK _3332_/D vssd1 vssd1 vccd1 vccd1 _3332_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1723__S _1937_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3263_ _3419_/CLK _3263_/D vssd1 vssd1 vccd1 vccd1 _3263_/Q sky130_fd_sc_hd__dfxtp_1
X_2214_ _2656_/A0 hold553/X _2218_/S vssd1 vssd1 vccd1 vccd1 _2214_/X sky130_fd_sc_hd__mux2_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3194_ _3194_/A0 hold229/X _3198_/S vssd1 vssd1 vccd1 vccd1 _3194_/X sky130_fd_sc_hd__mux2_1
X_2145_ _3718_/Q _2149_/B vssd1 vssd1 vccd1 vccd1 _2146_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_56_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2076_ _2076_/A _2497_/A _2076_/C vssd1 vssd1 vccd1 vccd1 _2076_/X sky130_fd_sc_hd__or3_1
XANTENNA__1678__B _1922_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2978_ hold707/X _3596_/Q _2987_/S vssd1 vssd1 vccd1 vccd1 _2978_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_71_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1929_ _3736_/Q _3214_/Q _3318_/Q _3336_/Q _1981_/S0 _1981_/S1 vssd1 vssd1 vccd1
+ vccd1 _1929_/X sky130_fd_sc_hd__mux4_1
XANTENNA__1694__A _2876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold730 _2547_/X vssd1 vssd1 vccd1 vccd1 _3490_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold741 _3394_/Q vssd1 vssd1 vccd1 vccd1 hold741/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold752 _2387_/X vssd1 vssd1 vccd1 vccd1 _3358_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold763 _3216_/Q vssd1 vssd1 vccd1 vccd1 hold763/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold796 _2635_/X vssd1 vssd1 vccd1 vccd1 _3565_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold774 _2394_/X vssd1 vssd1 vccd1 vccd1 _3364_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_394 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold785 _3695_/Q vssd1 vssd1 vccd1 vccd1 hold785/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2658__A0 _2658_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1795__S1 _1849_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2649__A0 _2355_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold90 hold90/A vssd1 vssd1 vccd1 vccd1 hold90/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2901_ _3137_/A _2944_/B _2900_/Y _3103_/A vssd1 vssd1 vccd1 vccd1 _2901_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_42_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2832_ _3596_/Q _2871_/A _2831_/Y _2876_/B vssd1 vssd1 vccd1 vccd1 _2832_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_45_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2763_ _2718_/B _2757_/X _2775_/A _2760_/X _2762_/X vssd1 vssd1 vccd1 vccd1 _2863_/B
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_41_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1714_ _2228_/A _2195_/B vssd1 vssd1 vccd1 vccd1 _2087_/B sky130_fd_sc_hd__nand2_4
X_2694_ _3596_/Q _2689_/B _2771_/A _2678_/X vssd1 vssd1 vccd1 vccd1 _2696_/A sky130_fd_sc_hd__a31oi_2
X_1645_ _2669_/A _1663_/B vssd1 vssd1 vccd1 vccd1 _1653_/C sky130_fd_sc_hd__or2_2
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3315_ _3692_/CLK _3315_/D vssd1 vssd1 vccd1 vccd1 _3315_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3246_ _3322_/CLK _3246_/D vssd1 vssd1 vccd1 vccd1 _3246_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3177_ _3177_/A _3181_/B vssd1 vssd1 vccd1 vccd1 _3177_/X sky130_fd_sc_hd__or2_1
XFILLER_0_83_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1863__A1 _2479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2128_ _3726_/Q _3714_/Q vssd1 vssd1 vccd1 vccd1 _2128_/Y sky130_fd_sc_hd__nor2_1
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2059_ _2076_/A _2955_/A _2076_/C _2058_/X _1979_/A vssd1 vssd1 vccd1 vccd1 _3627_/D
+ sky130_fd_sc_hd__o311a_1
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2812__A0 _2868_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout91_A _2091_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold560 _2243_/X vssd1 vssd1 vccd1 vccd1 _3273_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold571 _3640_/Q vssd1 vssd1 vccd1 vccd1 hold571/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold593 _3744_/Q vssd1 vssd1 vccd1 vccd1 hold593/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold582 _2624_/X vssd1 vssd1 vccd1 vccd1 _3556_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1777__S1 _2228_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1854__A1 _2244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3100_ _3099_/X _1704_/B _3100_/S vssd1 vssd1 vccd1 vccd1 _3100_/X sky130_fd_sc_hd__mux2_1
X_3031_ _3033_/B _3086_/A _3031_/C vssd1 vssd1 vccd1 vccd1 _3031_/X sky130_fd_sc_hd__and3b_1
XANTENNA__2098__A1 _3197_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_3_wb_clk_i clkbuf_leaf_5_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3387_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_73_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2815_ hold934/X _2730_/Y _2813_/X _2814_/X _2859_/A vssd1 vssd1 vccd1 vccd1 _2815_/X
+ sky130_fd_sc_hd__o221a_1
X_2746_ _2863_/A vssd1 vssd1 vccd1 vccd1 _2746_/Y sky130_fd_sc_hd__inv_2
X_2677_ _2675_/X _2677_/B vssd1 vssd1 vccd1 vccd1 _2788_/A sky130_fd_sc_hd__nand2b_2
XFILLER_0_41_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1781__B1 _2289_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1628_ _3033_/A _3030_/A vssd1 vssd1 vccd1 vccd1 _3026_/B sky130_fd_sc_hd__or2_1
XANTENNA__1911__S _2085_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2089__A1 hold908/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3229_ _3322_/CLK _3229_/D vssd1 vssd1 vccd1 vccd1 _3229_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1836__A1 _1889_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1931__S1 _1760_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold390 _2966_/X vssd1 vssd1 vccd1 vccd1 _3641_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_74_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2252__A1 _2653_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2600_ _3201_/A1 hold395/X _2604_/S vssd1 vssd1 vccd1 vccd1 _2600_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_82_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3580_ _3581_/CLK _3580_/D vssd1 vssd1 vccd1 vccd1 _3580_/Q sky130_fd_sc_hd__dfxtp_1
X_2531_ hold245/X _2357_/A _2534_/S vssd1 vssd1 vccd1 vccd1 _2531_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_11_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2462_ _3196_/A0 hold737/X _2464_/S vssd1 vssd1 vccd1 vccd1 _2462_/X sky130_fd_sc_hd__mux2_1
X_2393_ _2407_/A _2647_/A vssd1 vssd1 vccd1 vccd1 _2399_/S sky130_fd_sc_hd__nand2_4
XANTENNA__2400__B _3199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3014_ _3014_/A _3684_/Q _3045_/D vssd1 vssd1 vccd1 vccd1 _3014_/X sky130_fd_sc_hd__or3_1
XANTENNA__1818__B2 _2854_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout141_A _1988_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2729_ _2811_/A _2728_/X _2726_/Y _2876_/B vssd1 vssd1 vccd1 vccd1 _2729_/X sky130_fd_sc_hd__o211a_1
XANTENNA__1754__B1 _2228_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout111 _1625_/Y vssd1 vssd1 vccd1 vccd1 _2006_/A sky130_fd_sc_hd__buf_4
Xfanout122 _3349_/Q vssd1 vssd1 vccd1 vccd1 _2428_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout144 hold988/X vssd1 vssd1 vccd1 vccd1 _2797_/A sky130_fd_sc_hd__buf_4
Xfanout155 _3172_/C1 vssd1 vssd1 vccd1 vccd1 _3086_/A sky130_fd_sc_hd__clkbuf_2
Xfanout133 _1760_/A vssd1 vssd1 vccd1 vccd1 _1981_/S0 sky130_fd_sc_hd__buf_8
XANTENNA__1809__A1 _2087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2936__A1_N _2885_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2482__A1 _2353_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2038__A _2074_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1745__B1 _2085_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2220__B _2647_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2473__A1 _3193_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1962_ _3258_/Q _3270_/Q _2085_/B vssd1 vssd1 vccd1 vccd1 _1963_/B sky130_fd_sc_hd__mux2_1
X_1893_ _2006_/A _1893_/B vssd1 vssd1 vccd1 vccd1 _1893_/Y sky130_fd_sc_hd__nand2_1
X_3701_ _3702_/CLK _3701_/D vssd1 vssd1 vccd1 vccd1 _3701_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_50_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3632_ _3670_/CLK _3632_/D vssd1 vssd1 vccd1 vccd1 _3632_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_3_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3563_ _3575_/CLK _3563_/D vssd1 vssd1 vccd1 vccd1 _3563_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3494_ _3558_/CLK _3494_/D vssd1 vssd1 vccd1 vccd1 _3494_/Q sky130_fd_sc_hd__dfxtp_1
X_2514_ _2640_/A _2549_/A vssd1 vssd1 vccd1 vccd1 _2520_/S sky130_fd_sc_hd__nor2_2
X_2445_ _3193_/A0 hold575/X _2450_/S vssd1 vssd1 vccd1 vccd1 _2445_/X sky130_fd_sc_hd__mux2_1
X_2376_ hold115/X _2651_/A0 _2378_/S vssd1 vssd1 vccd1 vccd1 _2376_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_91_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1727__B1 _2087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2455__A1 _3203_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1966__B1 _2087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3168__C1 _3172_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2391__A0 _3197_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2230_ _2500_/B _2598_/A vssd1 vssd1 vccd1 vccd1 _2236_/S sky130_fd_sc_hd__nand2_2
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2885__B _2885_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2161_ _2161_/A _2161_/B vssd1 vssd1 vccd1 vccd1 _2164_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_88_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2092_ hold165/X _2091_/X _2100_/S vssd1 vssd1 vccd1 vccd1 _2092_/X sky130_fd_sc_hd__mux2_1
X_2994_ hold239/X _2994_/A1 _2999_/S vssd1 vssd1 vccd1 vccd1 _2994_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_56_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1945_ _3458_/Q _3590_/Q _2244_/B vssd1 vssd1 vccd1 vccd1 _1946_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_28_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1957__B1 _2006_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1876_ _3735_/Q _3213_/Q _3317_/Q _3335_/Q _1760_/A _1981_/S1 vssd1 vssd1 vccd1 vccd1
+ _1876_/X sky130_fd_sc_hd__mux4_1
Xhold912 _3688_/Q vssd1 vssd1 vccd1 vccd1 _2305_/A sky130_fd_sc_hd__clkbuf_2
X_3615_ _3676_/CLK _3615_/D vssd1 vssd1 vccd1 vccd1 _3615_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold901 _2349_/X vssd1 vssd1 vccd1 vccd1 _2350_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2382__A0 _3195_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3546_ _3558_/CLK hold48/X vssd1 vssd1 vccd1 vccd1 hold47/A sky130_fd_sc_hd__dfxtp_1
Xhold934 _3599_/Q vssd1 vssd1 vccd1 vccd1 hold934/X sky130_fd_sc_hd__buf_1
Xhold945 _3684_/Q vssd1 vssd1 vccd1 vccd1 _3045_/A sky130_fd_sc_hd__clkbuf_2
Xhold923 _3596_/Q vssd1 vssd1 vccd1 vccd1 hold923/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold956 _3331_/Q vssd1 vssd1 vccd1 vccd1 hold956/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold978 _3600_/Q vssd1 vssd1 vccd1 vccd1 hold978/X sky130_fd_sc_hd__buf_1
Xhold989 _2893_/Y vssd1 vssd1 vccd1 vccd1 hold989/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold967 _3140_/X vssd1 vssd1 vccd1 vccd1 _3706_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3477_ _3732_/CLK _3477_/D vssd1 vssd1 vccd1 vccd1 _3477_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2428_ _2480_/A _3351_/Q _2428_/C _2480_/C vssd1 vssd1 vccd1 vccd1 _3185_/B sky130_fd_sc_hd__or4_4
X_2359_ _2359_/A _2363_/B vssd1 vssd1 vccd1 vccd1 _2359_/X sky130_fd_sc_hd__or2_1
XANTENNA__2437__A1 _3108_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2912__A2 _2940_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1939__B1 _2428_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1730_ _1889_/A _1730_/B vssd1 vssd1 vccd1 vccd1 _1730_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__2061__C1 _1979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold208 _2191_/X vssd1 vssd1 vccd1 vccd1 _3233_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1661_ _3630_/Q _1663_/B _2669_/C _2742_/B vssd1 vssd1 vccd1 vccd1 _1662_/B sky130_fd_sc_hd__or4_1
X_3400_ _3725_/CLK _3400_/D vssd1 vssd1 vccd1 vccd1 _3400_/Q sky130_fd_sc_hd__dfxtp_1
Xhold219 _3496_/Q vssd1 vssd1 vccd1 vccd1 hold219/X sky130_fd_sc_hd__dlygate4sd3_1
X_3331_ _3447_/CLK _3331_/D vssd1 vssd1 vccd1 vccd1 _3331_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2116__A0 _2650_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3262_ _3665_/CLK _3262_/D vssd1 vssd1 vccd1 vccd1 _3262_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2667__A1 _2363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2213_ _2655_/A0 hold459/X _2218_/S vssd1 vssd1 vccd1 vccd1 _2213_/X sky130_fd_sc_hd__mux2_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3193_ _3193_/A0 hold541/X _3198_/S vssd1 vssd1 vccd1 vccd1 _3193_/X sky130_fd_sc_hd__mux2_1
X_2144_ _3707_/Q _2144_/B vssd1 vssd1 vccd1 vccd1 _2163_/B sky130_fd_sc_hd__xnor2_1
X_2075_ _2034_/B _2073_/Y _2074_/X _2495_/A vssd1 vssd1 vccd1 vccd1 _2075_/X sky130_fd_sc_hd__o211a_1
XANTENNA__2419__A1 _3197_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_334 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2977_ hold583/X _3595_/Q _2987_/S vssd1 vssd1 vccd1 vccd1 _2977_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1975__A _2867_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1928_ _2076_/A _2028_/S _1927_/Y _1979_/A vssd1 vssd1 vccd1 vccd1 _3607_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_71_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1859_ _2014_/A _1859_/B vssd1 vssd1 vccd1 vccd1 _1859_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_12_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold720 _2450_/X vssd1 vssd1 vccd1 vccd1 _3411_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold731 _3554_/Q vssd1 vssd1 vccd1 vccd1 hold731/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold742 _2431_/X vssd1 vssd1 vccd1 vccd1 _3394_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold753 _3359_/Q vssd1 vssd1 vccd1 vccd1 hold753/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold764 _2110_/X vssd1 vssd1 vccd1 vccd1 _3216_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold797 _3525_/Q vssd1 vssd1 vccd1 vccd1 hold797/X sky130_fd_sc_hd__dlygate4sd3_1
X_3529_ _3733_/CLK _3529_/D vssd1 vssd1 vccd1 vccd1 _3529_/Q sky130_fd_sc_hd__dfxtp_1
Xhold775 _3249_/Q vssd1 vssd1 vccd1 vccd1 hold775/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold786 _3107_/Y vssd1 vssd1 vccd1 vccd1 _3108_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_67_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2046__A _2046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_27_wb_clk_i clkbuf_3_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3745_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__1885__A _2245_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2043__C1 _1979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold80 hold80/A vssd1 vssd1 vccd1 vccd1 hold80/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold91 hold91/A vssd1 vssd1 vccd1 vccd1 hold91/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1872__A2 _2731_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2900_ _2944_/B _2900_/B vssd1 vssd1 vccd1 vccd1 _2900_/Y sky130_fd_sc_hd__nand2_1
X_2831_ _2871_/A _2863_/B vssd1 vssd1 vccd1 vccd1 _2831_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_26_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2585__A0 _2655_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2762_ _2762_/A _2809_/B _2762_/C vssd1 vssd1 vccd1 vccd1 _2762_/X sky130_fd_sc_hd__or3_1
XFILLER_0_84_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1713_ _2669_/A _1713_/B _2082_/C vssd1 vssd1 vccd1 vccd1 _1713_/X sky130_fd_sc_hd__or3_4
XFILLER_0_13_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2693_ _2771_/A vssd1 vssd1 vccd1 vccd1 _2705_/C sky130_fd_sc_hd__inv_2
XANTENNA__2337__A0 _3198_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1644_ _2712_/A _3627_/Q _2669_/B vssd1 vssd1 vccd1 vccd1 _2868_/B sky130_fd_sc_hd__or3_2
XANTENNA__2888__A1 _2876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3314_ _3692_/CLK _3314_/D vssd1 vssd1 vccd1 vccd1 _3314_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3245_ _3322_/CLK _3245_/D vssd1 vssd1 vccd1 vccd1 _3245_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3176_ _3711_/Q _3158_/Y hold886/X _3058_/A vssd1 vssd1 vccd1 vccd1 _3176_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_13_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2127_ _3725_/Q _2135_/B vssd1 vssd1 vccd1 vccd1 _2132_/C sky130_fd_sc_hd__nand2_1
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2058_ _2058_/A _2062_/B vssd1 vssd1 vccd1 vccd1 _2058_/X sky130_fd_sc_hd__or2_1
XFILLER_0_49_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2273__C1 _3058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1909__S _2085_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2576__A0 _2363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2040__A2 _2731_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold561 _3557_/Q vssd1 vssd1 vccd1 vccd1 hold561/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold572 _2965_/X vssd1 vssd1 vccd1 vccd1 _3640_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold550 _2449_/X vssd1 vssd1 vccd1 vccd1 _3410_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold594 _3204_/X vssd1 vssd1 vccd1 vccd1 _3744_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold583 _3652_/Q vssd1 vssd1 vccd1 vccd1 hold583/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout84_A _2475_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2567__A0 _2658_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3030_ _3030_/A _3678_/Q _3677_/Q _3080_/A vssd1 vssd1 vccd1 vccd1 _3033_/B sky130_fd_sc_hd__and4_1
XANTENNA_clkbuf_3_0__f_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2814_ _2797_/A hold759/X _2731_/X vssd1 vssd1 vccd1 vccd1 _2814_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_5_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2745_ _2738_/Y _2739_/X _2743_/X _2744_/X vssd1 vssd1 vccd1 vccd1 _2863_/A sky130_fd_sc_hd__o211a_1
X_2676_ _3598_/Q _2868_/C vssd1 vssd1 vccd1 vccd1 _2677_/B sky130_fd_sc_hd__or2_1
XFILLER_0_41_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1781__A1 _2245_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1627_ _1627_/A vssd1 vssd1 vccd1 vccd1 _1627_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2730__B1 _2854_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3228_ _3727_/CLK _3228_/D vssd1 vssd1 vccd1 vccd1 _3228_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2089__A2 _2084_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3159_ _3159_/A _3181_/B vssd1 vssd1 vccd1 vccd1 _3159_/X sky130_fd_sc_hd__or2_1
XFILLER_0_49_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold380 _2118_/X vssd1 vssd1 vccd1 vccd1 _3222_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold391 _3206_/Q vssd1 vssd1 vccd1 vccd1 hold391/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1080 _3617_/Q vssd1 vssd1 vccd1 vccd1 _2965_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_42_wb_clk_i clkbuf_3_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3727_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__3201__A1 _3201_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2530_ hold97/X _3201_/A1 _2534_/S vssd1 vssd1 vccd1 vccd1 hold98/A sky130_fd_sc_hd__mux2_1
XFILLER_0_23_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2461_ _2475_/A1 hold693/X _2464_/S vssd1 vssd1 vccd1 vccd1 _2461_/X sky130_fd_sc_hd__mux2_1
X_2392_ _3198_/A0 hold293/X _2392_/S vssd1 vssd1 vccd1 vccd1 _2392_/X sky130_fd_sc_hd__mux2_1
X_3013_ _3010_/B _3012_/X _3124_/A vssd1 vssd1 vccd1 vccd1 _3013_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2728_ _2701_/B hold908/X _2812_/S vssd1 vssd1 vccd1 vccd1 _2728_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1754__A1 _2289_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2659_ _2659_/A0 hold393/X _2660_/S vssd1 vssd1 vccd1 vccd1 _2659_/X sky130_fd_sc_hd__mux2_1
Xfanout112 _2244_/A vssd1 vssd1 vccd1 vccd1 _1889_/A sky130_fd_sc_hd__buf_4
Xfanout156 _3172_/C1 vssd1 vssd1 vccd1 vccd1 _3058_/A sky130_fd_sc_hd__buf_4
Xfanout145 hold988/X vssd1 vssd1 vccd1 vccd1 _2819_/A sky130_fd_sc_hd__buf_2
Xfanout134 hold1062/X vssd1 vssd1 vccd1 vccd1 _1760_/A sky130_fd_sc_hd__clkbuf_8
Xfanout123 _2289_/A vssd1 vssd1 vccd1 vccd1 _2085_/A sky130_fd_sc_hd__buf_6
XFILLER_0_69_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1893__A _2006_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3195__A0 _3195_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1745__A1 _3773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3700_ _3702_/CLK _3700_/D vssd1 vssd1 vccd1 vccd1 _3700_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1961_ _2085_/A _1961_/B vssd1 vssd1 vccd1 vccd1 _1961_/Y sky130_fd_sc_hd__nor2_1
X_1892_ _3457_/Q _3589_/Q _1996_/S vssd1 vssd1 vccd1 vccd1 _1893_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_50_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3631_ _3637_/CLK _3631_/D vssd1 vssd1 vccd1 vccd1 _3631_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3562_ _3585_/CLK _3562_/D vssd1 vssd1 vccd1 vccd1 _3562_/Q sky130_fd_sc_hd__dfxtp_1
X_2513_ hold283/X _2363_/A _2513_/S vssd1 vssd1 vccd1 vccd1 _2513_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_3_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3493_ _3735_/CLK _3493_/D vssd1 vssd1 vccd1 vccd1 _3493_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2444_ _2647_/A _2500_/B vssd1 vssd1 vccd1 vccd1 _2450_/S sky130_fd_sc_hd__nand2_2
XFILLER_0_59_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2375_ hold133/X _2650_/A0 _2378_/S vssd1 vssd1 vccd1 vccd1 _2375_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1742__S _2244_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1727__A1 _1889_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1966__A1 _2085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2160_ hold992/X _3096_/B _2159_/X _3157_/B vssd1 vssd1 vccd1 vccd1 _2160_/X sky130_fd_sc_hd__o31a_1
X_2091_ hold918/X _2084_/A _2099_/B1 hold943/X vssd1 vssd1 vccd1 vccd1 _2091_/X sky130_fd_sc_hd__a22o_4
XFILLER_0_45_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2685__B1_N _3594_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2993_ hold473/X _2195_/B _2999_/S vssd1 vssd1 vccd1 vccd1 _2993_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_90_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1944_ _2185_/C _1944_/B vssd1 vssd1 vccd1 vccd1 _1944_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_71_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1957__A1 _3771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1875_ _1979_/A _1875_/B vssd1 vssd1 vccd1 vccd1 _3606_/D sky130_fd_sc_hd__and2_1
XFILLER_0_9_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3614_ _3672_/CLK _3614_/D vssd1 vssd1 vccd1 vccd1 _3614_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold913 _3057_/Y vssd1 vssd1 vccd1 vccd1 _3688_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold902 _3631_/Q vssd1 vssd1 vccd1 vccd1 _1663_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_0_24_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3545_ _3545_/CLK _3545_/D vssd1 vssd1 vccd1 vccd1 _3545_/Q sky130_fd_sc_hd__dfxtp_1
Xhold935 _2815_/X vssd1 vssd1 vccd1 vccd1 _3599_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold946 _3044_/Y vssd1 vssd1 vccd1 vccd1 hold946/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold924 _2767_/X vssd1 vssd1 vccd1 vccd1 _3596_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3476_ _3732_/CLK _3476_/D vssd1 vssd1 vccd1 vccd1 _3476_/Q sky130_fd_sc_hd__dfxtp_1
Xhold979 _2827_/X vssd1 vssd1 vccd1 vccd1 _3600_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold957 _3705_/Q vssd1 vssd1 vccd1 vccd1 hold957/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold968 _3401_/Q vssd1 vssd1 vccd1 vccd1 hold968/X sky130_fd_sc_hd__dlygate4sd3_1
X_2427_ hold157/X _2660_/A0 _2427_/S vssd1 vssd1 vccd1 vccd1 _2427_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_86_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2358_ hold981/X _2351_/Y _2357_/X _3058_/A vssd1 vssd1 vccd1 vccd1 _3330_/D sky130_fd_sc_hd__o211a_1
X_2289_ _2289_/A _2289_/B _2289_/C _2480_/C vssd1 vssd1 vccd1 vccd1 _2612_/B sky130_fd_sc_hd__or4_4
XANTENNA__2437__A2 _2084_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1740__S0 _2289_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2842__C1 _2859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2373__A1 _2648_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2507__A _2612_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1939__A1 _1889_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1660_ _3626_/Q _3627_/Q vssd1 vssd1 vccd1 vccd1 _2742_/B sky130_fd_sc_hd__nand2_2
Xhold209 _3562_/Q vssd1 vssd1 vccd1 vccd1 hold209/X sky130_fd_sc_hd__dlygate4sd3_1
X_3330_ _3447_/CLK _3330_/D vssd1 vssd1 vccd1 vccd1 _3330_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3261_ _3743_/CLK _3261_/D vssd1 vssd1 vccd1 vccd1 _3261_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2212_ _2570_/A _2654_/A vssd1 vssd1 vccd1 vccd1 _2218_/S sky130_fd_sc_hd__nand2_4
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3192_ _3192_/A _3192_/B vssd1 vssd1 vccd1 vccd1 _3198_/S sky130_fd_sc_hd__or2_4
XFILLER_0_56_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2143_ _3719_/Q _2146_/A vssd1 vssd1 vccd1 vccd1 _2144_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2074_ _2074_/A _2497_/A _2076_/C vssd1 vssd1 vccd1 vccd1 _2074_/X sky130_fd_sc_hd__or3_1
XANTENNA__1722__S0 _1937_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2976_ hold407/X _3594_/Q _2987_/S vssd1 vssd1 vccd1 vccd1 _2976_/X sky130_fd_sc_hd__mux2_1
X_1927_ _2028_/S _1927_/B vssd1 vssd1 vccd1 vccd1 _1927_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_16_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1858_ _3256_/Q _3268_/Q _2085_/B vssd1 vssd1 vccd1 vccd1 _1859_/B sky130_fd_sc_hd__mux2_1
Xhold710 _2411_/X vssd1 vssd1 vccd1 vccd1 _3379_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold721 _3375_/Q vssd1 vssd1 vccd1 vccd1 hold721/X sky130_fd_sc_hd__dlygate4sd3_1
X_1789_ _2245_/B _1786_/X _1788_/X vssd1 vssd1 vccd1 vccd1 _1789_/Y sky130_fd_sc_hd__a21oi_1
Xhold732 _2622_/X vssd1 vssd1 vccd1 vccd1 _3554_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold754 _2388_/X vssd1 vssd1 vccd1 vccd1 _3359_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold743 _3321_/Q vssd1 vssd1 vccd1 vccd1 hold743/X sky130_fd_sc_hd__dlygate4sd3_1
X_3528_ _3728_/CLK hold94/X vssd1 vssd1 vccd1 vccd1 hold93/A sky130_fd_sc_hd__dfxtp_1
Xhold776 _2209_/X vssd1 vssd1 vccd1 vccd1 _3249_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold787 _3244_/Q vssd1 vssd1 vccd1 vccd1 hold787/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold765 _3246_/Q vssd1 vssd1 vccd1 vccd1 hold765/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold798 _2588_/X vssd1 vssd1 vccd1 vccd1 _3525_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3459_ _3745_/CLK _3459_/D vssd1 vssd1 vccd1 vccd1 _3459_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2815__C1 _2859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2594__A1 _2650_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold81 hold81/A vssd1 vssd1 vccd1 vccd1 hold81/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1952__S0 _2289_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold70 hold70/A vssd1 vssd1 vccd1 vccd1 hold70/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_47 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold92 hold92/A vssd1 vssd1 vccd1 vccd1 hold92/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_85_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2830_ hold943/X _2824_/X _2828_/X _2829_/X _2859_/A vssd1 vssd1 vccd1 vccd1 _2830_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_38_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2761_ _2755_/B _2755_/C _2704_/B vssd1 vssd1 vccd1 vccd1 _2762_/C sky130_fd_sc_hd__a21oi_1
XFILLER_0_5_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1712_ _1712_/A _2080_/A vssd1 vssd1 vccd1 vccd1 _2082_/C sky130_fd_sc_hd__nand2_4
X_2692_ _3597_/Q _2867_/C vssd1 vssd1 vccd1 vccd1 _2771_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_41_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1643_ _3628_/Q _1643_/B vssd1 vssd1 vccd1 vccd1 _2669_/B sky130_fd_sc_hd__or2_2
XFILLER_0_67_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2888__A2 _1696_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3313_ _3692_/CLK _3313_/D vssd1 vssd1 vccd1 vccd1 _3313_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3244_ _3322_/CLK _3244_/D vssd1 vssd1 vccd1 vccd1 _3244_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1750__S _1937_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3175_ _3175_/A _3181_/B vssd1 vssd1 vccd1 vccd1 _3175_/X sky130_fd_sc_hd__or2_1
X_2126_ _3725_/Q _2135_/B vssd1 vssd1 vccd1 vccd1 _2126_/Y sky130_fd_sc_hd__nor2_1
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2057_ _2074_/A _2955_/A _2076_/C _2056_/X _1979_/A vssd1 vssd1 vccd1 vccd1 _3626_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_76_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2959_ _2050_/A hold827/X _2959_/S vssd1 vssd1 vccd1 vccd1 _2959_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_32_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold540 _2200_/X vssd1 vssd1 vccd1 vccd1 _3238_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold562 _2625_/X vssd1 vssd1 vccd1 vccd1 _3557_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold551 _3269_/Q vssd1 vssd1 vccd1 vccd1 hold551/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold573 _3399_/Q vssd1 vssd1 vccd1 vccd1 hold573/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold584 _2977_/X vssd1 vssd1 vccd1 vccd1 _3652_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_49_wb_clk_i_A clkbuf_3_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold595 _3639_/Q vssd1 vssd1 vccd1 vccd1 hold595/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout77_A _2652_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1934__S0 _1937_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2264__A0 _3196_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput60 _3333_/Q vssd1 vssd1 vccd1 vccd1 io_out[28] sky130_fd_sc_hd__buf_12
XFILLER_0_53_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2813_ _2811_/A _2812_/X _2811_/Y _2876_/B vssd1 vssd1 vccd1 vccd1 _2813_/X sky130_fd_sc_hd__o211a_1
XANTENNA__2414__B _2612_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2558__A1 _3201_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2744_ _2704_/B _2740_/X _2809_/B _2723_/A _2736_/X vssd1 vssd1 vccd1 vccd1 _2744_/X
+ sky130_fd_sc_hd__o32a_1
X_2675_ _3598_/Q _2868_/C vssd1 vssd1 vccd1 vccd1 _2675_/X sky130_fd_sc_hd__and2_1
X_1626_ _1626_/A vssd1 vssd1 vccd1 vccd1 _1626_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2430__A _2619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3227_ _3727_/CLK _3227_/D vssd1 vssd1 vccd1 vccd1 _3227_/Q sky130_fd_sc_hd__dfxtp_1
X_3158_ _3158_/A _3158_/B vssd1 vssd1 vccd1 vccd1 _3158_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__2494__A0 _2653_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2109_ _3196_/A0 hold189/X _2111_/S vssd1 vssd1 vccd1 vccd1 _2109_/X sky130_fd_sc_hd__mux2_1
X_3089_ _3089_/A _3089_/B _3711_/Q vssd1 vssd1 vccd1 vccd1 _3089_/X sky130_fd_sc_hd__or3b_1
XFILLER_0_91_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2605__A _3192_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_5_wb_clk_i_A clkbuf_leaf_5_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold370 _2656_/X vssd1 vssd1 vccd1 vccd1 _3583_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold381 _3436_/Q vssd1 vssd1 vccd1 vccd1 hold381/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold392 _2090_/X vssd1 vssd1 vccd1 vccd1 _3206_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1907__S0 _2085_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1081 _3602_/Q vssd1 vssd1 vccd1 vccd1 _2984_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1070 _3608_/Q vssd1 vssd1 vccd1 vccd1 _2996_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_59_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_11_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3739_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_70_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1763__A2 _2022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2460_ _3194_/A0 hold333/X _2464_/S vssd1 vssd1 vccd1 vccd1 _2460_/X sky130_fd_sc_hd__mux2_1
X_2391_ _3197_/A0 hold563/X _2392_/S vssd1 vssd1 vccd1 vccd1 _2391_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_48_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3012_ _3014_/A _3684_/Q _3037_/D vssd1 vssd1 vccd1 vccd1 _3012_/X sky130_fd_sc_hd__or3_1
XFILLER_0_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout127_A _1849_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2727_ _3630_/Q _2868_/B _1676_/B vssd1 vssd1 vccd1 vccd1 _2812_/S sky130_fd_sc_hd__o21a_2
XFILLER_0_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2658_ _2658_/A0 hold303/X _2660_/S vssd1 vssd1 vccd1 vccd1 _2658_/X sky130_fd_sc_hd__mux2_1
X_2589_ _2361_/A hold791/X _2590_/S vssd1 vssd1 vccd1 vccd1 _2589_/X sky130_fd_sc_hd__mux2_1
Xfanout113 _2185_/A vssd1 vssd1 vccd1 vccd1 _2244_/A sky130_fd_sc_hd__buf_4
Xfanout102 _2083_/B vssd1 vssd1 vccd1 vccd1 _2854_/B sky130_fd_sc_hd__clkbuf_8
X_1609_ _3325_/Q vssd1 vssd1 vccd1 vccd1 _3772_/A sky130_fd_sc_hd__inv_2
Xfanout135 _3346_/Q vssd1 vssd1 vccd1 vccd1 _2000_/S0 sky130_fd_sc_hd__buf_8
Xfanout146 hold992/X vssd1 vssd1 vccd1 vccd1 _2876_/A sky130_fd_sc_hd__clkbuf_8
Xfanout124 _3348_/Q vssd1 vssd1 vccd1 vccd1 _2289_/A sky130_fd_sc_hd__buf_8
Xfanout157 input18/X vssd1 vssd1 vccd1 vccd1 _3172_/C1 sky130_fd_sc_hd__buf_4
XANTENNA__2467__A0 _3201_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2054__B _3157_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1681__A1 _1979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2245__A _2289_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1960_ hold51/A hold45/A hold91/A _3220_/Q _2085_/B _2014_/A vssd1 vssd1 vccd1 vccd1
+ _1961_/B sky130_fd_sc_hd__mux4_1
X_1891_ _2185_/C _1891_/B vssd1 vssd1 vccd1 vccd1 _1891_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_83_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3630_ _3668_/CLK _3630_/D vssd1 vssd1 vccd1 vccd1 _3630_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_36_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3561_ _3561_/CLK hold28/X vssd1 vssd1 vccd1 vccd1 hold27/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__3186__A1 _2353_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2512_ hold11/X _2361_/A _2513_/S vssd1 vssd1 vccd1 vccd1 hold12/A sky130_fd_sc_hd__mux2_1
XFILLER_0_59_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3492_ _3636_/CLK hold20/X vssd1 vssd1 vccd1 vccd1 hold19/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2443_ hold955/X _2653_/A0 _2443_/S vssd1 vssd1 vccd1 vccd1 _3405_/D sky130_fd_sc_hd__mux2_1
X_2374_ hold37/X _2355_/A _2378_/S vssd1 vssd1 vccd1 vccd1 hold38/A sky130_fd_sc_hd__mux2_1
XANTENNA__2449__A0 _3197_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2621__A0 _2656_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_hold992_A _3310_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output40_A _3613_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2090_ hold391/X _3193_/A0 _2100_/S vssd1 vssd1 vccd1 vccd1 _2090_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_0_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2992_ hold417/X _2480_/A _2992_/S vssd1 vssd1 vccd1 vccd1 _2992_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2603__A0 _2361_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1943_ _3530_/Q _3396_/Q _2244_/B vssd1 vssd1 vccd1 vccd1 _1944_/B sky130_fd_sc_hd__mux2_1
X_1874_ _2074_/A _1873_/X _2028_/S vssd1 vssd1 vccd1 vccd1 _1875_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3613_ _3662_/CLK _3613_/D vssd1 vssd1 vccd1 vccd1 _3613_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_3_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold903 _2077_/X vssd1 vssd1 vccd1 vccd1 _3631_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2906__A1 _2876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3544_ _3545_/CLK _3544_/D vssd1 vssd1 vccd1 vccd1 _3544_/Q sky130_fd_sc_hd__dfxtp_1
Xhold925 _3605_/Q vssd1 vssd1 vccd1 vccd1 hold925/X sky130_fd_sc_hd__buf_1
XFILLER_0_3_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold914 _3709_/Q vssd1 vssd1 vccd1 vccd1 hold914/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold936 _3704_/Q vssd1 vssd1 vccd1 vccd1 hold936/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_3475_ _3733_/CLK hold98/X vssd1 vssd1 vccd1 vccd1 hold97/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold947 _3046_/Y vssd1 vssd1 vccd1 vccd1 _3684_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold969 _3692_/Q vssd1 vssd1 vccd1 vccd1 _1600_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold958 _3138_/X vssd1 vssd1 vccd1 vccd1 _3705_/D sky130_fd_sc_hd__dlygate4sd3_1
X_2426_ hold309/X _2659_/A0 _2427_/S vssd1 vssd1 vccd1 vccd1 _2426_/X sky130_fd_sc_hd__mux2_1
X_2357_ _2357_/A _2363_/B vssd1 vssd1 vccd1 vccd1 _2357_/X sky130_fd_sc_hd__or2_1
XFILLER_0_19_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2288_ _2653_/A0 hold633/X _2288_/S vssd1 vssd1 vccd1 vccd1 _2288_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1989__A _2245_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2437__A3 _2084_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1740__S1 _2479_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2070__A1 _2195_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2070__B2 _2854_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2358__C1 _3058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2833__B1 _2940_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2061__A1 _2046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3260_ _3270_/CLK _3260_/D vssd1 vssd1 vccd1 vccd1 _3260_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3191_ hold59/X _2363_/A _3191_/S vssd1 vssd1 vccd1 vccd1 hold60/A sky130_fd_sc_hd__mux2_1
X_2211_ _2654_/A vssd1 vssd1 vccd1 vccd1 _2633_/B sky130_fd_sc_hd__inv_2
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2142_ _3708_/Q _2142_/B vssd1 vssd1 vccd1 vccd1 _2163_/A sky130_fd_sc_hd__xnor2_1
X_2073_ _2497_/A _2076_/C vssd1 vssd1 vccd1 vccd1 _2073_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_72_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1722__S1 _2245_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2975_ _1627_/A _3613_/Q _2987_/S vssd1 vssd1 vccd1 vccd1 _2975_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_29_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1926_ _1926_/A1 _1769_/Y _1925_/X _2854_/B vssd1 vssd1 vccd1 vccd1 _1927_/B sky130_fd_sc_hd__o22ai_1
X_1857_ _2289_/A _1857_/B vssd1 vssd1 vccd1 vccd1 _1857_/Y sky130_fd_sc_hd__nor2_1
Xhold711 _3555_/Q vssd1 vssd1 vccd1 vccd1 hold711/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold700 _2242_/X vssd1 vssd1 vccd1 vccd1 _3272_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3527_ _3539_/CLK _3527_/D vssd1 vssd1 vccd1 vccd1 _3527_/Q sky130_fd_sc_hd__dfxtp_1
X_1788_ _2006_/A _1787_/X _3348_/Q vssd1 vssd1 vccd1 vccd1 _1788_/X sky130_fd_sc_hd__a21o_1
Xhold733 _3385_/Q vssd1 vssd1 vccd1 vccd1 hold733/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold755 _3286_/Q vssd1 vssd1 vccd1 vccd1 hold755/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold722 _2406_/X vssd1 vssd1 vccd1 vccd1 _3375_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold744 _2337_/X vssd1 vssd1 vccd1 vccd1 _3321_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_39_wb_clk_i_A clkbuf_3_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold788 _2204_/X vssd1 vssd1 vccd1 vccd1 _3244_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold766 _2206_/X vssd1 vssd1 vccd1 vccd1 _3246_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold777 _3336_/Q vssd1 vssd1 vccd1 vccd1 hold777/X sky130_fd_sc_hd__dlygate4sd3_1
X_3458_ _3592_/CLK _3458_/D vssd1 vssd1 vccd1 vccd1 _3458_/Q sky130_fd_sc_hd__dfxtp_1
Xhold799 _3422_/Q vssd1 vssd1 vccd1 vccd1 hold799/X sky130_fd_sc_hd__dlygate4sd3_1
X_2409_ _2656_/A0 hold625/X _2413_/S vssd1 vssd1 vccd1 vccd1 _2409_/X sky130_fd_sc_hd__mux2_1
X_3389_ _3583_/CLK _3389_/D vssd1 vssd1 vccd1 vccd1 _3389_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2291__A1 _2648_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_36_wb_clk_i clkbuf_3_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3322_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_26_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold82 hold82/A vssd1 vssd1 vccd1 vccd1 hold82/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold60 hold60/A vssd1 vssd1 vccd1 vccd1 hold60/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 hold71/A vssd1 vssd1 vccd1 vccd1 hold71/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1952__S1 _2479_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold93 hold93/A vssd1 vssd1 vccd1 vccd1 hold93/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2237__B _2598_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2253__A _3192_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2760_ _2082_/D _2754_/A _2723_/A _2756_/B _2759_/Y vssd1 vssd1 vccd1 vccd1 _2760_/X
+ sky130_fd_sc_hd__o221a_1
X_1711_ _2876_/B _3311_/Q vssd1 vssd1 vccd1 vccd1 _1711_/X sky130_fd_sc_hd__and2_1
X_2691_ _3597_/Q _2867_/C vssd1 vssd1 vccd1 vccd1 _2691_/X sky130_fd_sc_hd__or2_1
XFILLER_0_41_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1642_ _2885_/B _2797_/A _1979_/A vssd1 vssd1 vccd1 vccd1 _1642_/X sky130_fd_sc_hd__and3_1
XFILLER_0_67_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3312_ _3649_/CLK _3312_/D vssd1 vssd1 vccd1 vccd1 _3312_/Q sky130_fd_sc_hd__dfxtp_1
X_3243_ _3649_/CLK _3243_/D vssd1 vssd1 vccd1 vccd1 _3243_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3174_ _2161_/A _3158_/Y _3173_/X _3058_/A vssd1 vssd1 vccd1 vccd1 _3174_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_83_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2428__A _2480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2125_ _3177_/A _2137_/A vssd1 vssd1 vccd1 vccd1 _2135_/B sky130_fd_sc_hd__and2_1
XFILLER_0_76_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2056_ _2717_/A _2062_/B vssd1 vssd1 vccd1 vccd1 _2056_/X sky130_fd_sc_hd__or2_1
XANTENNA__2273__A1 _2022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout157_A input18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2958_ _2046_/A hold815/X _2959_/S vssd1 vssd1 vccd1 vccd1 _2958_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1909_ _3257_/Q _3269_/Q _2085_/B vssd1 vssd1 vccd1 vccd1 _1910_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_4_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2889_ _2876_/A _2884_/Y _2948_/B _2892_/B _2883_/Y vssd1 vssd1 vccd1 vccd1 _2889_/Y
+ sky130_fd_sc_hd__o221ai_1
Xhold530 _2520_/X vssd1 vssd1 vccd1 vccd1 _3467_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold552 _2239_/X vssd1 vssd1 vccd1 vccd1 _3269_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold563 _3362_/Q vssd1 vssd1 vccd1 vccd1 hold563/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold541 _3734_/Q vssd1 vssd1 vccd1 vccd1 hold541/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold574 _2436_/X vssd1 vssd1 vccd1 vccd1 _3399_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold585 _3378_/Q vssd1 vssd1 vccd1 vccd1 hold585/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2733__C1 _2859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold596 _2964_/X vssd1 vssd1 vccd1 vccd1 _3639_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1934__S1 _2245_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2338__A _2619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput61 _2195_/B vssd1 vssd1 vccd1 vccd1 io_out[2] sky130_fd_sc_hd__buf_12
Xoutput50 _3296_/Q vssd1 vssd1 vccd1 vccd1 io_out[19] sky130_fd_sc_hd__buf_12
XANTENNA__2255__A1 _2656_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2812_ _2868_/D hold934/X _2812_/S vssd1 vssd1 vccd1 vccd1 _2812_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_26_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2743_ _2082_/D _2736_/A _2742_/X _2871_/A vssd1 vssd1 vccd1 vccd1 _2743_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_26_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_448 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2674_ _2868_/C _3598_/Q vssd1 vssd1 vccd1 vccd1 _2698_/B sky130_fd_sc_hd__and2b_1
X_1625_ _2185_/C vssd1 vssd1 vccd1 vccd1 _1625_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_1_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2730__A2 _2731_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3226_ _3723_/CLK _3226_/D vssd1 vssd1 vccd1 vccd1 _3226_/Q sky130_fd_sc_hd__dfxtp_2
X_3157_ _3224_/Q _3157_/B _3158_/B vssd1 vssd1 vccd1 vccd1 _3181_/B sky130_fd_sc_hd__and3_4
X_2108_ _3195_/A0 hold725/X _2111_/S vssd1 vssd1 vccd1 vccd1 _2108_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1997__A _2006_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3088_ _3118_/A _3096_/A _2311_/Y _3087_/X vssd1 vssd1 vccd1 vccd1 _3094_/S sky130_fd_sc_hd__o31a_1
X_2039_ _2031_/Y _2037_/X _2038_/X _2495_/A vssd1 vssd1 vccd1 vccd1 _3346_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_49_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1757__B1 _2195_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold371 _3523_/Q vssd1 vssd1 vccd1 vccd1 hold371/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold360 _2107_/X vssd1 vssd1 vccd1 vccd1 _3213_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold393 _3586_/Q vssd1 vssd1 vccd1 vccd1 hold393/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold382 _2482_/X vssd1 vssd1 vccd1 vccd1 _3436_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2485__A1 _3203_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1060 _3677_/Q vssd1 vssd1 vccd1 vccd1 _3024_/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2068__A _2495_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1907__S1 _2014_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1082 _3620_/Q vssd1 vssd1 vccd1 vccd1 _2968_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1693__C1 _1979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1071 _3350_/Q vssd1 vssd1 vccd1 vccd1 hold1071/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_59_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_hold918_A _3595_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_51_wb_clk_i clkbuf_3_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3676_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_2390_ _3196_/A0 hold789/X _2392_/S vssd1 vssd1 vccd1 vccd1 _2390_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_48_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3011_ _3682_/Q _3063_/B vssd1 vssd1 vccd1 vccd1 _3037_/D sky130_fd_sc_hd__nand2b_2
XANTENNA__2476__A1 _3196_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_60 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2726_ _2811_/A _2816_/B vssd1 vssd1 vccd1 vccd1 _2726_/Y sky130_fd_sc_hd__nand2_1
X_2657_ _3195_/A0 hold113/X _2660_/S vssd1 vssd1 vccd1 vccd1 _2657_/X sky130_fd_sc_hd__mux2_1
X_1608_ _3326_/Q vssd1 vssd1 vccd1 vccd1 _3773_/A sky130_fd_sc_hd__inv_2
X_2588_ _3203_/A1 hold797/X _2590_/S vssd1 vssd1 vccd1 vccd1 _2588_/X sky130_fd_sc_hd__mux2_1
Xfanout103 _1767_/Y vssd1 vssd1 vccd1 vccd1 _2731_/A2 sky130_fd_sc_hd__buf_6
Xfanout136 _3346_/Q vssd1 vssd1 vccd1 vccd1 _2289_/B sky130_fd_sc_hd__buf_4
Xfanout114 _1616_/Y vssd1 vssd1 vccd1 vccd1 _2876_/B sky130_fd_sc_hd__buf_4
Xfanout125 _1849_/S1 vssd1 vssd1 vccd1 vccd1 _1981_/S1 sky130_fd_sc_hd__clkbuf_8
Xfanout147 _2961_/A vssd1 vssd1 vccd1 vccd1 _3108_/A sky130_fd_sc_hd__buf_4
XANTENNA__2011__S0 _2085_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3209_ _3308_/CLK hold86/X vssd1 vssd1 vccd1 vccd1 hold85/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1978__A0 _2046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2351__A _2640_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2927__C1 _3103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1825__S0 _1981_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold190 _2109_/X vssd1 vssd1 vccd1 vccd1 _3215_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2245__B _2245_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1969__B1 _2195_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2630__A1 _2658_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1890_ _3529_/Q _3395_/Q _2244_/B vssd1 vssd1 vccd1 vccd1 _1891_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_24_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3560_ _3575_/CLK _3560_/D vssd1 vssd1 vccd1 vccd1 _3560_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2511_ hold121/X _3203_/A1 _2513_/S vssd1 vssd1 vccd1 vccd1 _2511_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2394__A0 _2655_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3491_ _3744_/CLK _3491_/D vssd1 vssd1 vccd1 vccd1 _3491_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2442_ hold971/X _2652_/A0 _2443_/S vssd1 vssd1 vccd1 vccd1 _3404_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_59_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2373_ hold197/X _2648_/A0 _2378_/S vssd1 vssd1 vccd1 vccd1 _2373_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_75_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2385__A0 _2660_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2709_ _2803_/B _2803_/C _2709_/C _2779_/A vssd1 vssd1 vccd1 vccd1 _2809_/A sky130_fd_sc_hd__and4_1
Xscrapcpu_170 vssd1 vssd1 vccd1 vccd1 scrapcpu_170/HI io_oeb[28] sky130_fd_sc_hd__conb_1
X_3689_ _3724_/CLK _3689_/D vssd1 vssd1 vccd1 vccd1 _3689_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2346__A _3108_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1820__C1 _1979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2991_ hold435/X _2228_/C _2992_/S vssd1 vssd1 vccd1 vccd1 _2991_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_56_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1942_ _2244_/A _1942_/B vssd1 vssd1 vccd1 vccd1 _1942_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_16_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1873_ _2994_/A1 _1769_/Y _1872_/X _2854_/B vssd1 vssd1 vccd1 vccd1 _1873_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_9_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3612_ _3649_/CLK _3612_/D vssd1 vssd1 vccd1 vccd1 _3612_/Q sky130_fd_sc_hd__dfxtp_4
Xhold904 _3598_/Q vssd1 vssd1 vccd1 vccd1 _2861_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_0_24_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_29_wb_clk_i_A clkbuf_3_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_3543_ _3543_/CLK _3543_/D vssd1 vssd1 vccd1 vccd1 _3543_/Q sky130_fd_sc_hd__dfxtp_1
Xhold926 _2848_/X vssd1 vssd1 vccd1 vccd1 _3605_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold915 _3146_/X vssd1 vssd1 vccd1 vccd1 _3709_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold937 _3162_/X vssd1 vssd1 vccd1 vccd1 _3716_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3474_ _3592_/CLK hold18/X vssd1 vssd1 vccd1 vccd1 hold17/A sky130_fd_sc_hd__dfxtp_1
Xhold948 _3714_/Q vssd1 vssd1 vccd1 vccd1 hold948/X sky130_fd_sc_hd__buf_1
Xhold959 _3618_/Q vssd1 vssd1 vccd1 vccd1 _2914_/B sky130_fd_sc_hd__buf_1
XANTENNA__2119__A0 _2653_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2425_ hold277/X _2658_/A0 _2427_/S vssd1 vssd1 vccd1 vccd1 _2425_/X sky130_fd_sc_hd__mux2_1
X_2356_ hold994/X _2351_/Y _2355_/X _3058_/A vssd1 vssd1 vccd1 vccd1 _3329_/D sky130_fd_sc_hd__o211a_1
X_2287_ _2361_/A hold577/X _2288_/S vssd1 vssd1 vccd1 vccd1 _2287_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_29_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1869__C1 _1922_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2076__A _2076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2061__A2 _2955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2015__S _2085_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2349__A0 _2653_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2210_ _2228_/A _2479_/B _2479_/C vssd1 vssd1 vccd1 vccd1 _2654_/A sky130_fd_sc_hd__and3_4
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3190_ hold81/X _2361_/A _3191_/S vssd1 vssd1 vccd1 vccd1 hold82/A sky130_fd_sc_hd__mux2_1
X_2141_ _2154_/B _2141_/B vssd1 vssd1 vccd1 vccd1 _2142_/B sky130_fd_sc_hd__or2_1
XFILLER_0_56_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2072_ _2067_/S _2070_/X _2071_/X _2495_/A vssd1 vssd1 vccd1 vccd1 _2072_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_72_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2974_ hold793/X _3612_/Q _2987_/S vssd1 vssd1 vccd1 vccd1 _2974_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2588__A0 _3203_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1925_ hold805/X _2731_/A2 _2867_/A _1713_/X vssd1 vssd1 vccd1 vccd1 _1925_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_16_104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_6_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3636_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_44_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1856_ _3304_/Q _3274_/Q _3206_/Q _3218_/Q _2085_/B _2014_/A vssd1 vssd1 vccd1 vccd1
+ _1857_/B sky130_fd_sc_hd__mux4_1
Xhold712 _2623_/X vssd1 vssd1 vccd1 vccd1 _3555_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1787_ _3461_/Q _3593_/Q _2244_/B vssd1 vssd1 vccd1 vccd1 _1787_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_71_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold701 _3509_/Q vssd1 vssd1 vccd1 vccd1 hold701/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3526_ _3561_/CLK _3526_/D vssd1 vssd1 vccd1 vccd1 _3526_/Q sky130_fd_sc_hd__dfxtp_1
Xhold723 _3516_/Q vssd1 vssd1 vccd1 vccd1 hold723/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold745 _3318_/Q vssd1 vssd1 vccd1 vccd1 hold745/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold734 _2418_/X vssd1 vssd1 vccd1 vccd1 _3385_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold767 _3673_/Q vssd1 vssd1 vccd1 vccd1 hold767/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold756 _2261_/X vssd1 vssd1 vccd1 vccd1 _3286_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold778 _2368_/X vssd1 vssd1 vccd1 vccd1 _3336_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3457_ _3745_/CLK _3457_/D vssd1 vssd1 vccd1 vccd1 _3457_/Q sky130_fd_sc_hd__dfxtp_1
Xhold789 _3361_/Q vssd1 vssd1 vccd1 vccd1 hold789/X sky130_fd_sc_hd__dlygate4sd3_1
X_2408_ _2655_/A0 hold127/X _2413_/S vssd1 vssd1 vccd1 vccd1 _2408_/X sky130_fd_sc_hd__mux2_1
X_3388_ _3735_/CLK _3388_/D vssd1 vssd1 vccd1 vccd1 _3388_/Q sky130_fd_sc_hd__dfxtp_1
X_2339_ _2648_/A0 _2619_/A _2647_/B _3108_/A vssd1 vssd1 vccd1 vccd1 _2339_/X sky130_fd_sc_hd__a31o_1
XANTENNA__2579__A0 _2656_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2751__A0 _2867_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold50 hold50/A vssd1 vssd1 vccd1 vccd1 hold50/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold61 hold61/A vssd1 vssd1 vccd1 vccd1 hold61/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 hold72/A vssd1 vssd1 vccd1 vccd1 hold72/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 hold83/A vssd1 vssd1 vccd1 vccd1 hold83/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 hold94/A vssd1 vssd1 vccd1 vccd1 hold94/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_85_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1710_ _1824_/A _1824_/B _3045_/B _2071_/D vssd1 vssd1 vccd1 vccd1 _1819_/A sky130_fd_sc_hd__or4_2
X_2690_ _3597_/Q _2867_/C vssd1 vssd1 vccd1 vccd1 _2690_/X sky130_fd_sc_hd__and2_1
X_1641_ _3045_/B _3048_/B _3096_/B vssd1 vssd1 vccd1 vccd1 _1685_/B sky130_fd_sc_hd__or3_4
XFILLER_0_41_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3311_ _3649_/CLK _3311_/D vssd1 vssd1 vccd1 vccd1 _3311_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3242_ _3637_/CLK _3242_/D vssd1 vssd1 vccd1 vccd1 _3242_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3173_ _3722_/Q _3181_/B vssd1 vssd1 vccd1 vccd1 _3173_/X sky130_fd_sc_hd__or2_1
X_2124_ _3175_/A _3722_/Q _2155_/A vssd1 vssd1 vccd1 vccd1 _2137_/A sky130_fd_sc_hd__and3_1
XFILLER_0_83_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2428__B _3351_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2055_ _2955_/A _2076_/C vssd1 vssd1 vccd1 vccd1 _2062_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_76_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2273__A2 _2245_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2444__A _2647_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2957_ _2076_/A _1922_/A _2959_/S vssd1 vssd1 vccd1 vccd1 _2957_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2025__A2 _1922_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2888_ _2876_/A _1696_/Y _2886_/A vssd1 vssd1 vccd1 vccd1 _2948_/B sky130_fd_sc_hd__o21ai_4
X_1908_ _2085_/A _1908_/B vssd1 vssd1 vccd1 vccd1 _1908_/Y sky130_fd_sc_hd__nor2_1
X_1839_ hold93/A _3394_/Q _2244_/B vssd1 vssd1 vccd1 vccd1 _1840_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_4_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold520 _2988_/X vssd1 vssd1 vccd1 vccd1 _3663_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold531 _3428_/Q vssd1 vssd1 vccd1 vccd1 hold531/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold553 _3251_/Q vssd1 vssd1 vccd1 vccd1 hold553/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold542 _3193_/X vssd1 vssd1 vccd1 vccd1 _3734_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold586 _2410_/X vssd1 vssd1 vccd1 vccd1 _3378_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3509_ _3739_/CLK _3509_/D vssd1 vssd1 vccd1 vccd1 _3509_/Q sky130_fd_sc_hd__dfxtp_1
Xhold564 _2391_/X vssd1 vssd1 vccd1 vccd1 _3362_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold575 _3406_/Q vssd1 vssd1 vccd1 vccd1 hold575/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold597 _3450_/Q vssd1 vssd1 vccd1 vccd1 hold597/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2619__A _2619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3185__A _3192_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput51 _3612_/Q vssd1 vssd1 vccd1 vccd1 io_out[1] sky130_fd_sc_hd__buf_12
Xoutput40 _3613_/Q vssd1 vssd1 vccd1 vccd1 io_out[0] sky130_fd_sc_hd__buf_12
Xoutput62 _3676_/Q vssd1 vssd1 vccd1 vccd1 io_out[30] sky130_fd_sc_hd__buf_12
XANTENNA__3204__A1 _2361_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2811_ _2811_/A _2843_/B vssd1 vssd1 vccd1 vccd1 _2811_/Y sky130_fd_sc_hd__nand2_1
X_2742_ _3628_/Q _2742_/B _2742_/C vssd1 vssd1 vccd1 vccd1 _2742_/X sky130_fd_sc_hd__or3_1
XFILLER_0_81_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3095__A _3108_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2673_ _2851_/A _2673_/B vssd1 vssd1 vccd1 vccd1 _2802_/A sky130_fd_sc_hd__or2_1
XFILLER_0_41_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1624_ _3348_/Q vssd1 vssd1 vccd1 vccd1 _2185_/A sky130_fd_sc_hd__inv_2
XANTENNA__2191__A1 _2652_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3225_ _3727_/CLK _3225_/D vssd1 vssd1 vccd1 vccd1 _3225_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3156_ hold948/X _3131_/X _3155_/X _3103_/A vssd1 vssd1 vccd1 vccd1 _3714_/D sky130_fd_sc_hd__o211a_1
X_3087_ _3677_/Q _3183_/B _2169_/B _2303_/X _3080_/A vssd1 vssd1 vccd1 vccd1 _3087_/X
+ sky130_fd_sc_hd__o221a_1
X_2107_ _3194_/A0 hold359/X _2111_/S vssd1 vssd1 vccd1 vccd1 _2107_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2038_ _2074_/A _2050_/B vssd1 vssd1 vccd1 vccd1 _2038_/X sky130_fd_sc_hd__or2_1
XFILLER_0_49_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1757__A1 _2480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold361 _3518_/Q vssd1 vssd1 vccd1 vccd1 hold361/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold350 _2973_/X vssd1 vssd1 vccd1 vccd1 _3648_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold372 _2586_/X vssd1 vssd1 vccd1 vccd1 _3523_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold394 _2659_/X vssd1 vssd1 vccd1 vccd1 _3586_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold383 _3580_/Q vssd1 vssd1 vccd1 vccd1 hold383/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout82_A _2359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1050 _3613_/Q vssd1 vssd1 vccd1 vccd1 _2874_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1072 _3601_/Q vssd1 vssd1 vccd1 vccd1 _2983_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1061 _3629_/Q vssd1 vssd1 vccd1 vccd1 _1643_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1083 _3615_/Q vssd1 vssd1 vccd1 vccd1 _2963_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2890__C1 _3103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2084__A _2084_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3198__A0 _3198_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_20_wb_clk_i clkbuf_3_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3570_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_3_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3010_ _3124_/A _3010_/B vssd1 vssd1 vccd1 vccd1 _3010_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_64_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3774_ _3774_/A vssd1 vssd1 vccd1 vccd1 _3774_/X sky130_fd_sc_hd__buf_1
XFILLER_0_89_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2725_ _2713_/X _2718_/X _2724_/X _2710_/Y vssd1 vssd1 vccd1 vccd1 _2816_/B sky130_fd_sc_hd__a31o_1
X_2656_ _2656_/A0 hold369/X _2660_/S vssd1 vssd1 vccd1 vccd1 _2656_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_14_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1607_ _3327_/Q vssd1 vssd1 vccd1 vccd1 _3774_/A sky130_fd_sc_hd__inv_2
X_2587_ _3195_/A0 hold769/X _2590_/S vssd1 vssd1 vccd1 vccd1 _2587_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_10_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout104 _1766_/Y vssd1 vssd1 vccd1 vccd1 _2940_/B2 sky130_fd_sc_hd__buf_4
XFILLER_0_1_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout115 _1616_/Y vssd1 vssd1 vccd1 vccd1 _1712_/A sky130_fd_sc_hd__buf_4
Xfanout126 _1849_/S1 vssd1 vssd1 vccd1 vccd1 _1760_/B sky130_fd_sc_hd__clkbuf_4
Xfanout137 _1954_/S vssd1 vssd1 vccd1 vccd1 _2085_/B sky130_fd_sc_hd__buf_6
Xfanout148 _1620_/Y vssd1 vssd1 vccd1 vccd1 _2961_/A sky130_fd_sc_hd__clkbuf_4
X_3208_ _3666_/CLK hold92/X vssd1 vssd1 vccd1 vccd1 hold91/A sky130_fd_sc_hd__dfxtp_1
X_3139_ _2904_/A _2886_/A _3137_/C vssd1 vssd1 vccd1 vccd1 _3139_/X sky130_fd_sc_hd__a21o_1
XANTENNA__2011__S1 _2014_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1825__S1 _1981_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold180 _2572_/X vssd1 vssd1 vccd1 vccd1 _3511_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold191 _3530_/Q vssd1 vssd1 vccd1 vccd1 hold191/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_34_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2245__C _2245_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2542__A _2619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3490_ _3744_/CLK _3490_/D vssd1 vssd1 vccd1 vccd1 _3490_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_19_wb_clk_i_A clkbuf_3_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_2510_ hold287/X _2357_/A _2513_/S vssd1 vssd1 vccd1 vccd1 _2510_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_11_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2441_ hold881/X _2651_/A0 _2443_/S vssd1 vssd1 vccd1 vccd1 _2441_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_11_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2372_ _2372_/A _2612_/B vssd1 vssd1 vccd1 vccd1 _2378_/S sky130_fd_sc_hd__nor2_2
XFILLER_0_78_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2708_ _2709_/C _2779_/A vssd1 vssd1 vccd1 vccd1 _2708_/Y sky130_fd_sc_hd__nand2_1
X_3688_ _3692_/CLK _3688_/D vssd1 vssd1 vccd1 vccd1 _3688_/Q sky130_fd_sc_hd__dfxtp_1
Xscrapcpu_160 vssd1 vssd1 vccd1 vccd1 scrapcpu_160/HI io_oeb[2] sky130_fd_sc_hd__conb_1
Xscrapcpu_171 vssd1 vssd1 vccd1 vccd1 scrapcpu_171/HI io_oeb[30] sky130_fd_sc_hd__conb_1
X_2639_ _2660_/A0 hold511/X _2639_/S vssd1 vssd1 vccd1 vccd1 _2639_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_84_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2376__A1 _2651_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1982__S0 _1760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2990_ hold589/X _2085_/A _2992_/S vssd1 vssd1 vccd1 vccd1 _2990_/X sky130_fd_sc_hd__mux2_1
X_1941_ _3730_/Q _3476_/Q hold5/A _3426_/Q _1996_/S _2185_/C vssd1 vssd1 vccd1 vccd1
+ _1942_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_56_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1811__B1 _2195_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1872_ hold239/X _2731_/A2 _2701_/B _1713_/X vssd1 vssd1 vccd1 vccd1 _1872_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_9_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3611_ _3646_/CLK _3611_/D vssd1 vssd1 vccd1 vccd1 _3611_/Q sky130_fd_sc_hd__dfxtp_1
X_3542_ _3587_/CLK _3542_/D vssd1 vssd1 vccd1 vccd1 _3542_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold916 _3243_/Q vssd1 vssd1 vccd1 vccd1 _1824_/A sky130_fd_sc_hd__clkbuf_2
Xhold905 _2799_/X vssd1 vssd1 vccd1 vccd1 _3598_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold927 _3707_/Q vssd1 vssd1 vccd1 vccd1 hold927/X sky130_fd_sc_hd__buf_1
X_3473_ _3744_/CLK _3473_/D vssd1 vssd1 vccd1 vccd1 _3473_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1616__A _2797_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold949 _3182_/X vssd1 vssd1 vccd1 vccd1 _3726_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold938 _3676_/Q vssd1 vssd1 vccd1 vccd1 _2885_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_51_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2424_ hold83/X _3195_/A0 _2427_/S vssd1 vssd1 vccd1 vccd1 hold84/A sky130_fd_sc_hd__mux2_1
XFILLER_0_86_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2355_ _2355_/A _2363_/B vssd1 vssd1 vccd1 vccd1 _2355_/X sky130_fd_sc_hd__or2_1
X_2286_ _2651_/A0 hold659/X _2288_/S vssd1 vssd1 vccd1 vccd1 _2286_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2827__C1 _2859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2530__A1 _3201_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2357__A _2357_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2833__A2 _1696_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2597__A1 _2099_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2140_ _3719_/Q _2146_/A _3720_/Q vssd1 vssd1 vccd1 vccd1 _2141_/B sky130_fd_sc_hd__a21oi_1
X_2071_ _2071_/A _2076_/A _3045_/B _2071_/D vssd1 vssd1 vccd1 vccd1 _2071_/X sky130_fd_sc_hd__or4_1
XFILLER_0_88_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2285__A0 _2650_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2973_ hold349/X _3625_/Q _2999_/S vssd1 vssd1 vccd1 vccd1 _2973_/X sky130_fd_sc_hd__mux2_1
X_1924_ _2687_/B vssd1 vssd1 vccd1 vccd1 _2867_/A sky130_fd_sc_hd__inv_2
XFILLER_0_29_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1855_ _2244_/A _1851_/Y _1853_/X _1854_/Y vssd1 vssd1 vccd1 vccd1 _1855_/X sky130_fd_sc_hd__a31o_1
X_1786_ _3533_/Q _3399_/Q _1996_/S vssd1 vssd1 vccd1 vccd1 _1786_/X sky130_fd_sc_hd__mux2_1
Xhold702 _2569_/X vssd1 vssd1 vccd1 vccd1 _3509_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3525_ _3561_/CLK _3525_/D vssd1 vssd1 vccd1 vccd1 _3525_/Q sky130_fd_sc_hd__dfxtp_1
Xhold735 _3354_/Q vssd1 vssd1 vccd1 vccd1 hold735/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold713 _3504_/Q vssd1 vssd1 vccd1 vccd1 hold713/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold724 _2578_/X vssd1 vssd1 vccd1 vccd1 _3516_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold746 _2334_/X vssd1 vssd1 vccd1 vccd1 _3318_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold757 _3527_/Q vssd1 vssd1 vccd1 vccd1 hold757/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold779 _3552_/Q vssd1 vssd1 vccd1 vccd1 hold779/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold768 _2998_/X vssd1 vssd1 vccd1 vccd1 _3673_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3456_ _3728_/CLK _3456_/D vssd1 vssd1 vccd1 vccd1 _3456_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1780__S _1937_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2512__A1 _2361_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2407_ _2407_/A _2598_/A vssd1 vssd1 vccd1 vccd1 _2413_/S sky130_fd_sc_hd__nand2_4
XFILLER_0_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3387_ _3387_/CLK _3387_/D vssd1 vssd1 vccd1 vccd1 _3387_/Q sky130_fd_sc_hd__dfxtp_1
X_2338_ _2619_/A _2647_/B vssd1 vssd1 vccd1 vccd1 _2349_/S sky130_fd_sc_hd__nand2_2
X_2269_ _2022_/A _2245_/C _2648_/A0 _2268_/X _3058_/A vssd1 vssd1 vccd1 vccd1 _3292_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_46_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2028__A0 _2050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2640__A _2640_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2200__A0 _2658_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2219__A_N _2000_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold40 hold40/A vssd1 vssd1 vccd1 vccd1 hold40/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 hold62/A vssd1 vssd1 vccd1 vccd1 hold62/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 hold51/A vssd1 vssd1 vccd1 vccd1 hold51/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 hold73/A vssd1 vssd1 vccd1 vccd1 hold73/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2087__A _2087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold84 hold84/A vssd1 vssd1 vccd1 vccd1 hold84/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 hold95/A vssd1 vssd1 vccd1 vccd1 hold95/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2267__B1 _2022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_45_wb_clk_i clkbuf_3_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3702_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_13_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1640_ _3045_/B _3048_/B _1640_/C vssd1 vssd1 vccd1 vccd1 _2960_/A sky130_fd_sc_hd__nor3_4
XANTENNA__2990__A1 _2085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3310_ _3649_/CLK _3310_/D vssd1 vssd1 vccd1 vccd1 _3310_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_21_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3241_ _3637_/CLK _3241_/D vssd1 vssd1 vccd1 vccd1 _3241_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3172_ _3709_/Q _3158_/Y hold873/X _3172_/C1 vssd1 vssd1 vccd1 vccd1 _3172_/X sky130_fd_sc_hd__o211a_1
X_2123_ _3721_/Q _2154_/B vssd1 vssd1 vccd1 vccd1 _2155_/A sky130_fd_sc_hd__and2_1
XANTENNA__2428__C _2428_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2054_ _2054_/A _3157_/B vssd1 vssd1 vccd1 vccd1 _2076_/C sky130_fd_sc_hd__nand2_2
XFILLER_0_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2273__A3 _2650_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2956_ _2074_/A _1870_/A _2959_/S vssd1 vssd1 vccd1 vccd1 _2956_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_32_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2887_ _2876_/A _1696_/Y _2886_/A vssd1 vssd1 vccd1 vccd1 _2935_/A sky130_fd_sc_hd__o21a_2
XFILLER_0_32_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1907_ hold55/A hold75/A _3207_/Q _3219_/Q _2085_/B _2014_/A vssd1 vssd1 vccd1 vccd1
+ _1908_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_89_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1838_ _1889_/A _1838_/B vssd1 vssd1 vccd1 vccd1 _1838_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_25_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold510 _2384_/X vssd1 vssd1 vccd1 vccd1 _3356_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold532 _2470_/X vssd1 vssd1 vccd1 vccd1 _3428_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold521 _3477_/Q vssd1 vssd1 vccd1 vccd1 hold521/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold554 _2214_/X vssd1 vssd1 vccd1 vccd1 _3251_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold543 _3270_/Q vssd1 vssd1 vccd1 vccd1 hold543/X sky130_fd_sc_hd__dlygate4sd3_1
X_1769_ _1713_/X _2731_/A2 _2854_/B vssd1 vssd1 vccd1 vccd1 _1769_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__2733__A1 hold908/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold1062_A _3346_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold587 _3427_/Q vssd1 vssd1 vccd1 vccd1 hold587/X sky130_fd_sc_hd__dlygate4sd3_1
X_3508_ _3545_/CLK _3508_/D vssd1 vssd1 vccd1 vccd1 _3508_/Q sky130_fd_sc_hd__dfxtp_1
Xhold565 _3655_/Q vssd1 vssd1 vccd1 vccd1 hold565/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold576 _2445_/X vssd1 vssd1 vccd1 vccd1 _3406_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3439_ _3539_/CLK _3439_/D vssd1 vssd1 vccd1 vccd1 _3439_/Q sky130_fd_sc_hd__dfxtp_1
Xhold598 _2501_/X vssd1 vssd1 vccd1 vccd1 _3450_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput30 _3621_/Q vssd1 vssd1 vccd1 vccd1 io_oeb[31] sky130_fd_sc_hd__buf_12
Xoutput41 _3401_/Q vssd1 vssd1 vccd1 vccd1 io_out[10] sky130_fd_sc_hd__buf_12
Xoutput52 _3297_/Q vssd1 vssd1 vccd1 vccd1 io_out[20] sky130_fd_sc_hd__buf_12
Xoutput63 _3692_/Q vssd1 vssd1 vccd1 vccd1 io_out[3] sky130_fd_sc_hd__buf_12
XANTENNA__2660__A0 _2660_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2810_ _2718_/B _2804_/Y _2805_/X _2807_/Y _2809_/X vssd1 vssd1 vccd1 vccd1 _2843_/B
+ sky130_fd_sc_hd__o311a_1
XANTENNA__2412__A0 _2659_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2741_ _2741_/A _2741_/B vssd1 vssd1 vccd1 vccd1 _2809_/B sky130_fd_sc_hd__or2_2
XFILLER_0_5_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2672_ _3599_/Q _2868_/D vssd1 vssd1 vccd1 vccd1 _2673_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1623_ _2195_/B vssd1 vssd1 vccd1 vccd1 _2228_/B sky130_fd_sc_hd__inv_2
XFILLER_0_1_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1624__A _3348_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3224_ _3702_/CLK _3224_/D vssd1 vssd1 vccd1 vccd1 _3224_/Q sky130_fd_sc_hd__dfxtp_1
.ends

