// This is the unpowered netlist.
module multiplexer (io_in_0,
    rst_scrapcpu,
    rst_vliw,
    rst_z80,
    wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    custom_settings,
    io_oeb,
    io_oeb_scrapcpu,
    io_oeb_vliw,
    io_oeb_z80,
    io_out,
    io_out_scrapcpu,
    io_out_vliw,
    io_out_z80,
    la_data_out,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o);
 input io_in_0;
 output rst_scrapcpu;
 output rst_vliw;
 output rst_z80;
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 output [31:0] custom_settings;
 output [37:0] io_oeb;
 input [35:0] io_oeb_scrapcpu;
 input [35:0] io_oeb_vliw;
 input [35:0] io_oeb_z80;
 output [37:0] io_out;
 input [35:0] io_out_scrapcpu;
 input [35:0] io_out_vliw;
 input [35:0] io_out_z80;
 output [39:0] la_data_out;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;

 wire net482;
 wire net479;
 wire net480;
 wire net483;
 wire net481;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire clknet_0_wb_clk_i;
 wire clknet_4_0_0_wb_clk_i;
 wire clknet_4_10_0_wb_clk_i;
 wire clknet_4_11_0_wb_clk_i;
 wire clknet_4_12_0_wb_clk_i;
 wire clknet_4_13_0_wb_clk_i;
 wire clknet_4_14_0_wb_clk_i;
 wire clknet_4_15_0_wb_clk_i;
 wire clknet_4_1_0_wb_clk_i;
 wire clknet_4_2_0_wb_clk_i;
 wire clknet_4_3_0_wb_clk_i;
 wire clknet_4_4_0_wb_clk_i;
 wire clknet_4_5_0_wb_clk_i;
 wire clknet_4_6_0_wb_clk_i;
 wire clknet_4_7_0_wb_clk_i;
 wire clknet_4_8_0_wb_clk_i;
 wire clknet_4_9_0_wb_clk_i;
 wire \design_select[0] ;
 wire \design_select[1] ;
 wire \design_select[2] ;
 wire \design_select[3] ;
 wire net1;
 wire net10;
 wire net100;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net101;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net102;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net103;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net104;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net105;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net106;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net107;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net108;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net109;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net11;
 wire net110;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net111;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net112;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net113;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net114;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net115;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net116;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net117;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net118;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net119;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net12;
 wire net120;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net121;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net122;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net123;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net124;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net125;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net126;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net48;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net79;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net8;
 wire net80;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net81;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net82;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net83;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net84;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net85;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net86;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net87;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net88;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net89;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net9;
 wire net90;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net91;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net92;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net93;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net94;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net95;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net96;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net97;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net98;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net99;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire \wb_counter[0] ;
 wire \wb_counter[10] ;
 wire \wb_counter[11] ;
 wire \wb_counter[12] ;
 wire \wb_counter[13] ;
 wire \wb_counter[14] ;
 wire \wb_counter[15] ;
 wire \wb_counter[16] ;
 wire \wb_counter[17] ;
 wire \wb_counter[18] ;
 wire \wb_counter[19] ;
 wire \wb_counter[1] ;
 wire \wb_counter[20] ;
 wire \wb_counter[21] ;
 wire \wb_counter[22] ;
 wire \wb_counter[23] ;
 wire \wb_counter[24] ;
 wire \wb_counter[26] ;
 wire \wb_counter[27] ;
 wire \wb_counter[28] ;
 wire \wb_counter[29] ;
 wire \wb_counter[2] ;
 wire \wb_counter[30] ;
 wire \wb_counter[31] ;
 wire \wb_counter[3] ;
 wire \wb_counter[4] ;
 wire \wb_counter[5] ;
 wire \wb_counter[6] ;
 wire \wb_counter[7] ;
 wire \wb_counter[8] ;
 wire \wb_counter[9] ;
 wire wb_feedback_delay;
 wire wb_override_act;
 wire wb_rst_override;
 wire \wbs_adr_delaybuff[0] ;
 wire \wbs_adr_delaybuff[1] ;
 wire \wbs_adr_delaybuff[2] ;
 wire \wbs_adr_delaybuff[3] ;
 wire \wbs_dat_delaybuff[0] ;
 wire \wbs_dat_delaybuff[10] ;
 wire \wbs_dat_delaybuff[11] ;
 wire \wbs_dat_delaybuff[12] ;
 wire \wbs_dat_delaybuff[13] ;
 wire \wbs_dat_delaybuff[14] ;
 wire \wbs_dat_delaybuff[15] ;
 wire \wbs_dat_delaybuff[16] ;
 wire \wbs_dat_delaybuff[17] ;
 wire \wbs_dat_delaybuff[18] ;
 wire \wbs_dat_delaybuff[19] ;
 wire \wbs_dat_delaybuff[1] ;
 wire \wbs_dat_delaybuff[20] ;
 wire \wbs_dat_delaybuff[21] ;
 wire \wbs_dat_delaybuff[22] ;
 wire \wbs_dat_delaybuff[23] ;
 wire \wbs_dat_delaybuff[24] ;
 wire \wbs_dat_delaybuff[25] ;
 wire \wbs_dat_delaybuff[26] ;
 wire \wbs_dat_delaybuff[27] ;
 wire \wbs_dat_delaybuff[28] ;
 wire \wbs_dat_delaybuff[29] ;
 wire \wbs_dat_delaybuff[2] ;
 wire \wbs_dat_delaybuff[30] ;
 wire \wbs_dat_delaybuff[31] ;
 wire \wbs_dat_delaybuff[3] ;
 wire \wbs_dat_delaybuff[4] ;
 wire \wbs_dat_delaybuff[5] ;
 wire \wbs_dat_delaybuff[6] ;
 wire \wbs_dat_delaybuff[7] ;
 wire \wbs_dat_delaybuff[8] ;
 wire \wbs_dat_delaybuff[9] ;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA__0396__A (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__0397__A0 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__0399__A_N (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA__0399__B (.DIODE(net580));
 sky130_fd_sc_hd__diode_2 ANTENNA__0399__C (.DIODE(net572));
 sky130_fd_sc_hd__diode_2 ANTENNA__0400__A (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__0400__B (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__0401__A_N (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA__0401__B (.DIODE(net572));
 sky130_fd_sc_hd__diode_2 ANTENNA__0401__C (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA__0402__A (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__0402__B (.DIODE(_0116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0403__A (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA__0403__B (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA__0403__C (.DIODE(net572));
 sky130_fd_sc_hd__diode_2 ANTENNA__0404__A (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__0404__B (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__0405__A1 (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA__0405__A2 (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA__0405__B1 (.DIODE(net572));
 sky130_fd_sc_hd__diode_2 ANTENNA__0406__A1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__0406__B1 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__0407__A1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__0407__A2 (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 ANTENNA__0408__A1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__0408__B1 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__0409__A1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__0409__A2 (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 ANTENNA__0410__A1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__0410__B1 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__0411__A1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__0411__A2 (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 ANTENNA__0412__A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__0412__B1 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__0413__A1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__0413__A2 (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 ANTENNA__0414__A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__0414__B1 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__0415__A1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__0415__A2 (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 ANTENNA__0416__A1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__0416__B1 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__0417__A1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__0417__A2 (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 ANTENNA__0418__A1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__0418__B1 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__0419__A1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__0419__A2 (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 ANTENNA__0420__A1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__0420__B1 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__0421__A1 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__0421__A2 (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 ANTENNA__0422__A1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__0422__B1 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__0423__A1 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__0423__A2 (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 ANTENNA__0424__A1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__0425__A1 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__0426__A1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__0427__A1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__0428__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__0429__A1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__0430__A1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__0431__A1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__0432__A1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__0433__A1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__0434__A1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__0435__A1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__0436__A1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__0437__A1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__0438__A1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__0439__A1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__0440__A1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__0440__B1 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__0441__A1 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__0441__A2 (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 ANTENNA__0442__A1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__0442__B1 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__0443__A1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__0444__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__0445__A1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__0446__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__0447__A1 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__0448__A1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__0449__A1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__0450__A1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__0451__A1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__0452__A1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__0453__A1 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__0454__A1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__0455__A1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__0456__A1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__0457__A1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__0457__A2 (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 ANTENNA__0458__A1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__0459__A1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__0460__B2 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__0461__A1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__0462__B2 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__0463__A1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__0464__B2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__0465__A1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__0466__B2 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__0467__A1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__0468__B2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__0469__A1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__0470__B2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__0471__A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__0472__B2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__0473__A1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__0474__B2 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__0475__A1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__0476__B2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__0477__A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__0478__B2 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__0479__A1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__0480__B2 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__0481__A1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__0482__B2 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__0483__A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__0484__B2 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__0485__A1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__0486__B2 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__0487__A1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__0488__B2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__0489__A1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__0490__B2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__0491__A1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__0492__A2 (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__0492__B1 (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__0492__B2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__0493__A1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__0493__A2 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__0494__A2 (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__0494__B1 (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__0494__B2 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__0495__A1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__0495__A2 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__0496__A2 (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__0496__B1 (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__0496__B2 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__0497__A1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__0497__A2 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__0498__B1 (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__0498__B2 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__0499__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__0499__A2 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__0500__B1 (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__0500__B2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__0501__A1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__0501__A2 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__0502__B1 (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__0502__B2 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__0503__A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__0503__A2 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__0504__B1 (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__0504__B2 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__0505__A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__0505__A2 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__0506__B1 (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__0506__B2 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__0507__A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__0507__A2 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__0508__B1 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA__0508__B2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__0509__A1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__0509__A2 (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA__0510__B1 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA__0510__B2 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__0511__A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__0511__A2 (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA__0512__B1 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA__0512__B2 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__0513__A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__0513__A2 (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA__0514__B1 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA__0514__B2 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__0515__A1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__0515__A2 (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA__0516__B1 (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__0516__B2 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__0517__A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__0517__A2 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__0518__B1 (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__0518__B2 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__0519__A1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__0519__A2 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__0520__B1 (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__0520__B2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__0521__A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__0521__A2 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__0522__B1 (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__0522__B2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__0523__A1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__0523__A2 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__0524__B1 (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__0524__B2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__0525__A1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__0525__A2 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__0526__B1 (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__0526__B2 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__0527__A1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__0527__A2 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__0528__B1 (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__0528__B2 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__0529__A1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__0529__A2 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA__0530__A2 (.DIODE(_0115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0530__B1 (.DIODE(_0117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0530__B2 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__0531__A1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__0531__A2 (.DIODE(_0116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0532__A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__0532__A2 (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__0532__B1 (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA__0533__A1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__0533__A2 (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA__0534__A1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__0534__A2 (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__0534__B1 (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA__0535__A1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__0536__A1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__0536__A2 (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__0536__B1 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA__0537__A1 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__0537__A2 (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA__0538__A1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__0538__A2 (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__0538__B1 (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA__0539__A1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__0540__A1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__0540__A2 (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__0540__B1 (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA__0541__A1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__0542__A1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__0542__A2 (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__0542__B1 (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA__0543__A1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__0544__A1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__0544__B1 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__0545__A1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__0545__A2 (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 ANTENNA__0546__A1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__0546__B1 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__0547__A1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__0547__A2 (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 ANTENNA__0548__A1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__0548__B1 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__0549__A1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__0549__A2 (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 ANTENNA__0551__A1 (.DIODE(net1172));
 sky130_fd_sc_hd__diode_2 ANTENNA__0553__A_N (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA__0553__B (.DIODE(_0191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0554__B (.DIODE(_0193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0555__B (.DIODE(_0193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0556__A (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__0556__B (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA__0557__A (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__0558__A (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__0559__B (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__0560__A2 (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__0561__B (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__0562__A2 (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__0563__B (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__0564__A2 (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__0565__B (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__0566__A2 (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__0567__B (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__0568__A1 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA__0568__A2 (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__0569__B (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__0570__A1 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA__0570__A2 (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__0571__B (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__0572__A2 (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__0573__B (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__0574__A2 (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__0575__B (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__0576__A2 (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__0577__B (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__0578__A2 (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__0579__B (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__0580__A2 (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__0581__B (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__0582__A2 (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__0583__B (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__0584__A2 (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__0585__B (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__0586__A2 (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__0587__B (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__0588__A2 (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__0589__B (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__0590__A2 (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__0591__B (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__0592__A2 (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__0593__B (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__0594__A1 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA__0594__A2 (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__0595__B (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__0596__A2 (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__0596__C1 (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 ANTENNA__0597__B (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__0598__A1 (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA__0598__A2 (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__0598__C1 (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 ANTENNA__0599__B (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__0600__A2 (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__0600__C1 (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 ANTENNA__0602__C1 (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 ANTENNA__0603__B (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__0604__A2 (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__0604__C1 (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 ANTENNA__0605__B (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__0606__A2 (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__0607__B (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__0608__A2 (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__0609__B (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__0610__A2 (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__0611__B (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__0612__A2 (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__0612__C1 (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 ANTENNA__0613__B (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__0614__A2 (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__0615__B (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__0616__A2 (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__0617__B (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__0618__A2 (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__0619__B (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__0620__A2 (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__0621__B (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA__0622__A2 (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__0622__C1 (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA__0624__B (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA__0625__C (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA__0626__A1 (.DIODE(net580));
 sky130_fd_sc_hd__diode_2 ANTENNA__0626__C1 (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 ANTENNA__0627__C (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA__0628__A1 (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA__0628__C1 (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 ANTENNA__0629__C (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA__0630__C1 (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 ANTENNA__0631__C (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA__0632__C1 (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 ANTENNA__0634__B (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA__0637__A1 (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA__0637__A2 (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA__0638__B (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA__0641__A1 (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA__0641__A2 (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA__0642__A (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA__0642__B (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA__0645__A1 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA__0645__A2 (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA__0646__A (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA__0646__B (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA__0649__A1 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA__0649__A2 (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA__0650__B (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA__0653__A1 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA__0653__A2 (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA__0654__B (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA__0657__A1 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA__0657__A2 (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA__0660__A1 (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA__0660__A2 (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA__0663__A1 (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA__0663__A2 (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA__0664__B (.DIODE(_0193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0665__C1 (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA__0666__A1 (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA__0667__A (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__0668__C1 (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA__0669__A1 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA__0670__A (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__0671__C1 (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA__0672__A1 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA__0673__A (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__0674__C1 (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA__0675__A2 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__0676__A (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__0677__C1 (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA__0678__A1 (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA__0679__A (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__0680__C1 (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA__0681__A1 (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA__0682__A (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__0683__C1 (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA__0684__A1 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA__0685__A (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__0686__C1 (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA__0687__A1 (.DIODE(net766));
 sky130_fd_sc_hd__diode_2 ANTENNA__0688__A (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__0689__A2 (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__0689__C1 (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA__0690__A1 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA__0691__A (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__0692__A2 (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__0692__C1 (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA__0693__A1 (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA__0693__A2 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__0694__A (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__0695__A2 (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__0695__C1 (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA__0696__A1 (.DIODE(net748));
 sky130_fd_sc_hd__diode_2 ANTENNA__0696__A2 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__0697__A (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__0698__A2 (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__0698__C1 (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA__0699__A1 (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA__0699__A2 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__0700__A (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__0701__A2 (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__0702__A1 (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA__0702__A2 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__0703__A (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__0704__A2 (.DIODE(net1081));
 sky130_fd_sc_hd__diode_2 ANTENNA__0705__A1 (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA__0706__A (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__0707__A2 (.DIODE(net1081));
 sky130_fd_sc_hd__diode_2 ANTENNA__0708__A1 (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA__0708__A2 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__0709__A (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__0710__A2 (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__0711__A1 (.DIODE(net742));
 sky130_fd_sc_hd__diode_2 ANTENNA__0711__A2 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__0712__A (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__0713__A2 (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__0714__A1 (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA__0714__A2 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__0715__A (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__0716__A2 (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__0716__C1 (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA__0717__A1 (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA__0717__A2 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__0718__A (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__0719__A2 (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__0719__B1 (.DIODE(_0237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0720__A1 (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA__0720__A2 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__0721__A (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__0722__A2 (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__0722__B1 (.DIODE(_0237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0723__A1 (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA__0723__A2 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__0724__A (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__0725__A2 (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__0726__A1 (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA__0726__A2 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__0727__A (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__0728__A2 (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__0728__C1 (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA__0729__A1 (.DIODE(net745));
 sky130_fd_sc_hd__diode_2 ANTENNA__0729__A2 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__0730__A (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__0731__A2 (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__0731__C1 (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA__0732__A1 (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA__0732__A2 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__0733__A (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__0734__A2 (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__0734__C1 (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA__0735__A1 (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA__0735__A2 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__0736__A (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__0740__B (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__0741__A2 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__0744__B1 (.DIODE(_0309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0745__A2 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__0747__B (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__0748__A1 (.DIODE(_0309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0751__B1 (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__0752__A2 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__0752__C1 (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA__0754__A (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__0755__A1 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA__0755__A2 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__0758__B1 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__0759__A1 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA__0759__A2 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__0762__B1 (.DIODE(_0309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0763__A2 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__0767__B1 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__0768__A2 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__0771__B1 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__0772__A2 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__0775__B1 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__0776__A2 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__0778__A (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__0779__A2 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__0783__B1 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__0784__A2 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__0787__B1 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__0788__A2 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__0791__B1 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__0792__A2 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__0795__B1 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__0796__A2 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__0800__B1 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__0801__A2 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__0803__A (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__0804__A2 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__0808__B1 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__0809__A1 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA__0809__A2 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__0812__B1 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__0813__A2 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__0813__C1 (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 ANTENNA__0816__C1 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__0817__A1 (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA__0817__A2 (.DIODE(_0309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0818__A (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__0821__A (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__0822__A2 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__0822__C1 (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 ANTENNA__0825__B1 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__0826__A2 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__0826__C1 (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 ANTENNA__0829__B1 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__0830__A2 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__0830__C1 (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 ANTENNA__0833__B1 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__0834__A2 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__0837__B1 (.DIODE(_0309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0838__A2 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__0839__A (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__0840__B (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__0841__A1 (.DIODE(_0309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0841__C1 (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA__0842__B (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__0843__A2 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__0844__B1 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__0845__A2 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__0847__B (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__0848__A1 (.DIODE(_0309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0851__B1 (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__0852__A2 (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__0855__B (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__0856__A1 (.DIODE(_0309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0858__B (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__0859__A1 (.DIODE(_0309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0862__B (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__0863__A1 (.DIODE(_0309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0863__C1 (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA__0864__C (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA__0865__C1 (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 ANTENNA__0867__A (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__0979__D (.DIODE(net507));
 sky130_fd_sc_hd__diode_2 ANTENNA__0982__D (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA__0983__D (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA__0984__D (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA__0985__D (.DIODE(net529));
 sky130_fd_sc_hd__diode_2 ANTENNA__0986__D (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA__0987__D (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA__1007__D (.DIODE(net487));
 sky130_fd_sc_hd__diode_2 ANTENNA__1013__A (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA__1014__A (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA__1015__A (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__1016__A (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__1017__A (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__1018__A (.DIODE(net582));
 sky130_fd_sc_hd__diode_2 ANTENNA__1019__A (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__1020__A (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__1021__A (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__1022__A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__1023__A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__1024__A (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__1025__A (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__1026__A (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__1027__A (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__1028__A (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__1029__A (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__1030__A (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__1031__A (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__1032__A (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__1033__A (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__1034__A (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__1035__A (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__1036__A (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__1037__A (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__1038__A (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__1039__A (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__1040__A (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__1041__A (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__1042__A (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__1043__A (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__1044__A (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__1045__A (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__1046__A (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA__1047__A (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__1048__A (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__1049__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout437_A (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout438_A (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout439_A (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout441_A (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout443_A (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout447_A (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout452_A (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout453_A (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout454_A (.DIODE(net565));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout455_A (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout456_A (.DIODE(net565));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout457_A (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout458_A (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout459_A (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout460_A (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout461_A (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout462_A (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout463_A (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout464_A (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout466_A (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout467_A (.DIODE(_0237_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout468_A (.DIODE(_0237_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout469_A (.DIODE(net1081));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout470_A (.DIODE(net1081));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout471_A (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout472_A (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout473_A (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout474_A (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout475_A (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold101_A (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold145_A (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold154_A (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold157_A (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold164_A (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold187_A (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold206_A (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold211_A (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold216_A (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold236_A (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold244_A (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold24_A (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold26_A (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold28_A (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold30_A (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold312_A (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold32_A (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold336_A (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold36_A (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold394_A (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold398_A (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold40_A (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold548_A (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold559_A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold572_A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold575_A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold578_A (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold581_A (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold584_A (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold591_A (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold594_A (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold600_A (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold603_A (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold606_A (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold609_A (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold612_A (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold614_A (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold618_A (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold621_A (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold624_A (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold627_A (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold630_A (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold634_A (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold689_A (.DIODE(_0191_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold690_A (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold78_A (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold82_A (.DIODE(_0117_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold83_A (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold85_A (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold89_A (.DIODE(_0114_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold90_A (.DIODE(_0116_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold91_A (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold92_A (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold97_A (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold98_A (.DIODE(_0115_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold99_A (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_output258_A (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA_output259_A (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_output260_A (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_output261_A (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_output262_A (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_output263_A (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_output264_A (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_output265_A (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_output266_A (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_output267_A (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA_output268_A (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_output269_A (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA_output270_A (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_output271_A (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_output272_A (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA_output273_A (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_output274_A (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA_output275_A (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA_output276_A (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA_output277_A (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA_output278_A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA_output279_A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA_output280_A (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA_output281_A (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA_output282_A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_output283_A (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_output284_A (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_output285_A (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_output286_A (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA_output287_A (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA_output288_A (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA_output289_A (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA_output290_A (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA_output291_A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_output292_A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA_output293_A (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_output294_A (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA_output295_A (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA_output296_A (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_output297_A (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA_output298_A (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_output299_A (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA_output300_A (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_output301_A (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA_output302_A (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_output303_A (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA_output304_A (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA_output305_A (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA_output306_A (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA_output307_A (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_output308_A (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA_output309_A (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA_output310_A (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA_output311_A (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_output312_A (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_output313_A (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA_output314_A (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_output315_A (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_output316_A (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA_output317_A (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_output318_A (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA_output319_A (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_output320_A (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA_output321_A (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_output322_A (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_output323_A (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_output324_A (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_output325_A (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA_output326_A (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_output327_A (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_output328_A (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA_output329_A (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA_output330_A (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_output331_A (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA_output332_A (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA_output333_A (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA_output334_A (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_output335_A (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA_output336_A (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA_output337_A (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA_output338_A (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA_output339_A (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_output340_A (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_output341_A (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_output342_A (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_output343_A (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_output344_A (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA_output345_A (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_output346_A (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_output347_A (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA_output348_A (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA_output349_A (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA_output350_A (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA_output351_A (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA_output352_A (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA_output353_A (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA_output354_A (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA_output355_A (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA_output356_A (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA_output357_A (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA_output358_A (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA_output359_A (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA_output360_A (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA_output361_A (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA_output362_A (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_output363_A (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA_output364_A (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA_output365_A (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_output366_A (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA_output367_A (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA_output368_A (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA_output369_A (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA_output370_A (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA_output371_A (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA_output372_A (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA_output374_A (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA_output375_A (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA_output376_A (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA_output377_A (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_output378_A (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_output379_A (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA_output380_A (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA_output381_A (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA_output382_A (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA_output383_A (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA_output385_A (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA_output386_A (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_output387_A (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA_output388_A (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_output389_A (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA_output390_A (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA_output391_A (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA_output392_A (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_output393_A (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA_output396_A (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA_output397_A (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA_output398_A (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA_output399_A (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA_output400_A (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA_output401_A (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA_output402_A (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_output404_A (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_output405_A (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_output406_A (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA_output408_A (.DIODE(net754));
 sky130_fd_sc_hd__diode_2 ANTENNA_output409_A (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_output410_A (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_output411_A (.DIODE(net766));
 sky130_fd_sc_hd__diode_2 ANTENNA_output412_A (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_output413_A (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA_output414_A (.DIODE(net748));
 sky130_fd_sc_hd__diode_2 ANTENNA_output415_A (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_output416_A (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_output417_A (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_output418_A (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_output419_A (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_output420_A (.DIODE(net742));
 sky130_fd_sc_hd__diode_2 ANTENNA_output421_A (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_output422_A (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA_output423_A (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_output424_A (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA_output425_A (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_output426_A (.DIODE(net745));
 sky130_fd_sc_hd__diode_2 ANTENNA_output427_A (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA_output428_A (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_output429_A (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_output430_A (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_output431_A (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_output432_A (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_output433_A (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_output434_A (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA_output435_A (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_output436_A (.DIODE(net787));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_86 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_6 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_198_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_199_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_200_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_201_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_201_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_204_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_205_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_205_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_206_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_206_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_207_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_207_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_208_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_208_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_209_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_210_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_210_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_210_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_214_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_215_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_215_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_216_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_216_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_216_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_218_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_218_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_218_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_218_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_218_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_218_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_218_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_218_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_218_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_220_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_220_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_220_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_220_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_220_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_220_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_220_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_220_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_220_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_221_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_221_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_221_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_221_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_221_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_221_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_221_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_221_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_222_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_222_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_223_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_223_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_223_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_224_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_224_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_224_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_224_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_224_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_225_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_225_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_226_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_226_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_226_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_226_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_226_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_227_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_227_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_227_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_227_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_227_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_228_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_228_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_229_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_230_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_230_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_231_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_231_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_231_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_231_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_232_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_232_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_233_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_233_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_233_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_233_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_233_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_234_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_234_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_235_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_235_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_235_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_235_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_235_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_236_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_236_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_236_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_237_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_237_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_237_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_237_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_238_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_239_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_239_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_239_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_239_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_239_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_239_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_240_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_240_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_240_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_240_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_241_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_241_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_241_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_241_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_241_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_242_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_242_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_242_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_242_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_243_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_243_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_243_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_243_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_243_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_244_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_244_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_244_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_244_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_244_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_245_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_245_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_245_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_245_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_245_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_246_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_246_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_246_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_246_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_247_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_247_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_247_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_247_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_247_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_247_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_248_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_248_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_248_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_249_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_249_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_249_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_249_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_249_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_250_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_250_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_250_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_250_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_250_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_250_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_251_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_251_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_251_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_252_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_252_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_252_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_252_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_253_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_253_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_253_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_253_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_253_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_253_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_253_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_254_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_254_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_254_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_254_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_255_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_255_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_255_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_255_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_255_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_255_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_256_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_256_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_256_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_256_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_256_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_256_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_256_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_257_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_257_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_257_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_257_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_257_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_258_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_258_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_258_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_258_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_258_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_259_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_259_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_259_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_259_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_259_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_259_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_259_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_260_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_260_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_260_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_260_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_260_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_260_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_260_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_261_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_261_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_261_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_261_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_261_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_261_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_262_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_262_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_262_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_262_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_263_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_263_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_263_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_263_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_264_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_264_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_264_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_264_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_264_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_265_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_265_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_265_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_265_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_265_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_266_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_266_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_266_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_267_16 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_267_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_267_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_267_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_267_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_268_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_268_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_268_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_268_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_268_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_269_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_269_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_270_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_270_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_270_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_270_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_270_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_271_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_271_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_271_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_271_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_271_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_271_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_272_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_273_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_273_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_273_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_273_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_273_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_273_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_274_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_274_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_274_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_274_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_274_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_274_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_274_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_275_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_275_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_275_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_275_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_275_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_276_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_276_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_276_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_276_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_276_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_277_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_277_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_277_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_277_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_277_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_277_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_278_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_278_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_278_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_279_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_279_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_279_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_279_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_279_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_280_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_280_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_280_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_280_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_280_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_281_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_281_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_281_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_281_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_281_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_282_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_282_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_282_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_282_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_283_16 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_283_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_283_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_284_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_284_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_284_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_285_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_285_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_285_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_285_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_285_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_285_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_285_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_285_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_285_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_285_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_285_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_285_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_285_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_285_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_285_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_285_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_285_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_286_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_286_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_286_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_286_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_286_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_286_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_286_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_286_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_286_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_286_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_286_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_286_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_286_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_286_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_286_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_286_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_286_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_286_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_286_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_286_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_287_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_287_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_287_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_287_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_287_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_287_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_287_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_287_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_287_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_287_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_287_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_287_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_287_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_287_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_287_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_287_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_287_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_287_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_287_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_287_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_288_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_288_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_288_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_288_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_288_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_288_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_288_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_288_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_288_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_288_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_288_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_288_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_288_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_288_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_288_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_288_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_288_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_289_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_289_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_289_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_289_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_289_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_289_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_289_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_289_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_289_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_289_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_289_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_289_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_289_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_289_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_289_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_289_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_290_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_290_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_290_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_290_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_290_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_290_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_290_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_290_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_290_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_290_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_290_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_290_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_290_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_290_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_291_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_291_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_291_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_291_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_291_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_291_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_291_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_291_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_291_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_291_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_291_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_291_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_291_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_291_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_291_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_292_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_292_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_292_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_292_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_292_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_292_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_292_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_292_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_292_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_292_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_292_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_292_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_292_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_292_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_293_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_293_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_293_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_293_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_293_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_293_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_293_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_293_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_293_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_293_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_293_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_293_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_293_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_293_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_294_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_294_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_294_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_294_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_294_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_294_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_294_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_294_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_294_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_294_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_294_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_294_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_294_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_294_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_295_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_295_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_295_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_295_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_295_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_295_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_295_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_295_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_295_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_295_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_295_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_295_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_295_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_295_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_295_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_296_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_296_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_296_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_296_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_296_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_296_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_296_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_296_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_296_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_296_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_296_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_296_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_296_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_296_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_297_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_297_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_297_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_297_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_297_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_297_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_297_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_297_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_297_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_297_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_297_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_297_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_297_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_297_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_297_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_298_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_298_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_298_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_298_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_298_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_298_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_298_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_298_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_298_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_298_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_298_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_298_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_298_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_298_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_299_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_299_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_299_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_299_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_299_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_299_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_299_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_300_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_300_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_300_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_300_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_300_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_300_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_300_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_300_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_300_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_300_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_300_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_300_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_300_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_300_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_301_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_301_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_301_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_301_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_301_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_301_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_301_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_301_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_301_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_301_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_301_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_301_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_301_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_301_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_301_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_302_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_302_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_302_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_302_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_302_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_302_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_302_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_302_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_302_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_302_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_302_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_302_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_302_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_302_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_303_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_303_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_303_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_303_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_303_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_303_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_303_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_303_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_303_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_303_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_303_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_303_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_303_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_303_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_303_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_304_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_304_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_304_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_304_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_304_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_304_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_304_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_304_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_304_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_304_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_304_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_304_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_304_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_304_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_305_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_305_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_305_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_305_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_305_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_305_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_305_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_305_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_305_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_305_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_305_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_305_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_305_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_305_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_306_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_306_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_306_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_306_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_306_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_306_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_306_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_306_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_306_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_306_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_306_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_306_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_306_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_306_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_307_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_307_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_307_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_307_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_307_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_307_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_307_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_307_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_308_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_308_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_308_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_308_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_308_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_308_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_308_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_308_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_308_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_308_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_308_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_308_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_308_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_308_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_309_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_309_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_309_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_309_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_309_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_309_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_309_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_309_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_309_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_309_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_309_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_309_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_309_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_309_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_309_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_310_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_310_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_310_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_310_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_310_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_310_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_310_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_310_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_310_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_310_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_310_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_310_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_310_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_310_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_311_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_311_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_311_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_311_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_311_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_311_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_311_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_311_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_311_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_311_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_311_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_311_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_311_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_311_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_312_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_312_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_312_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_312_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_312_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_312_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_312_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_312_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_312_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_312_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_312_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_312_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_312_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_312_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_313_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_313_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_313_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_313_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_313_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_313_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_313_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_313_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_313_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_313_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_313_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_313_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_313_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_313_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_313_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_314_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_314_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_314_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_314_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_314_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_314_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_314_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_314_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_314_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_314_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_314_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_314_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_314_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_314_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_315_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_315_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_315_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_315_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_315_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_315_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_315_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_315_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_315_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_315_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_315_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_315_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_315_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_315_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_315_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_316_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_316_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_316_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_316_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_316_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_316_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_316_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_316_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_316_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_316_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_316_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_316_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_316_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_316_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_317_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_317_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_317_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_317_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_317_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_317_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_317_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_317_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_317_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_317_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_317_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_317_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_317_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_317_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_318_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_318_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_318_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_318_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_318_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_318_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_318_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_318_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_318_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_318_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_318_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_318_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_318_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_318_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_319_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_319_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_319_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_319_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_319_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_319_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_319_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_319_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_319_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_319_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_319_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_319_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_319_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_319_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_319_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_320_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_320_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_320_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_320_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_320_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_320_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_320_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_320_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_320_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_320_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_320_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_320_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_320_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_320_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_321_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_321_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_321_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_321_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_321_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_321_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_321_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_321_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_321_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_321_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_321_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_321_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_321_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_321_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_321_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_322_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_322_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_322_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_322_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_322_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_322_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_322_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_322_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_322_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_322_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_322_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_322_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_322_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_322_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_322_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_323_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_323_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_323_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_323_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_323_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_323_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_323_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_323_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_323_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_323_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_323_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_323_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_323_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_323_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_324_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_324_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_324_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_324_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_324_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_324_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_324_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_324_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_324_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_324_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_324_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_324_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_324_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_324_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_324_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_325_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_325_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_325_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_325_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_325_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_325_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_325_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_325_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_325_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_325_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_325_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_325_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_325_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_325_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_325_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_325_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_326_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_326_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_326_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_326_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_326_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_326_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_326_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_326_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_326_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_326_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_326_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_326_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_326_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_326_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_326_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_327_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_327_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_327_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_327_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_327_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_327_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_327_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_327_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_327_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_327_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_327_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_327_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_327_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_327_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_327_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_327_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_328_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_328_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_328_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_328_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_328_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_328_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_328_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_328_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_328_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_328_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_328_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_328_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_328_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_328_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_328_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_329_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_329_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_329_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_329_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_329_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_329_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_329_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_329_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_329_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_329_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_329_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_329_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_329_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_329_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_329_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_330_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_330_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_330_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_330_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_330_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_330_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_330_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_330_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_330_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_330_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_330_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_330_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_330_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_330_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_330_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_331_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_331_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_331_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_331_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_331_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_331_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_331_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_331_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_331_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_331_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_331_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_331_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_331_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_331_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_331_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_331_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_332_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_332_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_332_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_332_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_332_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_332_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_332_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_332_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_332_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_332_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_332_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_332_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_332_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_332_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_332_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_333_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_333_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_333_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_333_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_333_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_333_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_333_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_333_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_333_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_333_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_333_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_333_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_333_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_333_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_333_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_333_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_334_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_334_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_334_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_334_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_334_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_334_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_334_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_334_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_334_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_334_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_334_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_334_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_334_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_334_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_334_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_335_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_335_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_335_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_335_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_335_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_335_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_335_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_335_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_335_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_335_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_335_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_335_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_335_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_335_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_335_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_336_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_336_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_336_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_336_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_336_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_336_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_336_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_336_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_336_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_336_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_336_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_336_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_336_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_336_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_336_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_337_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_337_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_337_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_337_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_337_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_337_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_337_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_337_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_337_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_337_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_337_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_337_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_337_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_337_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_337_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_338_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_338_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_338_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_338_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_338_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_338_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_338_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_338_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_338_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_338_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_338_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_338_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_338_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_338_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_338_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_339_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_339_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_339_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_339_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_339_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_339_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_339_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_339_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_339_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_339_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_339_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_339_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_339_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_339_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_339_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_339_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_340_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_340_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_340_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_340_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_340_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_340_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_340_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_340_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_340_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_340_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_340_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_340_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_340_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_340_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_340_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_341_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_341_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_341_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_341_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_341_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_341_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_341_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_341_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_341_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_341_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_341_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_341_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_341_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_341_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_341_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_342_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_342_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_342_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_342_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_342_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_342_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_342_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_342_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_342_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_342_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_342_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_342_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_342_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_342_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_343_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_343_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_343_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_343_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_343_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_343_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_343_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_343_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_343_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_343_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_343_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_343_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_343_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_343_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_343_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_344_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_344_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_344_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_344_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_344_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_344_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_344_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_344_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_344_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_344_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_344_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_344_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_344_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_344_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_345_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_345_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_345_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_345_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_345_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_345_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_345_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_345_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_345_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_345_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_345_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_345_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_345_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_345_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_345_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_346_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_346_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_346_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_346_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_346_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_346_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_346_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_346_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_346_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_346_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_346_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_346_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_346_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_346_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_346_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_347_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_347_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_347_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_347_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_347_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_347_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_347_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_347_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_347_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_347_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_347_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_347_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_347_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_347_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_347_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_348_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_348_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_348_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_348_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_348_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_348_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_348_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_348_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_348_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_348_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_348_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_348_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_348_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_348_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_348_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_349_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_349_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_349_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_349_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_349_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_349_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_349_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_349_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_349_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_349_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_349_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_349_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_349_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_349_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_350_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_350_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_350_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_350_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_350_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_350_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_350_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_350_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_350_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_350_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_350_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_350_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_350_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_350_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_350_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_351_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_351_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_351_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_351_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_351_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_351_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_351_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_351_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_351_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_351_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_351_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_351_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_351_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_351_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_351_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_352_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_352_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_352_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_352_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_352_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_352_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_352_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_352_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_352_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_352_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_352_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_352_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_352_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_352_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_353_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_353_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_353_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_353_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_353_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_353_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_353_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_353_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_353_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_353_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_353_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_353_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_353_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_353_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_353_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_354_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_354_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_354_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_354_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_354_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_354_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_354_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_354_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_354_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_354_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_354_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_354_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_354_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_354_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_354_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_355_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_355_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_355_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_355_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_355_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_355_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_355_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_355_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_355_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_355_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_355_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_355_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_355_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_355_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_355_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_356_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_356_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_356_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_356_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_356_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_356_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_356_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_356_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_356_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_356_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_356_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_356_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_356_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_356_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_356_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_356_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_357_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_357_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_357_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_357_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_357_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_357_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_357_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_357_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_357_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_357_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_357_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_357_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_357_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_357_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_357_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_357_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_357_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_357_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_357_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_358_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_358_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_358_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_358_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_358_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_358_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_358_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_358_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_358_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_358_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_358_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_358_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_358_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_358_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_358_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_358_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_358_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_358_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_358_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_358_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_358_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_358_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_358_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_358_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_358_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_358_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_358_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_358_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_358_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_358_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_358_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_358_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_358_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_358_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_358_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_358_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_358_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_358_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_358_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_358_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_358_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_358_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_358_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_358_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_358_36 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_358_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_358_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_358_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_358_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_358_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_358_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_358_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_358_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_358_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_358_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_358_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_358_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_358_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_186 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_348 ();
 sky130_fd_sc_hd__decap_3 PHY_349 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_350 ();
 sky130_fd_sc_hd__decap_3 PHY_351 ();
 sky130_fd_sc_hd__decap_3 PHY_352 ();
 sky130_fd_sc_hd__decap_3 PHY_353 ();
 sky130_fd_sc_hd__decap_3 PHY_354 ();
 sky130_fd_sc_hd__decap_3 PHY_355 ();
 sky130_fd_sc_hd__decap_3 PHY_356 ();
 sky130_fd_sc_hd__decap_3 PHY_357 ();
 sky130_fd_sc_hd__decap_3 PHY_358 ();
 sky130_fd_sc_hd__decap_3 PHY_359 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_360 ();
 sky130_fd_sc_hd__decap_3 PHY_361 ();
 sky130_fd_sc_hd__decap_3 PHY_362 ();
 sky130_fd_sc_hd__decap_3 PHY_363 ();
 sky130_fd_sc_hd__decap_3 PHY_364 ();
 sky130_fd_sc_hd__decap_3 PHY_365 ();
 sky130_fd_sc_hd__decap_3 PHY_366 ();
 sky130_fd_sc_hd__decap_3 PHY_367 ();
 sky130_fd_sc_hd__decap_3 PHY_368 ();
 sky130_fd_sc_hd__decap_3 PHY_369 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_370 ();
 sky130_fd_sc_hd__decap_3 PHY_371 ();
 sky130_fd_sc_hd__decap_3 PHY_372 ();
 sky130_fd_sc_hd__decap_3 PHY_373 ();
 sky130_fd_sc_hd__decap_3 PHY_374 ();
 sky130_fd_sc_hd__decap_3 PHY_375 ();
 sky130_fd_sc_hd__decap_3 PHY_376 ();
 sky130_fd_sc_hd__decap_3 PHY_377 ();
 sky130_fd_sc_hd__decap_3 PHY_378 ();
 sky130_fd_sc_hd__decap_3 PHY_379 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_380 ();
 sky130_fd_sc_hd__decap_3 PHY_381 ();
 sky130_fd_sc_hd__decap_3 PHY_382 ();
 sky130_fd_sc_hd__decap_3 PHY_383 ();
 sky130_fd_sc_hd__decap_3 PHY_384 ();
 sky130_fd_sc_hd__decap_3 PHY_385 ();
 sky130_fd_sc_hd__decap_3 PHY_386 ();
 sky130_fd_sc_hd__decap_3 PHY_387 ();
 sky130_fd_sc_hd__decap_3 PHY_388 ();
 sky130_fd_sc_hd__decap_3 PHY_389 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_390 ();
 sky130_fd_sc_hd__decap_3 PHY_391 ();
 sky130_fd_sc_hd__decap_3 PHY_392 ();
 sky130_fd_sc_hd__decap_3 PHY_393 ();
 sky130_fd_sc_hd__decap_3 PHY_394 ();
 sky130_fd_sc_hd__decap_3 PHY_395 ();
 sky130_fd_sc_hd__decap_3 PHY_396 ();
 sky130_fd_sc_hd__decap_3 PHY_397 ();
 sky130_fd_sc_hd__decap_3 PHY_398 ();
 sky130_fd_sc_hd__decap_3 PHY_399 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_400 ();
 sky130_fd_sc_hd__decap_3 PHY_401 ();
 sky130_fd_sc_hd__decap_3 PHY_402 ();
 sky130_fd_sc_hd__decap_3 PHY_403 ();
 sky130_fd_sc_hd__decap_3 PHY_404 ();
 sky130_fd_sc_hd__decap_3 PHY_405 ();
 sky130_fd_sc_hd__decap_3 PHY_406 ();
 sky130_fd_sc_hd__decap_3 PHY_407 ();
 sky130_fd_sc_hd__decap_3 PHY_408 ();
 sky130_fd_sc_hd__decap_3 PHY_409 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_410 ();
 sky130_fd_sc_hd__decap_3 PHY_411 ();
 sky130_fd_sc_hd__decap_3 PHY_412 ();
 sky130_fd_sc_hd__decap_3 PHY_413 ();
 sky130_fd_sc_hd__decap_3 PHY_414 ();
 sky130_fd_sc_hd__decap_3 PHY_415 ();
 sky130_fd_sc_hd__decap_3 PHY_416 ();
 sky130_fd_sc_hd__decap_3 PHY_417 ();
 sky130_fd_sc_hd__decap_3 PHY_418 ();
 sky130_fd_sc_hd__decap_3 PHY_419 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_420 ();
 sky130_fd_sc_hd__decap_3 PHY_421 ();
 sky130_fd_sc_hd__decap_3 PHY_422 ();
 sky130_fd_sc_hd__decap_3 PHY_423 ();
 sky130_fd_sc_hd__decap_3 PHY_424 ();
 sky130_fd_sc_hd__decap_3 PHY_425 ();
 sky130_fd_sc_hd__decap_3 PHY_426 ();
 sky130_fd_sc_hd__decap_3 PHY_427 ();
 sky130_fd_sc_hd__decap_3 PHY_428 ();
 sky130_fd_sc_hd__decap_3 PHY_429 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_430 ();
 sky130_fd_sc_hd__decap_3 PHY_431 ();
 sky130_fd_sc_hd__decap_3 PHY_432 ();
 sky130_fd_sc_hd__decap_3 PHY_433 ();
 sky130_fd_sc_hd__decap_3 PHY_434 ();
 sky130_fd_sc_hd__decap_3 PHY_435 ();
 sky130_fd_sc_hd__decap_3 PHY_436 ();
 sky130_fd_sc_hd__decap_3 PHY_437 ();
 sky130_fd_sc_hd__decap_3 PHY_438 ();
 sky130_fd_sc_hd__decap_3 PHY_439 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_440 ();
 sky130_fd_sc_hd__decap_3 PHY_441 ();
 sky130_fd_sc_hd__decap_3 PHY_442 ();
 sky130_fd_sc_hd__decap_3 PHY_443 ();
 sky130_fd_sc_hd__decap_3 PHY_444 ();
 sky130_fd_sc_hd__decap_3 PHY_445 ();
 sky130_fd_sc_hd__decap_3 PHY_446 ();
 sky130_fd_sc_hd__decap_3 PHY_447 ();
 sky130_fd_sc_hd__decap_3 PHY_448 ();
 sky130_fd_sc_hd__decap_3 PHY_449 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_450 ();
 sky130_fd_sc_hd__decap_3 PHY_451 ();
 sky130_fd_sc_hd__decap_3 PHY_452 ();
 sky130_fd_sc_hd__decap_3 PHY_453 ();
 sky130_fd_sc_hd__decap_3 PHY_454 ();
 sky130_fd_sc_hd__decap_3 PHY_455 ();
 sky130_fd_sc_hd__decap_3 PHY_456 ();
 sky130_fd_sc_hd__decap_3 PHY_457 ();
 sky130_fd_sc_hd__decap_3 PHY_458 ();
 sky130_fd_sc_hd__decap_3 PHY_459 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_460 ();
 sky130_fd_sc_hd__decap_3 PHY_461 ();
 sky130_fd_sc_hd__decap_3 PHY_462 ();
 sky130_fd_sc_hd__decap_3 PHY_463 ();
 sky130_fd_sc_hd__decap_3 PHY_464 ();
 sky130_fd_sc_hd__decap_3 PHY_465 ();
 sky130_fd_sc_hd__decap_3 PHY_466 ();
 sky130_fd_sc_hd__decap_3 PHY_467 ();
 sky130_fd_sc_hd__decap_3 PHY_468 ();
 sky130_fd_sc_hd__decap_3 PHY_469 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_470 ();
 sky130_fd_sc_hd__decap_3 PHY_471 ();
 sky130_fd_sc_hd__decap_3 PHY_472 ();
 sky130_fd_sc_hd__decap_3 PHY_473 ();
 sky130_fd_sc_hd__decap_3 PHY_474 ();
 sky130_fd_sc_hd__decap_3 PHY_475 ();
 sky130_fd_sc_hd__decap_3 PHY_476 ();
 sky130_fd_sc_hd__decap_3 PHY_477 ();
 sky130_fd_sc_hd__decap_3 PHY_478 ();
 sky130_fd_sc_hd__decap_3 PHY_479 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_480 ();
 sky130_fd_sc_hd__decap_3 PHY_481 ();
 sky130_fd_sc_hd__decap_3 PHY_482 ();
 sky130_fd_sc_hd__decap_3 PHY_483 ();
 sky130_fd_sc_hd__decap_3 PHY_484 ();
 sky130_fd_sc_hd__decap_3 PHY_485 ();
 sky130_fd_sc_hd__decap_3 PHY_486 ();
 sky130_fd_sc_hd__decap_3 PHY_487 ();
 sky130_fd_sc_hd__decap_3 PHY_488 ();
 sky130_fd_sc_hd__decap_3 PHY_489 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_490 ();
 sky130_fd_sc_hd__decap_3 PHY_491 ();
 sky130_fd_sc_hd__decap_3 PHY_492 ();
 sky130_fd_sc_hd__decap_3 PHY_493 ();
 sky130_fd_sc_hd__decap_3 PHY_494 ();
 sky130_fd_sc_hd__decap_3 PHY_495 ();
 sky130_fd_sc_hd__decap_3 PHY_496 ();
 sky130_fd_sc_hd__decap_3 PHY_497 ();
 sky130_fd_sc_hd__decap_3 PHY_498 ();
 sky130_fd_sc_hd__decap_3 PHY_499 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_500 ();
 sky130_fd_sc_hd__decap_3 PHY_501 ();
 sky130_fd_sc_hd__decap_3 PHY_502 ();
 sky130_fd_sc_hd__decap_3 PHY_503 ();
 sky130_fd_sc_hd__decap_3 PHY_504 ();
 sky130_fd_sc_hd__decap_3 PHY_505 ();
 sky130_fd_sc_hd__decap_3 PHY_506 ();
 sky130_fd_sc_hd__decap_3 PHY_507 ();
 sky130_fd_sc_hd__decap_3 PHY_508 ();
 sky130_fd_sc_hd__decap_3 PHY_509 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_510 ();
 sky130_fd_sc_hd__decap_3 PHY_511 ();
 sky130_fd_sc_hd__decap_3 PHY_512 ();
 sky130_fd_sc_hd__decap_3 PHY_513 ();
 sky130_fd_sc_hd__decap_3 PHY_514 ();
 sky130_fd_sc_hd__decap_3 PHY_515 ();
 sky130_fd_sc_hd__decap_3 PHY_516 ();
 sky130_fd_sc_hd__decap_3 PHY_517 ();
 sky130_fd_sc_hd__decap_3 PHY_518 ();
 sky130_fd_sc_hd__decap_3 PHY_519 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_520 ();
 sky130_fd_sc_hd__decap_3 PHY_521 ();
 sky130_fd_sc_hd__decap_3 PHY_522 ();
 sky130_fd_sc_hd__decap_3 PHY_523 ();
 sky130_fd_sc_hd__decap_3 PHY_524 ();
 sky130_fd_sc_hd__decap_3 PHY_525 ();
 sky130_fd_sc_hd__decap_3 PHY_526 ();
 sky130_fd_sc_hd__decap_3 PHY_527 ();
 sky130_fd_sc_hd__decap_3 PHY_528 ();
 sky130_fd_sc_hd__decap_3 PHY_529 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_530 ();
 sky130_fd_sc_hd__decap_3 PHY_531 ();
 sky130_fd_sc_hd__decap_3 PHY_532 ();
 sky130_fd_sc_hd__decap_3 PHY_533 ();
 sky130_fd_sc_hd__decap_3 PHY_534 ();
 sky130_fd_sc_hd__decap_3 PHY_535 ();
 sky130_fd_sc_hd__decap_3 PHY_536 ();
 sky130_fd_sc_hd__decap_3 PHY_537 ();
 sky130_fd_sc_hd__decap_3 PHY_538 ();
 sky130_fd_sc_hd__decap_3 PHY_539 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_540 ();
 sky130_fd_sc_hd__decap_3 PHY_541 ();
 sky130_fd_sc_hd__decap_3 PHY_542 ();
 sky130_fd_sc_hd__decap_3 PHY_543 ();
 sky130_fd_sc_hd__decap_3 PHY_544 ();
 sky130_fd_sc_hd__decap_3 PHY_545 ();
 sky130_fd_sc_hd__decap_3 PHY_546 ();
 sky130_fd_sc_hd__decap_3 PHY_547 ();
 sky130_fd_sc_hd__decap_3 PHY_548 ();
 sky130_fd_sc_hd__decap_3 PHY_549 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_550 ();
 sky130_fd_sc_hd__decap_3 PHY_551 ();
 sky130_fd_sc_hd__decap_3 PHY_552 ();
 sky130_fd_sc_hd__decap_3 PHY_553 ();
 sky130_fd_sc_hd__decap_3 PHY_554 ();
 sky130_fd_sc_hd__decap_3 PHY_555 ();
 sky130_fd_sc_hd__decap_3 PHY_556 ();
 sky130_fd_sc_hd__decap_3 PHY_557 ();
 sky130_fd_sc_hd__decap_3 PHY_558 ();
 sky130_fd_sc_hd__decap_3 PHY_559 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_560 ();
 sky130_fd_sc_hd__decap_3 PHY_561 ();
 sky130_fd_sc_hd__decap_3 PHY_562 ();
 sky130_fd_sc_hd__decap_3 PHY_563 ();
 sky130_fd_sc_hd__decap_3 PHY_564 ();
 sky130_fd_sc_hd__decap_3 PHY_565 ();
 sky130_fd_sc_hd__decap_3 PHY_566 ();
 sky130_fd_sc_hd__decap_3 PHY_567 ();
 sky130_fd_sc_hd__decap_3 PHY_568 ();
 sky130_fd_sc_hd__decap_3 PHY_569 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_570 ();
 sky130_fd_sc_hd__decap_3 PHY_571 ();
 sky130_fd_sc_hd__decap_3 PHY_572 ();
 sky130_fd_sc_hd__decap_3 PHY_573 ();
 sky130_fd_sc_hd__decap_3 PHY_574 ();
 sky130_fd_sc_hd__decap_3 PHY_575 ();
 sky130_fd_sc_hd__decap_3 PHY_576 ();
 sky130_fd_sc_hd__decap_3 PHY_577 ();
 sky130_fd_sc_hd__decap_3 PHY_578 ();
 sky130_fd_sc_hd__decap_3 PHY_579 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_580 ();
 sky130_fd_sc_hd__decap_3 PHY_581 ();
 sky130_fd_sc_hd__decap_3 PHY_582 ();
 sky130_fd_sc_hd__decap_3 PHY_583 ();
 sky130_fd_sc_hd__decap_3 PHY_584 ();
 sky130_fd_sc_hd__decap_3 PHY_585 ();
 sky130_fd_sc_hd__decap_3 PHY_586 ();
 sky130_fd_sc_hd__decap_3 PHY_587 ();
 sky130_fd_sc_hd__decap_3 PHY_588 ();
 sky130_fd_sc_hd__decap_3 PHY_589 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_590 ();
 sky130_fd_sc_hd__decap_3 PHY_591 ();
 sky130_fd_sc_hd__decap_3 PHY_592 ();
 sky130_fd_sc_hd__decap_3 PHY_593 ();
 sky130_fd_sc_hd__decap_3 PHY_594 ();
 sky130_fd_sc_hd__decap_3 PHY_595 ();
 sky130_fd_sc_hd__decap_3 PHY_596 ();
 sky130_fd_sc_hd__decap_3 PHY_597 ();
 sky130_fd_sc_hd__decap_3 PHY_598 ();
 sky130_fd_sc_hd__decap_3 PHY_599 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_600 ();
 sky130_fd_sc_hd__decap_3 PHY_601 ();
 sky130_fd_sc_hd__decap_3 PHY_602 ();
 sky130_fd_sc_hd__decap_3 PHY_603 ();
 sky130_fd_sc_hd__decap_3 PHY_604 ();
 sky130_fd_sc_hd__decap_3 PHY_605 ();
 sky130_fd_sc_hd__decap_3 PHY_606 ();
 sky130_fd_sc_hd__decap_3 PHY_607 ();
 sky130_fd_sc_hd__decap_3 PHY_608 ();
 sky130_fd_sc_hd__decap_3 PHY_609 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_610 ();
 sky130_fd_sc_hd__decap_3 PHY_611 ();
 sky130_fd_sc_hd__decap_3 PHY_612 ();
 sky130_fd_sc_hd__decap_3 PHY_613 ();
 sky130_fd_sc_hd__decap_3 PHY_614 ();
 sky130_fd_sc_hd__decap_3 PHY_615 ();
 sky130_fd_sc_hd__decap_3 PHY_616 ();
 sky130_fd_sc_hd__decap_3 PHY_617 ();
 sky130_fd_sc_hd__decap_3 PHY_618 ();
 sky130_fd_sc_hd__decap_3 PHY_619 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_620 ();
 sky130_fd_sc_hd__decap_3 PHY_621 ();
 sky130_fd_sc_hd__decap_3 PHY_622 ();
 sky130_fd_sc_hd__decap_3 PHY_623 ();
 sky130_fd_sc_hd__decap_3 PHY_624 ();
 sky130_fd_sc_hd__decap_3 PHY_625 ();
 sky130_fd_sc_hd__decap_3 PHY_626 ();
 sky130_fd_sc_hd__decap_3 PHY_627 ();
 sky130_fd_sc_hd__decap_3 PHY_628 ();
 sky130_fd_sc_hd__decap_3 PHY_629 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_630 ();
 sky130_fd_sc_hd__decap_3 PHY_631 ();
 sky130_fd_sc_hd__decap_3 PHY_632 ();
 sky130_fd_sc_hd__decap_3 PHY_633 ();
 sky130_fd_sc_hd__decap_3 PHY_634 ();
 sky130_fd_sc_hd__decap_3 PHY_635 ();
 sky130_fd_sc_hd__decap_3 PHY_636 ();
 sky130_fd_sc_hd__decap_3 PHY_637 ();
 sky130_fd_sc_hd__decap_3 PHY_638 ();
 sky130_fd_sc_hd__decap_3 PHY_639 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_640 ();
 sky130_fd_sc_hd__decap_3 PHY_641 ();
 sky130_fd_sc_hd__decap_3 PHY_642 ();
 sky130_fd_sc_hd__decap_3 PHY_643 ();
 sky130_fd_sc_hd__decap_3 PHY_644 ();
 sky130_fd_sc_hd__decap_3 PHY_645 ();
 sky130_fd_sc_hd__decap_3 PHY_646 ();
 sky130_fd_sc_hd__decap_3 PHY_647 ();
 sky130_fd_sc_hd__decap_3 PHY_648 ();
 sky130_fd_sc_hd__decap_3 PHY_649 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_650 ();
 sky130_fd_sc_hd__decap_3 PHY_651 ();
 sky130_fd_sc_hd__decap_3 PHY_652 ();
 sky130_fd_sc_hd__decap_3 PHY_653 ();
 sky130_fd_sc_hd__decap_3 PHY_654 ();
 sky130_fd_sc_hd__decap_3 PHY_655 ();
 sky130_fd_sc_hd__decap_3 PHY_656 ();
 sky130_fd_sc_hd__decap_3 PHY_657 ();
 sky130_fd_sc_hd__decap_3 PHY_658 ();
 sky130_fd_sc_hd__decap_3 PHY_659 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_660 ();
 sky130_fd_sc_hd__decap_3 PHY_661 ();
 sky130_fd_sc_hd__decap_3 PHY_662 ();
 sky130_fd_sc_hd__decap_3 PHY_663 ();
 sky130_fd_sc_hd__decap_3 PHY_664 ();
 sky130_fd_sc_hd__decap_3 PHY_665 ();
 sky130_fd_sc_hd__decap_3 PHY_666 ();
 sky130_fd_sc_hd__decap_3 PHY_667 ();
 sky130_fd_sc_hd__decap_3 PHY_668 ();
 sky130_fd_sc_hd__decap_3 PHY_669 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_670 ();
 sky130_fd_sc_hd__decap_3 PHY_671 ();
 sky130_fd_sc_hd__decap_3 PHY_672 ();
 sky130_fd_sc_hd__decap_3 PHY_673 ();
 sky130_fd_sc_hd__decap_3 PHY_674 ();
 sky130_fd_sc_hd__decap_3 PHY_675 ();
 sky130_fd_sc_hd__decap_3 PHY_676 ();
 sky130_fd_sc_hd__decap_3 PHY_677 ();
 sky130_fd_sc_hd__decap_3 PHY_678 ();
 sky130_fd_sc_hd__decap_3 PHY_679 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_680 ();
 sky130_fd_sc_hd__decap_3 PHY_681 ();
 sky130_fd_sc_hd__decap_3 PHY_682 ();
 sky130_fd_sc_hd__decap_3 PHY_683 ();
 sky130_fd_sc_hd__decap_3 PHY_684 ();
 sky130_fd_sc_hd__decap_3 PHY_685 ();
 sky130_fd_sc_hd__decap_3 PHY_686 ();
 sky130_fd_sc_hd__decap_3 PHY_687 ();
 sky130_fd_sc_hd__decap_3 PHY_688 ();
 sky130_fd_sc_hd__decap_3 PHY_689 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_690 ();
 sky130_fd_sc_hd__decap_3 PHY_691 ();
 sky130_fd_sc_hd__decap_3 PHY_692 ();
 sky130_fd_sc_hd__decap_3 PHY_693 ();
 sky130_fd_sc_hd__decap_3 PHY_694 ();
 sky130_fd_sc_hd__decap_3 PHY_695 ();
 sky130_fd_sc_hd__decap_3 PHY_696 ();
 sky130_fd_sc_hd__decap_3 PHY_697 ();
 sky130_fd_sc_hd__decap_3 PHY_698 ();
 sky130_fd_sc_hd__decap_3 PHY_699 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_700 ();
 sky130_fd_sc_hd__decap_3 PHY_701 ();
 sky130_fd_sc_hd__decap_3 PHY_702 ();
 sky130_fd_sc_hd__decap_3 PHY_703 ();
 sky130_fd_sc_hd__decap_3 PHY_704 ();
 sky130_fd_sc_hd__decap_3 PHY_705 ();
 sky130_fd_sc_hd__decap_3 PHY_706 ();
 sky130_fd_sc_hd__decap_3 PHY_707 ();
 sky130_fd_sc_hd__decap_3 PHY_708 ();
 sky130_fd_sc_hd__decap_3 PHY_709 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_710 ();
 sky130_fd_sc_hd__decap_3 PHY_711 ();
 sky130_fd_sc_hd__decap_3 PHY_712 ();
 sky130_fd_sc_hd__decap_3 PHY_713 ();
 sky130_fd_sc_hd__decap_3 PHY_714 ();
 sky130_fd_sc_hd__decap_3 PHY_715 ();
 sky130_fd_sc_hd__decap_3 PHY_716 ();
 sky130_fd_sc_hd__decap_3 PHY_717 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__inv_2 _0396_ (.A(net477),
    .Y(_0113_));
 sky130_fd_sc_hd__mux2_8 _0397_ (.A0(net1),
    .A1(net1116),
    .S(net847),
    .X(net394));
 sky130_fd_sc_hd__nor2_1 _0398_ (.A(net586),
    .B(net571),
    .Y(_0114_));
 sky130_fd_sc_hd__and3b_2 _0399_ (.A_N(net559),
    .B(net580),
    .C(net572),
    .X(_0115_));
 sky130_fd_sc_hd__and2_1 _0400_ (.A(net394),
    .B(net464),
    .X(net403));
 sky130_fd_sc_hd__and3b_4 _0401_ (.A_N(net564),
    .B(net572),
    .C(net559),
    .X(_0116_));
 sky130_fd_sc_hd__and2_2 _0402_ (.A(net394),
    .B(_0116_),
    .X(net401));
 sky130_fd_sc_hd__and3_2 _0403_ (.A(net559),
    .B(net564),
    .C(net572),
    .X(_0117_));
 sky130_fd_sc_hd__and2_2 _0404_ (.A(net394),
    .B(net456),
    .X(net402));
 sky130_fd_sc_hd__o21ai_1 _0405_ (.A1(net559),
    .A2(net564),
    .B1(net572),
    .Y(_0118_));
 sky130_fd_sc_hd__a22o_1 _0406_ (.A1(net109),
    .A2(net466),
    .B1(net456),
    .B2(net73),
    .X(_0119_));
 sky130_fd_sc_hd__a211o_4 _0407_ (.A1(net37),
    .A2(net461),
    .B1(net451),
    .C1(_0119_),
    .X(net291));
 sky130_fd_sc_hd__a22o_1 _0408_ (.A1(net75),
    .A2(net466),
    .B1(net456),
    .B2(net39),
    .X(_0120_));
 sky130_fd_sc_hd__a211o_4 _0409_ (.A1(net3),
    .A2(net461),
    .B1(net451),
    .C1(_0120_),
    .X(net292));
 sky130_fd_sc_hd__a22o_1 _0410_ (.A1(net76),
    .A2(net466),
    .B1(net456),
    .B2(net40),
    .X(_0121_));
 sky130_fd_sc_hd__a211o_4 _0411_ (.A1(net4),
    .A2(net461),
    .B1(net451),
    .C1(_0121_),
    .X(net293));
 sky130_fd_sc_hd__a22o_1 _0412_ (.A1(net77),
    .A2(net466),
    .B1(net456),
    .B2(net41),
    .X(_0122_));
 sky130_fd_sc_hd__a211o_4 _0413_ (.A1(net5),
    .A2(net461),
    .B1(net451),
    .C1(_0122_),
    .X(net294));
 sky130_fd_sc_hd__a22o_1 _0414_ (.A1(net78),
    .A2(net466),
    .B1(net456),
    .B2(net42),
    .X(_0123_));
 sky130_fd_sc_hd__a211o_4 _0415_ (.A1(net6),
    .A2(net461),
    .B1(net450),
    .C1(_0123_),
    .X(net295));
 sky130_fd_sc_hd__a22o_1 _0416_ (.A1(net79),
    .A2(net466),
    .B1(net456),
    .B2(net43),
    .X(_0124_));
 sky130_fd_sc_hd__a211o_4 _0417_ (.A1(net7),
    .A2(net461),
    .B1(net450),
    .C1(_0124_),
    .X(net296));
 sky130_fd_sc_hd__a22o_1 _0418_ (.A1(net80),
    .A2(net466),
    .B1(net456),
    .B2(net44),
    .X(_0125_));
 sky130_fd_sc_hd__a211o_4 _0419_ (.A1(net8),
    .A2(net461),
    .B1(net450),
    .C1(_0125_),
    .X(net297));
 sky130_fd_sc_hd__a22o_1 _0420_ (.A1(net81),
    .A2(net466),
    .B1(net456),
    .B2(net45),
    .X(_0126_));
 sky130_fd_sc_hd__a211o_4 _0421_ (.A1(net9),
    .A2(net461),
    .B1(net450),
    .C1(_0126_),
    .X(net298));
 sky130_fd_sc_hd__a22o_1 _0422_ (.A1(net82),
    .A2(net466),
    .B1(net456),
    .B2(net46),
    .X(_0127_));
 sky130_fd_sc_hd__a211o_4 _0423_ (.A1(net10),
    .A2(net461),
    .B1(net450),
    .C1(_0127_),
    .X(net299));
 sky130_fd_sc_hd__a22o_1 _0424_ (.A1(net83),
    .A2(net465),
    .B1(net455),
    .B2(net47),
    .X(_0128_));
 sky130_fd_sc_hd__a211o_4 _0425_ (.A1(net11),
    .A2(net460),
    .B1(net450),
    .C1(_0128_),
    .X(net301));
 sky130_fd_sc_hd__a22o_1 _0426_ (.A1(net84),
    .A2(net465),
    .B1(net455),
    .B2(net48),
    .X(_0129_));
 sky130_fd_sc_hd__a211o_4 _0427_ (.A1(net12),
    .A2(net460),
    .B1(net450),
    .C1(_0129_),
    .X(net302));
 sky130_fd_sc_hd__a22o_1 _0428_ (.A1(net86),
    .A2(net465),
    .B1(net455),
    .B2(net50),
    .X(_0130_));
 sky130_fd_sc_hd__a211o_4 _0429_ (.A1(net14),
    .A2(net460),
    .B1(net450),
    .C1(_0130_),
    .X(net303));
 sky130_fd_sc_hd__a22o_1 _0430_ (.A1(net87),
    .A2(net465),
    .B1(net455),
    .B2(net51),
    .X(_0131_));
 sky130_fd_sc_hd__a211o_4 _0431_ (.A1(net15),
    .A2(net460),
    .B1(net450),
    .C1(_0131_),
    .X(net304));
 sky130_fd_sc_hd__a22o_1 _0432_ (.A1(net88),
    .A2(net465),
    .B1(net455),
    .B2(net52),
    .X(_0132_));
 sky130_fd_sc_hd__a211o_4 _0433_ (.A1(net16),
    .A2(net460),
    .B1(net450),
    .C1(_0132_),
    .X(net305));
 sky130_fd_sc_hd__a22o_1 _0434_ (.A1(net89),
    .A2(net465),
    .B1(net455),
    .B2(net53),
    .X(_0133_));
 sky130_fd_sc_hd__a211o_4 _0435_ (.A1(net17),
    .A2(net460),
    .B1(net450),
    .C1(_0133_),
    .X(net306));
 sky130_fd_sc_hd__a22o_1 _0436_ (.A1(net90),
    .A2(net465),
    .B1(net455),
    .B2(net54),
    .X(_0134_));
 sky130_fd_sc_hd__a211o_4 _0437_ (.A1(net18),
    .A2(net460),
    .B1(net449),
    .C1(_0134_),
    .X(net307));
 sky130_fd_sc_hd__a22o_1 _0438_ (.A1(net91),
    .A2(net465),
    .B1(net455),
    .B2(net55),
    .X(_0135_));
 sky130_fd_sc_hd__a211o_4 _0439_ (.A1(net19),
    .A2(net460),
    .B1(net449),
    .C1(_0135_),
    .X(net308));
 sky130_fd_sc_hd__a22o_1 _0440_ (.A1(net92),
    .A2(net466),
    .B1(net456),
    .B2(net56),
    .X(_0136_));
 sky130_fd_sc_hd__a211o_4 _0441_ (.A1(net20),
    .A2(net461),
    .B1(net449),
    .C1(_0136_),
    .X(net309));
 sky130_fd_sc_hd__a22o_1 _0442_ (.A1(net93),
    .A2(net466),
    .B1(net456),
    .B2(net57),
    .X(_0137_));
 sky130_fd_sc_hd__a211o_4 _0443_ (.A1(net21),
    .A2(net460),
    .B1(net449),
    .C1(_0137_),
    .X(net310));
 sky130_fd_sc_hd__a22o_1 _0444_ (.A1(net94),
    .A2(net465),
    .B1(net455),
    .B2(net58),
    .X(_0138_));
 sky130_fd_sc_hd__a211o_4 _0445_ (.A1(net22),
    .A2(net460),
    .B1(net449),
    .C1(_0138_),
    .X(net312));
 sky130_fd_sc_hd__a22o_1 _0446_ (.A1(net95),
    .A2(net465),
    .B1(net455),
    .B2(net59),
    .X(_0139_));
 sky130_fd_sc_hd__a211o_4 _0447_ (.A1(net23),
    .A2(net460),
    .B1(net449),
    .C1(_0139_),
    .X(net313));
 sky130_fd_sc_hd__a22o_1 _0448_ (.A1(net97),
    .A2(net465),
    .B1(net455),
    .B2(net61),
    .X(_0140_));
 sky130_fd_sc_hd__a211o_4 _0449_ (.A1(net25),
    .A2(net460),
    .B1(net449),
    .C1(_0140_),
    .X(net314));
 sky130_fd_sc_hd__a22o_1 _0450_ (.A1(net98),
    .A2(net465),
    .B1(net455),
    .B2(net62),
    .X(_0141_));
 sky130_fd_sc_hd__a211o_4 _0451_ (.A1(net26),
    .A2(net460),
    .B1(net449),
    .C1(_0141_),
    .X(net315));
 sky130_fd_sc_hd__a22o_1 _0452_ (.A1(net99),
    .A2(net465),
    .B1(net455),
    .B2(net63),
    .X(_0142_));
 sky130_fd_sc_hd__a211o_4 _0453_ (.A1(net27),
    .A2(net460),
    .B1(net449),
    .C1(_0142_),
    .X(net316));
 sky130_fd_sc_hd__a22o_1 _0454_ (.A1(net100),
    .A2(net465),
    .B1(net455),
    .B2(net64),
    .X(_0143_));
 sky130_fd_sc_hd__a211o_4 _0455_ (.A1(net28),
    .A2(net460),
    .B1(net449),
    .C1(_0143_),
    .X(net317));
 sky130_fd_sc_hd__a22o_1 _0456_ (.A1(net101),
    .A2(net465),
    .B1(net455),
    .B2(net65),
    .X(_0144_));
 sky130_fd_sc_hd__a211o_4 _0457_ (.A1(net29),
    .A2(net461),
    .B1(net449),
    .C1(_0144_),
    .X(net318));
 sky130_fd_sc_hd__a22o_1 _0458_ (.A1(net102),
    .A2(net465),
    .B1(net455),
    .B2(net66),
    .X(_0145_));
 sky130_fd_sc_hd__a211o_4 _0459_ (.A1(net30),
    .A2(net460),
    .B1(net449),
    .C1(_0145_),
    .X(net319));
 sky130_fd_sc_hd__a22o_1 _0460_ (.A1(net182),
    .A2(net462),
    .B1(net452),
    .B2(net146),
    .X(_0146_));
 sky130_fd_sc_hd__a21o_4 _0461_ (.A1(net110),
    .A2(net457),
    .B1(_0146_),
    .X(net336));
 sky130_fd_sc_hd__a22o_1 _0462_ (.A1(net193),
    .A2(net462),
    .B1(net452),
    .B2(net157),
    .X(_0147_));
 sky130_fd_sc_hd__a21o_4 _0463_ (.A1(net121),
    .A2(net457),
    .B1(_0147_),
    .X(net347));
 sky130_fd_sc_hd__a22o_1 _0464_ (.A1(net204),
    .A2(net462),
    .B1(net452),
    .B2(net168),
    .X(_0148_));
 sky130_fd_sc_hd__a21o_4 _0465_ (.A1(net132),
    .A2(net457),
    .B1(_0148_),
    .X(net357));
 sky130_fd_sc_hd__a22o_1 _0466_ (.A1(net211),
    .A2(net462),
    .B1(net452),
    .B2(net175),
    .X(_0149_));
 sky130_fd_sc_hd__a21o_4 _0467_ (.A1(net139),
    .A2(net457),
    .B1(_0149_),
    .X(net358));
 sky130_fd_sc_hd__a22o_1 _0468_ (.A1(net212),
    .A2(net462),
    .B1(net452),
    .B2(net176),
    .X(_0150_));
 sky130_fd_sc_hd__a21o_4 _0469_ (.A1(net140),
    .A2(net457),
    .B1(_0150_),
    .X(net359));
 sky130_fd_sc_hd__a22o_1 _0470_ (.A1(net213),
    .A2(net462),
    .B1(net452),
    .B2(net177),
    .X(_0151_));
 sky130_fd_sc_hd__a21o_4 _0471_ (.A1(net141),
    .A2(net457),
    .B1(_0151_),
    .X(net360));
 sky130_fd_sc_hd__a22o_1 _0472_ (.A1(net214),
    .A2(net462),
    .B1(net452),
    .B2(net178),
    .X(_0152_));
 sky130_fd_sc_hd__a21o_4 _0473_ (.A1(net142),
    .A2(net457),
    .B1(_0152_),
    .X(net361));
 sky130_fd_sc_hd__a22o_1 _0474_ (.A1(net215),
    .A2(net462),
    .B1(net452),
    .B2(net179),
    .X(_0153_));
 sky130_fd_sc_hd__a21o_4 _0475_ (.A1(net143),
    .A2(net457),
    .B1(_0153_),
    .X(net362));
 sky130_fd_sc_hd__a22o_1 _0476_ (.A1(net216),
    .A2(net462),
    .B1(net452),
    .B2(net180),
    .X(_0154_));
 sky130_fd_sc_hd__a21o_4 _0477_ (.A1(net144),
    .A2(net457),
    .B1(_0154_),
    .X(net326));
 sky130_fd_sc_hd__a22o_1 _0478_ (.A1(net217),
    .A2(net462),
    .B1(net452),
    .B2(net181),
    .X(_0155_));
 sky130_fd_sc_hd__a21o_4 _0479_ (.A1(net145),
    .A2(net457),
    .B1(_0155_),
    .X(net327));
 sky130_fd_sc_hd__a22o_1 _0480_ (.A1(net183),
    .A2(net462),
    .B1(net452),
    .B2(net147),
    .X(_0156_));
 sky130_fd_sc_hd__a21o_4 _0481_ (.A1(net111),
    .A2(net457),
    .B1(_0156_),
    .X(net328));
 sky130_fd_sc_hd__a22o_1 _0482_ (.A1(net184),
    .A2(net462),
    .B1(net452),
    .B2(net148),
    .X(_0157_));
 sky130_fd_sc_hd__a21o_4 _0483_ (.A1(net112),
    .A2(net457),
    .B1(_0157_),
    .X(net329));
 sky130_fd_sc_hd__a22o_1 _0484_ (.A1(net185),
    .A2(net462),
    .B1(net452),
    .B2(net149),
    .X(_0158_));
 sky130_fd_sc_hd__a21o_4 _0485_ (.A1(net113),
    .A2(net457),
    .B1(_0158_),
    .X(net330));
 sky130_fd_sc_hd__a22o_1 _0486_ (.A1(net186),
    .A2(net462),
    .B1(net452),
    .B2(net150),
    .X(_0159_));
 sky130_fd_sc_hd__a21o_4 _0487_ (.A1(net114),
    .A2(net457),
    .B1(_0159_),
    .X(net331));
 sky130_fd_sc_hd__a22o_1 _0488_ (.A1(net187),
    .A2(net462),
    .B1(net452),
    .B2(net151),
    .X(_0160_));
 sky130_fd_sc_hd__a21o_4 _0489_ (.A1(net115),
    .A2(net457),
    .B1(_0160_),
    .X(net332));
 sky130_fd_sc_hd__a22o_1 _0490_ (.A1(net188),
    .A2(net462),
    .B1(net452),
    .B2(net152),
    .X(_0161_));
 sky130_fd_sc_hd__a21o_4 _0491_ (.A1(net116),
    .A2(net457),
    .B1(_0161_),
    .X(net333));
 sky130_fd_sc_hd__a22o_1 _0492_ (.A1(net189),
    .A2(net464),
    .B1(net453),
    .B2(net153),
    .X(_0162_));
 sky130_fd_sc_hd__a21o_4 _0493_ (.A1(net117),
    .A2(net458),
    .B1(_0162_),
    .X(net334));
 sky130_fd_sc_hd__a22o_1 _0494_ (.A1(net190),
    .A2(net464),
    .B1(net453),
    .B2(net154),
    .X(_0163_));
 sky130_fd_sc_hd__a21o_4 _0495_ (.A1(net118),
    .A2(net458),
    .B1(_0163_),
    .X(net335));
 sky130_fd_sc_hd__a22o_1 _0496_ (.A1(net191),
    .A2(net464),
    .B1(net453),
    .B2(net155),
    .X(_0164_));
 sky130_fd_sc_hd__a21o_4 _0497_ (.A1(net119),
    .A2(net458),
    .B1(_0164_),
    .X(net337));
 sky130_fd_sc_hd__a22o_1 _0498_ (.A1(net192),
    .A2(net463),
    .B1(net453),
    .B2(net156),
    .X(_0165_));
 sky130_fd_sc_hd__a21o_4 _0499_ (.A1(net120),
    .A2(net458),
    .B1(_0165_),
    .X(net338));
 sky130_fd_sc_hd__a22o_1 _0500_ (.A1(net194),
    .A2(net463),
    .B1(net453),
    .B2(net158),
    .X(_0166_));
 sky130_fd_sc_hd__a21o_4 _0501_ (.A1(net122),
    .A2(net458),
    .B1(_0166_),
    .X(net339));
 sky130_fd_sc_hd__a22o_1 _0502_ (.A1(net195),
    .A2(net463),
    .B1(net453),
    .B2(net159),
    .X(_0167_));
 sky130_fd_sc_hd__a21o_4 _0503_ (.A1(net123),
    .A2(net458),
    .B1(_0167_),
    .X(net340));
 sky130_fd_sc_hd__a22o_1 _0504_ (.A1(net196),
    .A2(net463),
    .B1(net453),
    .B2(net160),
    .X(_0168_));
 sky130_fd_sc_hd__a21o_4 _0505_ (.A1(net124),
    .A2(net458),
    .B1(_0168_),
    .X(net341));
 sky130_fd_sc_hd__a22o_1 _0506_ (.A1(net197),
    .A2(net463),
    .B1(net453),
    .B2(net161),
    .X(_0169_));
 sky130_fd_sc_hd__a21o_4 _0507_ (.A1(net125),
    .A2(net458),
    .B1(_0169_),
    .X(net342));
 sky130_fd_sc_hd__a22o_1 _0508_ (.A1(net198),
    .A2(net463),
    .B1(net454),
    .B2(net162),
    .X(_0170_));
 sky130_fd_sc_hd__a21o_4 _0509_ (.A1(net126),
    .A2(net459),
    .B1(_0170_),
    .X(net343));
 sky130_fd_sc_hd__a22o_1 _0510_ (.A1(net199),
    .A2(net463),
    .B1(net454),
    .B2(net163),
    .X(_0171_));
 sky130_fd_sc_hd__a21o_4 _0511_ (.A1(net127),
    .A2(net459),
    .B1(_0171_),
    .X(net344));
 sky130_fd_sc_hd__a22o_1 _0512_ (.A1(net200),
    .A2(net463),
    .B1(net454),
    .B2(net164),
    .X(_0172_));
 sky130_fd_sc_hd__a21o_4 _0513_ (.A1(net128),
    .A2(net459),
    .B1(_0172_),
    .X(net345));
 sky130_fd_sc_hd__a22o_1 _0514_ (.A1(net201),
    .A2(net463),
    .B1(net454),
    .B2(net165),
    .X(_0173_));
 sky130_fd_sc_hd__a21o_4 _0515_ (.A1(net129),
    .A2(net459),
    .B1(_0173_),
    .X(net346));
 sky130_fd_sc_hd__a22o_1 _0516_ (.A1(net202),
    .A2(net463),
    .B1(net453),
    .B2(net166),
    .X(_0174_));
 sky130_fd_sc_hd__a21o_4 _0517_ (.A1(net130),
    .A2(net458),
    .B1(_0174_),
    .X(net348));
 sky130_fd_sc_hd__a22o_1 _0518_ (.A1(net203),
    .A2(net463),
    .B1(net453),
    .B2(net167),
    .X(_0175_));
 sky130_fd_sc_hd__a21o_4 _0519_ (.A1(net131),
    .A2(net458),
    .B1(_0175_),
    .X(net349));
 sky130_fd_sc_hd__a22o_1 _0520_ (.A1(net205),
    .A2(net463),
    .B1(net453),
    .B2(net169),
    .X(_0176_));
 sky130_fd_sc_hd__a21o_4 _0521_ (.A1(net133),
    .A2(net458),
    .B1(_0176_),
    .X(net350));
 sky130_fd_sc_hd__a22o_1 _0522_ (.A1(net206),
    .A2(net463),
    .B1(net453),
    .B2(net170),
    .X(_0177_));
 sky130_fd_sc_hd__a21o_4 _0523_ (.A1(net134),
    .A2(net458),
    .B1(_0177_),
    .X(net351));
 sky130_fd_sc_hd__a22o_1 _0524_ (.A1(net207),
    .A2(net463),
    .B1(net453),
    .B2(net171),
    .X(_0178_));
 sky130_fd_sc_hd__a21o_4 _0525_ (.A1(net135),
    .A2(net458),
    .B1(_0178_),
    .X(net352));
 sky130_fd_sc_hd__a22o_1 _0526_ (.A1(net208),
    .A2(net463),
    .B1(net453),
    .B2(net172),
    .X(_0179_));
 sky130_fd_sc_hd__a21o_4 _0527_ (.A1(net136),
    .A2(net458),
    .B1(_0179_),
    .X(net353));
 sky130_fd_sc_hd__a22o_1 _0528_ (.A1(net209),
    .A2(net463),
    .B1(net453),
    .B2(net173),
    .X(_0180_));
 sky130_fd_sc_hd__a21o_4 _0529_ (.A1(net137),
    .A2(net458),
    .B1(_0180_),
    .X(net354));
 sky130_fd_sc_hd__a22o_1 _0530_ (.A1(net210),
    .A2(_0115_),
    .B1(_0117_),
    .B2(net174),
    .X(_0181_));
 sky130_fd_sc_hd__a21o_4 _0531_ (.A1(net138),
    .A2(_0116_),
    .B1(_0181_),
    .X(net355));
 sky130_fd_sc_hd__a22o_1 _0532_ (.A1(net74),
    .A2(net464),
    .B1(net566),
    .B2(net38),
    .X(_0182_));
 sky130_fd_sc_hd__a211o_4 _0533_ (.A1(net2),
    .A2(net459),
    .B1(net560),
    .C1(net567),
    .X(net300));
 sky130_fd_sc_hd__a22o_1 _0534_ (.A1(net85),
    .A2(net464),
    .B1(net566),
    .B2(net49),
    .X(_0183_));
 sky130_fd_sc_hd__a211o_4 _0535_ (.A1(net13),
    .A2(net574),
    .B1(net560),
    .C1(_0183_),
    .X(net311));
 sky130_fd_sc_hd__a22o_1 _0536_ (.A1(net96),
    .A2(net464),
    .B1(net454),
    .B2(net60),
    .X(_0184_));
 sky130_fd_sc_hd__a211o_4 _0537_ (.A1(net24),
    .A2(net459),
    .B1(net560),
    .C1(_0184_),
    .X(net320));
 sky130_fd_sc_hd__a22o_1 _0538_ (.A1(net103),
    .A2(net464),
    .B1(net566),
    .B2(net67),
    .X(_0185_));
 sky130_fd_sc_hd__a211o_4 _0539_ (.A1(net31),
    .A2(net574),
    .B1(net451),
    .C1(_0185_),
    .X(net321));
 sky130_fd_sc_hd__a22o_1 _0540_ (.A1(net104),
    .A2(net464),
    .B1(net566),
    .B2(net68),
    .X(_0186_));
 sky130_fd_sc_hd__a211o_4 _0541_ (.A1(net32),
    .A2(net574),
    .B1(net451),
    .C1(_0186_),
    .X(net322));
 sky130_fd_sc_hd__a22o_1 _0542_ (.A1(net105),
    .A2(net464),
    .B1(net566),
    .B2(net69),
    .X(_0187_));
 sky130_fd_sc_hd__a211o_4 _0543_ (.A1(net33),
    .A2(net574),
    .B1(net451),
    .C1(_0187_),
    .X(net323));
 sky130_fd_sc_hd__a22o_1 _0544_ (.A1(net106),
    .A2(net466),
    .B1(net456),
    .B2(net70),
    .X(_0188_));
 sky130_fd_sc_hd__a211o_4 _0545_ (.A1(net34),
    .A2(net461),
    .B1(net451),
    .C1(_0188_),
    .X(net324));
 sky130_fd_sc_hd__a22o_1 _0546_ (.A1(net107),
    .A2(net466),
    .B1(net456),
    .B2(net71),
    .X(_0189_));
 sky130_fd_sc_hd__a211o_4 _0547_ (.A1(net35),
    .A2(net461),
    .B1(net451),
    .C1(_0189_),
    .X(net325));
 sky130_fd_sc_hd__a22o_1 _0548_ (.A1(net108),
    .A2(net466),
    .B1(net456),
    .B2(net72),
    .X(_0190_));
 sky130_fd_sc_hd__a211o_4 _0549_ (.A1(net36),
    .A2(net461),
    .B1(net451),
    .C1(_0190_),
    .X(net290));
 sky130_fd_sc_hd__and2_2 _0550_ (.A(net256),
    .B(net223),
    .X(_0191_));
 sky130_fd_sc_hd__mux2_1 _0551_ (.A0(net604),
    .A1(net1172),
    .S(net474),
    .X(_0000_));
 sky130_fd_sc_hd__nand3b_1 _0552_ (.A_N(net856),
    .B(net1080),
    .C(net1174),
    .Y(_0192_));
 sky130_fd_sc_hd__and3b_1 _0553_ (.A_N(net923),
    .B(_0191_),
    .C(net604),
    .X(_0193_));
 sky130_fd_sc_hd__and2_1 _0554_ (.A(net870),
    .B(_0193_),
    .X(_0194_));
 sky130_fd_sc_hd__nand2_1 _0555_ (.A(net870),
    .B(_0193_),
    .Y(_0195_));
 sky130_fd_sc_hd__nand2_1 _0556_ (.A(net257),
    .B(net871),
    .Y(_0196_));
 sky130_fd_sc_hd__nor2_1 _0557_ (.A(net469),
    .B(net872),
    .Y(_0197_));
 sky130_fd_sc_hd__or2_1 _0558_ (.A(net469),
    .B(net1180),
    .X(_0198_));
 sky130_fd_sc_hd__or2_1 _0559_ (.A(net1031),
    .B(net443),
    .X(_0199_));
 sky130_fd_sc_hd__o211a_1 _0560_ (.A1(net845),
    .A2(net441),
    .B1(net1032),
    .C1(net473),
    .X(_0001_));
 sky130_fd_sc_hd__or2_1 _0561_ (.A(net1110),
    .B(net444),
    .X(_0200_));
 sky130_fd_sc_hd__o211a_1 _0562_ (.A1(net854),
    .A2(net442),
    .B1(net1111),
    .C1(net473),
    .X(_0002_));
 sky130_fd_sc_hd__or2_1 _0563_ (.A(net1113),
    .B(net444),
    .X(_0201_));
 sky130_fd_sc_hd__o211a_1 _0564_ (.A1(net852),
    .A2(net442),
    .B1(net1114),
    .C1(net473),
    .X(_0003_));
 sky130_fd_sc_hd__or2_1 _0565_ (.A(net699),
    .B(net444),
    .X(_0202_));
 sky130_fd_sc_hd__o211a_1 _0566_ (.A1(net697),
    .A2(net442),
    .B1(net700),
    .C1(net471),
    .X(_0004_));
 sky130_fd_sc_hd__or2_1 _0567_ (.A(net819),
    .B(net444),
    .X(_0203_));
 sky130_fd_sc_hd__o211a_1 _0568_ (.A1(net817),
    .A2(net442),
    .B1(net820),
    .C1(net471),
    .X(_0005_));
 sky130_fd_sc_hd__or2_1 _0569_ (.A(net1095),
    .B(net444),
    .X(_0204_));
 sky130_fd_sc_hd__o211a_1 _0570_ (.A1(net793),
    .A2(net442),
    .B1(net1096),
    .C1(net472),
    .X(_0006_));
 sky130_fd_sc_hd__or2_1 _0571_ (.A(net1104),
    .B(net444),
    .X(_0205_));
 sky130_fd_sc_hd__o211a_1 _0572_ (.A1(net864),
    .A2(net442),
    .B1(net1105),
    .C1(net471),
    .X(_0007_));
 sky130_fd_sc_hd__or2_1 _0573_ (.A(net1101),
    .B(net444),
    .X(_0206_));
 sky130_fd_sc_hd__o211a_1 _0574_ (.A1(net666),
    .A2(net442),
    .B1(net1102),
    .C1(net471),
    .X(_0008_));
 sky130_fd_sc_hd__or2_1 _0575_ (.A(net670),
    .B(net444),
    .X(_0207_));
 sky130_fd_sc_hd__o211a_1 _0576_ (.A1(net664),
    .A2(net442),
    .B1(net671),
    .C1(net471),
    .X(_0009_));
 sky130_fd_sc_hd__or2_1 _0577_ (.A(net1064),
    .B(net444),
    .X(_0208_));
 sky130_fd_sc_hd__o211a_1 _0578_ (.A1(net631),
    .A2(net442),
    .B1(net1065),
    .C1(net471),
    .X(_0010_));
 sky130_fd_sc_hd__or2_1 _0579_ (.A(net647),
    .B(net444),
    .X(_0209_));
 sky130_fd_sc_hd__o211a_1 _0580_ (.A1(net645),
    .A2(net442),
    .B1(net648),
    .C1(net471),
    .X(_0011_));
 sky130_fd_sc_hd__or2_1 _0581_ (.A(net1074),
    .B(net444),
    .X(_0210_));
 sky130_fd_sc_hd__o211a_1 _0582_ (.A1(net650),
    .A2(net442),
    .B1(net1075),
    .C1(net471),
    .X(_0012_));
 sky130_fd_sc_hd__or2_1 _0583_ (.A(net640),
    .B(net444),
    .X(_0211_));
 sky130_fd_sc_hd__o211a_1 _0584_ (.A1(net626),
    .A2(net442),
    .B1(net641),
    .C1(net471),
    .X(_0013_));
 sky130_fd_sc_hd__or2_1 _0585_ (.A(net1097),
    .B(net444),
    .X(_0212_));
 sky130_fd_sc_hd__o211a_1 _0586_ (.A1(net577),
    .A2(net442),
    .B1(net1098),
    .C1(net473),
    .X(_0014_));
 sky130_fd_sc_hd__or2_1 _0587_ (.A(net628),
    .B(net444),
    .X(_0213_));
 sky130_fd_sc_hd__o211a_1 _0588_ (.A1(net616),
    .A2(net442),
    .B1(net629),
    .C1(net473),
    .X(_0015_));
 sky130_fd_sc_hd__or2_1 _0589_ (.A(net637),
    .B(net444),
    .X(_0214_));
 sky130_fd_sc_hd__o211a_1 _0590_ (.A1(net614),
    .A2(net442),
    .B1(net638),
    .C1(net473),
    .X(_0016_));
 sky130_fd_sc_hd__or2_1 _0591_ (.A(net1061),
    .B(net443),
    .X(_0215_));
 sky130_fd_sc_hd__o211a_1 _0592_ (.A1(net608),
    .A2(net441),
    .B1(net1062),
    .C1(net473),
    .X(_0017_));
 sky130_fd_sc_hd__or2_1 _0593_ (.A(net1092),
    .B(net443),
    .X(_0216_));
 sky130_fd_sc_hd__o211a_1 _0594_ (.A1(net702),
    .A2(net441),
    .B1(net1093),
    .C1(net473),
    .X(_0018_));
 sky130_fd_sc_hd__or2_1 _0595_ (.A(net1086),
    .B(net443),
    .X(_0217_));
 sky130_fd_sc_hd__o211a_1 _0596_ (.A1(net681),
    .A2(net441),
    .B1(net1087),
    .C1(net475),
    .X(_0019_));
 sky130_fd_sc_hd__or2_1 _0597_ (.A(net795),
    .B(net443),
    .X(_0218_));
 sky130_fd_sc_hd__o211a_1 _0598_ (.A1(net714),
    .A2(net441),
    .B1(net796),
    .C1(net475),
    .X(_0020_));
 sky130_fd_sc_hd__or2_1 _0599_ (.A(net1067),
    .B(net443),
    .X(_0219_));
 sky130_fd_sc_hd__o211a_1 _0600_ (.A1(net704),
    .A2(net441),
    .B1(net1068),
    .C1(net475),
    .X(_0021_));
 sky130_fd_sc_hd__or2_1 _0601_ (.A(net694),
    .B(_0197_),
    .X(_0220_));
 sky130_fd_sc_hd__o211a_1 _0602_ (.A1(net692),
    .A2(_0198_),
    .B1(net695),
    .C1(net475),
    .X(_0022_));
 sky130_fd_sc_hd__or2_1 _0603_ (.A(net689),
    .B(net443),
    .X(_0221_));
 sky130_fd_sc_hd__o211a_1 _0604_ (.A1(net683),
    .A2(net441),
    .B1(net690),
    .C1(net475),
    .X(_0023_));
 sky130_fd_sc_hd__or2_1 _0605_ (.A(net719),
    .B(net443),
    .X(_0222_));
 sky130_fd_sc_hd__o211a_1 _0606_ (.A1(net717),
    .A2(net441),
    .B1(net720),
    .C1(net474),
    .X(_0024_));
 sky130_fd_sc_hd__or2_1 _0607_ (.A(net727),
    .B(net443),
    .X(_0223_));
 sky130_fd_sc_hd__o211a_1 _0608_ (.A1(net725),
    .A2(net441),
    .B1(net728),
    .C1(net474),
    .X(_0025_));
 sky130_fd_sc_hd__or2_1 _0609_ (.A(net1107),
    .B(net443),
    .X(_0224_));
 sky130_fd_sc_hd__o211a_1 _0610_ (.A1(net643),
    .A2(net441),
    .B1(net1108),
    .C1(net474),
    .X(_0026_));
 sky130_fd_sc_hd__or2_1 _0611_ (.A(net1083),
    .B(net443),
    .X(_0225_));
 sky130_fd_sc_hd__o211a_1 _0612_ (.A1(net668),
    .A2(net441),
    .B1(net1084),
    .C1(net475),
    .X(_0027_));
 sky130_fd_sc_hd__or2_1 _0613_ (.A(net1077),
    .B(net443),
    .X(_0226_));
 sky130_fd_sc_hd__o211a_1 _0614_ (.A1(net606),
    .A2(net441),
    .B1(net1078),
    .C1(net474),
    .X(_0028_));
 sky130_fd_sc_hd__or2_1 _0615_ (.A(net1058),
    .B(net443),
    .X(_0227_));
 sky130_fd_sc_hd__o211a_1 _0616_ (.A1(net652),
    .A2(net441),
    .B1(net1059),
    .C1(net474),
    .X(_0029_));
 sky130_fd_sc_hd__or2_1 _0617_ (.A(net1042),
    .B(net443),
    .X(_0228_));
 sky130_fd_sc_hd__o211a_1 _0618_ (.A1(net618),
    .A2(net441),
    .B1(net1043),
    .C1(net474),
    .X(_0030_));
 sky130_fd_sc_hd__or2_1 _0619_ (.A(net1089),
    .B(net443),
    .X(_0229_));
 sky130_fd_sc_hd__o211a_1 _0620_ (.A1(net620),
    .A2(net441),
    .B1(net1090),
    .C1(net474),
    .X(_0031_));
 sky130_fd_sc_hd__or2_1 _0621_ (.A(net1055),
    .B(net443),
    .X(_0230_));
 sky130_fd_sc_hd__o211a_1 _0622_ (.A1(net662),
    .A2(net441),
    .B1(net1056),
    .C1(net476),
    .X(_0032_));
 sky130_fd_sc_hd__or3b_1 _0623_ (.A(net856),
    .B(net1080),
    .C_N(net1174),
    .X(_0231_));
 sky130_fd_sc_hd__nor2_1 _0624_ (.A(net872),
    .B(net857),
    .Y(_0232_));
 sky130_fd_sc_hd__or3_1 _0625_ (.A(net885),
    .B(net872),
    .C(net857),
    .X(_0233_));
 sky130_fd_sc_hd__o211a_1 _0626_ (.A1(net580),
    .A2(net873),
    .B1(net886),
    .C1(net475),
    .X(_0033_));
 sky130_fd_sc_hd__or3_1 _0627_ (.A(net697),
    .B(_0196_),
    .C(net857),
    .X(_0234_));
 sky130_fd_sc_hd__o211a_1 _0628_ (.A1(net584),
    .A2(_0232_),
    .B1(net858),
    .C1(net475),
    .X(_0034_));
 sky130_fd_sc_hd__or3_1 _0629_ (.A(net881),
    .B(net872),
    .C(net857),
    .X(_0235_));
 sky130_fd_sc_hd__o211a_1 _0630_ (.A1(net594),
    .A2(net873),
    .B1(net882),
    .C1(net475),
    .X(_0035_));
 sky130_fd_sc_hd__or3_1 _0631_ (.A(net877),
    .B(net872),
    .C(net857),
    .X(_0236_));
 sky130_fd_sc_hd__o211a_1 _0632_ (.A1(net596),
    .A2(net873),
    .B1(net878),
    .C1(net475),
    .X(_0036_));
 sky130_fd_sc_hd__or3b_4 _0633_ (.A(net856),
    .B(net1119),
    .C_N(net1080),
    .X(_0237_));
 sky130_fd_sc_hd__or2_1 _0634_ (.A(net847),
    .B(net857),
    .X(_0238_));
 sky130_fd_sc_hd__o221a_1 _0635_ (.A1(net1031),
    .A2(net470),
    .B1(net468),
    .B2(net814),
    .C1(_0238_),
    .X(_0239_));
 sky130_fd_sc_hd__or2_1 _0636_ (.A(net447),
    .B(net1128),
    .X(_0240_));
 sky130_fd_sc_hd__o211a_1 _0637_ (.A1(net830),
    .A2(net871),
    .B1(_0240_),
    .C1(net472),
    .X(_0037_));
 sky130_fd_sc_hd__or2_1 _0638_ (.A(net556),
    .B(net857),
    .X(_0241_));
 sky130_fd_sc_hd__o221a_1 _0639_ (.A1(net1110),
    .A2(net470),
    .B1(net468),
    .B2(net860),
    .C1(_0241_),
    .X(_0242_));
 sky130_fd_sc_hd__or2_1 _0640_ (.A(net447),
    .B(net1130),
    .X(_0243_));
 sky130_fd_sc_hd__o211a_1 _0641_ (.A1(net828),
    .A2(net871),
    .B1(_0243_),
    .C1(net472),
    .X(_0038_));
 sky130_fd_sc_hd__or2_1 _0642_ (.A(net564),
    .B(net857),
    .X(_0244_));
 sky130_fd_sc_hd__o221a_1 _0643_ (.A1(net1113),
    .A2(net470),
    .B1(net468),
    .B2(net888),
    .C1(_0244_),
    .X(_0245_));
 sky130_fd_sc_hd__or2_1 _0644_ (.A(net447),
    .B(net1133),
    .X(_0246_));
 sky130_fd_sc_hd__o211a_1 _0645_ (.A1(net826),
    .A2(net871),
    .B1(_0246_),
    .C1(net472),
    .X(_0039_));
 sky130_fd_sc_hd__or2_1 _0646_ (.A(net559),
    .B(net857),
    .X(_0247_));
 sky130_fd_sc_hd__o221a_1 _0647_ (.A1(net699),
    .A2(net470),
    .B1(net468),
    .B2(net1015),
    .C1(_0247_),
    .X(_0248_));
 sky130_fd_sc_hd__or2_1 _0648_ (.A(net447),
    .B(net1082),
    .X(_0249_));
 sky130_fd_sc_hd__o211a_1 _0649_ (.A1(net824),
    .A2(net871),
    .B1(_0249_),
    .C1(net472),
    .X(_0040_));
 sky130_fd_sc_hd__or2_1 _0650_ (.A(net594),
    .B(net857),
    .X(_0250_));
 sky130_fd_sc_hd__o221a_1 _0651_ (.A1(net819),
    .A2(net470),
    .B1(net468),
    .B2(net1045),
    .C1(_0250_),
    .X(_0251_));
 sky130_fd_sc_hd__or2_1 _0652_ (.A(net447),
    .B(net1120),
    .X(_0252_));
 sky130_fd_sc_hd__o211a_1 _0653_ (.A1(net835),
    .A2(net871),
    .B1(_0252_),
    .C1(net472),
    .X(_0041_));
 sky130_fd_sc_hd__or2_1 _0654_ (.A(net596),
    .B(net857),
    .X(_0253_));
 sky130_fd_sc_hd__o221a_1 _0655_ (.A1(net1095),
    .A2(net470),
    .B1(net468),
    .B2(net801),
    .C1(_0253_),
    .X(_0254_));
 sky130_fd_sc_hd__or2_1 _0656_ (.A(net447),
    .B(net1124),
    .X(_0255_));
 sky130_fd_sc_hd__o211a_1 _0657_ (.A1(net837),
    .A2(net871),
    .B1(_0255_),
    .C1(net472),
    .X(_0042_));
 sky130_fd_sc_hd__o22a_1 _0658_ (.A1(net1104),
    .A2(net470),
    .B1(net468),
    .B2(net866),
    .X(_0256_));
 sky130_fd_sc_hd__or2_1 _0659_ (.A(net447),
    .B(net1122),
    .X(_0257_));
 sky130_fd_sc_hd__o211a_1 _0660_ (.A1(net839),
    .A2(net871),
    .B1(_0257_),
    .C1(net472),
    .X(_0043_));
 sky130_fd_sc_hd__o22a_1 _0661_ (.A1(net1101),
    .A2(net470),
    .B1(net468),
    .B2(net677),
    .X(_0258_));
 sky130_fd_sc_hd__or2_1 _0662_ (.A(net447),
    .B(net1126),
    .X(_0259_));
 sky130_fd_sc_hd__o211a_1 _0663_ (.A1(net822),
    .A2(net871),
    .B1(_0259_),
    .C1(net472),
    .X(_0044_));
 sky130_fd_sc_hd__and3_1 _0664_ (.A(net870),
    .B(_0193_),
    .C(_0231_),
    .X(_0260_));
 sky130_fd_sc_hd__o221a_1 _0665_ (.A1(net670),
    .A2(net470),
    .B1(net468),
    .B2(net1038),
    .C1(net445),
    .X(_0261_));
 sky130_fd_sc_hd__a21oi_1 _0666_ (.A1(net790),
    .A2(net447),
    .B1(_0261_),
    .Y(_0262_));
 sky130_fd_sc_hd__nor2_1 _0667_ (.A(net477),
    .B(net791),
    .Y(_0045_));
 sky130_fd_sc_hd__o221a_1 _0668_ (.A1(net1064),
    .A2(net470),
    .B1(net468),
    .B2(net633),
    .C1(net445),
    .X(_0263_));
 sky130_fd_sc_hd__a21oi_1 _0669_ (.A1(net787),
    .A2(net447),
    .B1(_0263_),
    .Y(_0264_));
 sky130_fd_sc_hd__nor2_1 _0670_ (.A(net477),
    .B(net788),
    .Y(_0046_));
 sky130_fd_sc_hd__o221a_1 _0671_ (.A1(net647),
    .A2(net470),
    .B1(net468),
    .B2(net1023),
    .C1(net445),
    .X(_0265_));
 sky130_fd_sc_hd__a21oi_1 _0672_ (.A1(net811),
    .A2(net447),
    .B1(_0265_),
    .Y(_0266_));
 sky130_fd_sc_hd__nor2_1 _0673_ (.A(net477),
    .B(net812),
    .Y(_0047_));
 sky130_fd_sc_hd__o221a_1 _0674_ (.A1(net1074),
    .A2(net470),
    .B1(net468),
    .B2(net658),
    .C1(net445),
    .X(_0267_));
 sky130_fd_sc_hd__a21oi_1 _0675_ (.A1(net730),
    .A2(net448),
    .B1(_0267_),
    .Y(_0268_));
 sky130_fd_sc_hd__nor2_1 _0676_ (.A(net477),
    .B(net731),
    .Y(_0048_));
 sky130_fd_sc_hd__o221a_1 _0677_ (.A1(net640),
    .A2(net470),
    .B1(net468),
    .B2(net1070),
    .C1(net445),
    .X(_0269_));
 sky130_fd_sc_hd__a21oi_1 _0678_ (.A1(net754),
    .A2(net447),
    .B1(_0269_),
    .Y(_0270_));
 sky130_fd_sc_hd__nor2_1 _0679_ (.A(net477),
    .B(net755),
    .Y(_0049_));
 sky130_fd_sc_hd__o221a_1 _0680_ (.A1(net1097),
    .A2(net470),
    .B1(net468),
    .B2(net622),
    .C1(net445),
    .X(_0271_));
 sky130_fd_sc_hd__a21oi_1 _0681_ (.A1(net757),
    .A2(net447),
    .B1(net1238),
    .Y(_0272_));
 sky130_fd_sc_hd__nor2_1 _0682_ (.A(net477),
    .B(net758),
    .Y(_0050_));
 sky130_fd_sc_hd__o221a_1 _0683_ (.A1(net628),
    .A2(net470),
    .B1(net468),
    .B2(net1034),
    .C1(net445),
    .X(_0273_));
 sky130_fd_sc_hd__a21oi_1 _0684_ (.A1(net808),
    .A2(net447),
    .B1(_0273_),
    .Y(_0274_));
 sky130_fd_sc_hd__nor2_1 _0685_ (.A(net477),
    .B(net809),
    .Y(_0051_));
 sky130_fd_sc_hd__o221a_1 _0686_ (.A1(net637),
    .A2(net470),
    .B1(net468),
    .B2(net1019),
    .C1(net445),
    .X(_0275_));
 sky130_fd_sc_hd__a21oi_1 _0687_ (.A1(net766),
    .A2(net447),
    .B1(_0275_),
    .Y(_0276_));
 sky130_fd_sc_hd__nor2_1 _0688_ (.A(net477),
    .B(net767),
    .Y(_0052_));
 sky130_fd_sc_hd__o221a_1 _0689_ (.A1(net1061),
    .A2(net469),
    .B1(net467),
    .B2(net610),
    .C1(net445),
    .X(_0277_));
 sky130_fd_sc_hd__a21oi_1 _0690_ (.A1(net805),
    .A2(net447),
    .B1(_0277_),
    .Y(_0278_));
 sky130_fd_sc_hd__nor2_1 _0691_ (.A(net477),
    .B(net806),
    .Y(_0053_));
 sky130_fd_sc_hd__o221a_1 _0692_ (.A1(net1092),
    .A2(net469),
    .B1(net467),
    .B2(net706),
    .C1(net445),
    .X(_0279_));
 sky130_fd_sc_hd__a21oi_1 _0693_ (.A1(net781),
    .A2(net448),
    .B1(_0279_),
    .Y(_0280_));
 sky130_fd_sc_hd__nor2_1 _0694_ (.A(net477),
    .B(net782),
    .Y(_0054_));
 sky130_fd_sc_hd__o221a_1 _0695_ (.A1(net1086),
    .A2(net469),
    .B1(net467),
    .B2(net685),
    .C1(net445),
    .X(_0281_));
 sky130_fd_sc_hd__a21oi_1 _0696_ (.A1(net748),
    .A2(net448),
    .B1(_0281_),
    .Y(_0282_));
 sky130_fd_sc_hd__nor2_1 _0697_ (.A(net477),
    .B(net749),
    .Y(_0055_));
 sky130_fd_sc_hd__o221a_1 _0698_ (.A1(net795),
    .A2(net469),
    .B1(net467),
    .B2(net1166),
    .C1(net445),
    .X(_0283_));
 sky130_fd_sc_hd__a21oi_1 _0699_ (.A1(net760),
    .A2(net448),
    .B1(_0283_),
    .Y(_0284_));
 sky130_fd_sc_hd__nor2_1 _0700_ (.A(net477),
    .B(net761),
    .Y(_0056_));
 sky130_fd_sc_hd__o221a_1 _0701_ (.A1(net1067),
    .A2(net469),
    .B1(net467),
    .B2(net710),
    .C1(net446),
    .X(_0285_));
 sky130_fd_sc_hd__a21oi_1 _0702_ (.A1(net775),
    .A2(net448),
    .B1(_0285_),
    .Y(_0286_));
 sky130_fd_sc_hd__nor2_1 _0703_ (.A(net477),
    .B(net776),
    .Y(_0057_));
 sky130_fd_sc_hd__o221a_1 _0704_ (.A1(net694),
    .A2(net1081),
    .B1(net467),
    .B2(net1051),
    .C1(net446),
    .X(_0287_));
 sky130_fd_sc_hd__a21oi_1 _0705_ (.A1(net763),
    .A2(_0195_),
    .B1(_0287_),
    .Y(_0288_));
 sky130_fd_sc_hd__nor2_1 _0706_ (.A(net477),
    .B(net764),
    .Y(_0058_));
 sky130_fd_sc_hd__o221a_1 _0707_ (.A1(net689),
    .A2(net1081),
    .B1(net467),
    .B2(net1047),
    .C1(net446),
    .X(_0289_));
 sky130_fd_sc_hd__a21oi_1 _0708_ (.A1(net778),
    .A2(net448),
    .B1(_0289_),
    .Y(_0290_));
 sky130_fd_sc_hd__nor2_1 _0709_ (.A(net477),
    .B(net779),
    .Y(_0059_));
 sky130_fd_sc_hd__o221a_1 _0710_ (.A1(net719),
    .A2(net469),
    .B1(net467),
    .B2(net1027),
    .C1(net446),
    .X(_0291_));
 sky130_fd_sc_hd__a21oi_1 _0711_ (.A1(net742),
    .A2(net448),
    .B1(_0291_),
    .Y(_0292_));
 sky130_fd_sc_hd__nor2_1 _0712_ (.A(net478),
    .B(net743),
    .Y(_0060_));
 sky130_fd_sc_hd__o221a_1 _0713_ (.A1(net727),
    .A2(net469),
    .B1(net467),
    .B2(net841),
    .C1(net446),
    .X(_0293_));
 sky130_fd_sc_hd__a21oi_1 _0714_ (.A1(net772),
    .A2(net448),
    .B1(_0293_),
    .Y(_0294_));
 sky130_fd_sc_hd__nor2_1 _0715_ (.A(net478),
    .B(net773),
    .Y(_0061_));
 sky130_fd_sc_hd__o221a_1 _0716_ (.A1(net1107),
    .A2(net469),
    .B1(net467),
    .B2(net1173),
    .C1(net445),
    .X(_0295_));
 sky130_fd_sc_hd__a21oi_1 _0717_ (.A1(net751),
    .A2(net448),
    .B1(_0295_),
    .Y(_0296_));
 sky130_fd_sc_hd__nor2_1 _0718_ (.A(net478),
    .B(net752),
    .Y(_0062_));
 sky130_fd_sc_hd__o221a_1 _0719_ (.A1(net1083),
    .A2(net469),
    .B1(_0237_),
    .B2(net673),
    .C1(net446),
    .X(_0297_));
 sky130_fd_sc_hd__a21oi_1 _0720_ (.A1(net784),
    .A2(net448),
    .B1(_0297_),
    .Y(_0298_));
 sky130_fd_sc_hd__nor2_1 _0721_ (.A(net478),
    .B(net785),
    .Y(_0063_));
 sky130_fd_sc_hd__o221a_1 _0722_ (.A1(net1077),
    .A2(net469),
    .B1(_0237_),
    .B2(net722),
    .C1(net446),
    .X(_0299_));
 sky130_fd_sc_hd__a21oi_1 _0723_ (.A1(net739),
    .A2(net448),
    .B1(_0299_),
    .Y(_0300_));
 sky130_fd_sc_hd__nor2_1 _0724_ (.A(net478),
    .B(net740),
    .Y(_0064_));
 sky130_fd_sc_hd__o221a_1 _0725_ (.A1(net1058),
    .A2(net469),
    .B1(net467),
    .B2(net654),
    .C1(net446),
    .X(_0301_));
 sky130_fd_sc_hd__a21oi_1 _0726_ (.A1(net798),
    .A2(net448),
    .B1(_0301_),
    .Y(_0302_));
 sky130_fd_sc_hd__nor2_1 _0727_ (.A(net478),
    .B(net799),
    .Y(_0065_));
 sky130_fd_sc_hd__o221a_1 _0728_ (.A1(net1042),
    .A2(net469),
    .B1(net467),
    .B2(net733),
    .C1(net445),
    .X(_0303_));
 sky130_fd_sc_hd__a21oi_1 _0729_ (.A1(net745),
    .A2(net448),
    .B1(_0303_),
    .Y(_0304_));
 sky130_fd_sc_hd__nor2_1 _0730_ (.A(net478),
    .B(net746),
    .Y(_0066_));
 sky130_fd_sc_hd__o221a_1 _0731_ (.A1(net1089),
    .A2(net469),
    .B1(net467),
    .B2(net832),
    .C1(net445),
    .X(_0305_));
 sky130_fd_sc_hd__a21oi_1 _0732_ (.A1(net769),
    .A2(net448),
    .B1(_0305_),
    .Y(_0306_));
 sky130_fd_sc_hd__nor2_1 _0733_ (.A(net478),
    .B(net770),
    .Y(_0067_));
 sky130_fd_sc_hd__o221a_1 _0734_ (.A1(net1055),
    .A2(net469),
    .B1(net467),
    .B2(net849),
    .C1(net445),
    .X(_0307_));
 sky130_fd_sc_hd__a21oi_1 _0735_ (.A1(net736),
    .A2(net448),
    .B1(_0307_),
    .Y(_0308_));
 sky130_fd_sc_hd__nor2_1 _0736_ (.A(net478),
    .B(net737),
    .Y(_0068_));
 sky130_fd_sc_hd__and2_1 _0737_ (.A(net604),
    .B(net474),
    .X(_0069_));
 sky130_fd_sc_hd__nor2_4 _0738_ (.A(net1180),
    .B(net467),
    .Y(_0309_));
 sky130_fd_sc_hd__or2_1 _0739_ (.A(net1180),
    .B(net467),
    .X(_0310_));
 sky130_fd_sc_hd__nand2_1 _0740_ (.A(net814),
    .B(net438),
    .Y(_0311_));
 sky130_fd_sc_hd__o211a_1 _0741_ (.A1(net845),
    .A2(net438),
    .B1(net815),
    .C1(net473),
    .X(_0070_));
 sky130_fd_sc_hd__nand2_1 _0742_ (.A(net814),
    .B(net860),
    .Y(_0312_));
 sky130_fd_sc_hd__or2_1 _0743_ (.A(net814),
    .B(net860),
    .X(_0313_));
 sky130_fd_sc_hd__a21o_1 _0744_ (.A1(net861),
    .A2(_0313_),
    .B1(_0309_),
    .X(_0314_));
 sky130_fd_sc_hd__o211a_1 _0745_ (.A1(net854),
    .A2(net438),
    .B1(net862),
    .C1(net473),
    .X(_0071_));
 sky130_fd_sc_hd__xnor2_1 _0746_ (.A(net888),
    .B(net861),
    .Y(_0315_));
 sky130_fd_sc_hd__or2_1 _0747_ (.A(net885),
    .B(net438),
    .X(_0316_));
 sky130_fd_sc_hd__o211a_1 _0748_ (.A1(_0309_),
    .A2(net889),
    .B1(_0316_),
    .C1(net473),
    .X(_0072_));
 sky130_fd_sc_hd__and4_2 _0749_ (.A(net814),
    .B(net860),
    .C(net1132),
    .D(net1015),
    .X(_0317_));
 sky130_fd_sc_hd__a31oi_1 _0750_ (.A1(net814),
    .A2(net860),
    .A3(net888),
    .B1(net1015),
    .Y(_0318_));
 sky130_fd_sc_hd__o21ai_1 _0751_ (.A1(_0317_),
    .A2(net1016),
    .B1(net440),
    .Y(_0319_));
 sky130_fd_sc_hd__o211a_1 _0752_ (.A1(net697),
    .A2(net438),
    .B1(net1017),
    .C1(net476),
    .X(_0073_));
 sky130_fd_sc_hd__xnor2_1 _0753_ (.A(net1045),
    .B(_0317_),
    .Y(_0320_));
 sky130_fd_sc_hd__nand2_1 _0754_ (.A(net437),
    .B(net1046),
    .Y(_0321_));
 sky130_fd_sc_hd__o211a_1 _0755_ (.A1(net817),
    .A2(net437),
    .B1(_0321_),
    .C1(net472),
    .X(_0074_));
 sky130_fd_sc_hd__a21oi_1 _0756_ (.A1(\wb_counter[4] ),
    .A2(_0317_),
    .B1(net801),
    .Y(_0322_));
 sky130_fd_sc_hd__and3_1 _0757_ (.A(net1045),
    .B(net801),
    .C(_0317_),
    .X(_0323_));
 sky130_fd_sc_hd__o21ai_1 _0758_ (.A1(net802),
    .A2(_0323_),
    .B1(net437),
    .Y(_0324_));
 sky130_fd_sc_hd__o211a_1 _0759_ (.A1(net793),
    .A2(net437),
    .B1(net803),
    .C1(net472),
    .X(_0075_));
 sky130_fd_sc_hd__or2_1 _0760_ (.A(net866),
    .B(_0323_),
    .X(_0325_));
 sky130_fd_sc_hd__nand2_1 _0761_ (.A(net866),
    .B(_0323_),
    .Y(_0326_));
 sky130_fd_sc_hd__a21o_1 _0762_ (.A1(_0325_),
    .A2(net867),
    .B1(_0309_),
    .X(_0327_));
 sky130_fd_sc_hd__o211a_1 _0763_ (.A1(net864),
    .A2(net437),
    .B1(net868),
    .C1(net471),
    .X(_0076_));
 sky130_fd_sc_hd__a21oi_1 _0764_ (.A1(\wb_counter[6] ),
    .A2(_0323_),
    .B1(net677),
    .Y(_0328_));
 sky130_fd_sc_hd__and4_1 _0765_ (.A(net1045),
    .B(net801),
    .C(net866),
    .D(net677),
    .X(_0329_));
 sky130_fd_sc_hd__and2_1 _0766_ (.A(_0317_),
    .B(_0329_),
    .X(_0330_));
 sky130_fd_sc_hd__o21ai_1 _0767_ (.A1(net678),
    .A2(_0330_),
    .B1(net437),
    .Y(_0331_));
 sky130_fd_sc_hd__o211a_1 _0768_ (.A1(net666),
    .A2(net437),
    .B1(net679),
    .C1(net471),
    .X(_0077_));
 sky130_fd_sc_hd__nor2_1 _0769_ (.A(net1038),
    .B(_0330_),
    .Y(_0332_));
 sky130_fd_sc_hd__and3_1 _0770_ (.A(net1038),
    .B(_0317_),
    .C(_0329_),
    .X(_0333_));
 sky130_fd_sc_hd__o21ai_1 _0771_ (.A1(net1039),
    .A2(_0333_),
    .B1(net437),
    .Y(_0334_));
 sky130_fd_sc_hd__o211a_1 _0772_ (.A1(net664),
    .A2(net437),
    .B1(net1040),
    .C1(net471),
    .X(_0078_));
 sky130_fd_sc_hd__nor2_1 _0773_ (.A(net633),
    .B(_0333_),
    .Y(_0335_));
 sky130_fd_sc_hd__and2_1 _0774_ (.A(net633),
    .B(_0333_),
    .X(_0336_));
 sky130_fd_sc_hd__o21ai_1 _0775_ (.A1(net634),
    .A2(_0336_),
    .B1(net437),
    .Y(_0337_));
 sky130_fd_sc_hd__o211a_1 _0776_ (.A1(net631),
    .A2(net437),
    .B1(net635),
    .C1(net471),
    .X(_0079_));
 sky130_fd_sc_hd__xnor2_1 _0777_ (.A(net1023),
    .B(_0336_),
    .Y(_0338_));
 sky130_fd_sc_hd__nand2_1 _0778_ (.A(net437),
    .B(net1024),
    .Y(_0339_));
 sky130_fd_sc_hd__o211a_1 _0779_ (.A1(net645),
    .A2(net437),
    .B1(net1025),
    .C1(net471),
    .X(_0080_));
 sky130_fd_sc_hd__a21oi_1 _0780_ (.A1(\wb_counter[10] ),
    .A2(_0336_),
    .B1(net658),
    .Y(_0340_));
 sky130_fd_sc_hd__and4_1 _0781_ (.A(net1038),
    .B(net633),
    .C(net1023),
    .D(net658),
    .X(_0341_));
 sky130_fd_sc_hd__and3_1 _0782_ (.A(_0317_),
    .B(_0329_),
    .C(_0341_),
    .X(_0342_));
 sky130_fd_sc_hd__o21ai_1 _0783_ (.A1(net659),
    .A2(_0342_),
    .B1(net437),
    .Y(_0343_));
 sky130_fd_sc_hd__o211a_1 _0784_ (.A1(net650),
    .A2(net437),
    .B1(net660),
    .C1(net471),
    .X(_0081_));
 sky130_fd_sc_hd__nor2_1 _0785_ (.A(net1070),
    .B(_0342_),
    .Y(_0344_));
 sky130_fd_sc_hd__and2_1 _0786_ (.A(net1070),
    .B(_0342_),
    .X(_0345_));
 sky130_fd_sc_hd__o21ai_1 _0787_ (.A1(net1071),
    .A2(_0345_),
    .B1(net438),
    .Y(_0346_));
 sky130_fd_sc_hd__o211a_1 _0788_ (.A1(net626),
    .A2(net437),
    .B1(net1072),
    .C1(net471),
    .X(_0082_));
 sky130_fd_sc_hd__nor2_1 _0789_ (.A(net622),
    .B(_0345_),
    .Y(_0347_));
 sky130_fd_sc_hd__and3_1 _0790_ (.A(net1070),
    .B(net622),
    .C(_0342_),
    .X(_0348_));
 sky130_fd_sc_hd__o21ai_1 _0791_ (.A1(net623),
    .A2(_0348_),
    .B1(net438),
    .Y(_0349_));
 sky130_fd_sc_hd__o211a_1 _0792_ (.A1(net577),
    .A2(net438),
    .B1(net624),
    .C1(net473),
    .X(_0083_));
 sky130_fd_sc_hd__nor2_1 _0793_ (.A(net1034),
    .B(_0348_),
    .Y(_0350_));
 sky130_fd_sc_hd__and2_1 _0794_ (.A(net1034),
    .B(_0348_),
    .X(_0351_));
 sky130_fd_sc_hd__o21ai_1 _0795_ (.A1(net1035),
    .A2(_0351_),
    .B1(net438),
    .Y(_0352_));
 sky130_fd_sc_hd__o211a_1 _0796_ (.A1(net616),
    .A2(net438),
    .B1(net1036),
    .C1(net473),
    .X(_0084_));
 sky130_fd_sc_hd__nor2_1 _0797_ (.A(net1019),
    .B(_0351_),
    .Y(_0353_));
 sky130_fd_sc_hd__and4_1 _0798_ (.A(\wb_counter[12] ),
    .B(net622),
    .C(net1034),
    .D(net1019),
    .X(_0354_));
 sky130_fd_sc_hd__and4_2 _0799_ (.A(_0317_),
    .B(_0329_),
    .C(_0341_),
    .D(_0354_),
    .X(_0355_));
 sky130_fd_sc_hd__o21ai_1 _0800_ (.A1(net1020),
    .A2(_0355_),
    .B1(net438),
    .Y(_0356_));
 sky130_fd_sc_hd__o211a_1 _0801_ (.A1(net614),
    .A2(net438),
    .B1(net1021),
    .C1(net473),
    .X(_0085_));
 sky130_fd_sc_hd__xnor2_1 _0802_ (.A(net610),
    .B(_0355_),
    .Y(_0357_));
 sky130_fd_sc_hd__nand2_1 _0803_ (.A(net438),
    .B(net611),
    .Y(_0358_));
 sky130_fd_sc_hd__o211a_1 _0804_ (.A1(net1138),
    .A2(net438),
    .B1(net612),
    .C1(net473),
    .X(_0086_));
 sky130_fd_sc_hd__a21oi_1 _0805_ (.A1(net610),
    .A2(_0355_),
    .B1(net706),
    .Y(_0359_));
 sky130_fd_sc_hd__and2_1 _0806_ (.A(net610),
    .B(net706),
    .X(_0360_));
 sky130_fd_sc_hd__and2_1 _0807_ (.A(_0355_),
    .B(_0360_),
    .X(_0361_));
 sky130_fd_sc_hd__o21ai_1 _0808_ (.A1(net707),
    .A2(_0361_),
    .B1(net439),
    .Y(_0362_));
 sky130_fd_sc_hd__o211a_1 _0809_ (.A1(net702),
    .A2(net438),
    .B1(net708),
    .C1(net473),
    .X(_0087_));
 sky130_fd_sc_hd__nor2_1 _0810_ (.A(net685),
    .B(_0361_),
    .Y(_0363_));
 sky130_fd_sc_hd__and3_1 _0811_ (.A(net685),
    .B(_0355_),
    .C(_0360_),
    .X(_0364_));
 sky130_fd_sc_hd__o21ai_1 _0812_ (.A1(net686),
    .A2(_0364_),
    .B1(net439),
    .Y(_0365_));
 sky130_fd_sc_hd__o211a_1 _0813_ (.A1(net681),
    .A2(net439),
    .B1(net687),
    .C1(net475),
    .X(_0088_));
 sky130_fd_sc_hd__and2_1 _0814_ (.A(net685),
    .B(net1166),
    .X(_0366_));
 sky130_fd_sc_hd__nand2_1 _0815_ (.A(_0361_),
    .B(_0366_),
    .Y(_0367_));
 sky130_fd_sc_hd__o211a_1 _0816_ (.A1(net1166),
    .A2(_0364_),
    .B1(_0367_),
    .C1(net439),
    .X(_0368_));
 sky130_fd_sc_hd__a21oi_1 _0817_ (.A1(net714),
    .A2(_0309_),
    .B1(_0368_),
    .Y(_0369_));
 sky130_fd_sc_hd__nor2_1 _0818_ (.A(net478),
    .B(net715),
    .Y(_0089_));
 sky130_fd_sc_hd__and4_1 _0819_ (.A(net710),
    .B(_0355_),
    .C(_0360_),
    .D(_0366_),
    .X(_0370_));
 sky130_fd_sc_hd__xor2_1 _0820_ (.A(net710),
    .B(_0367_),
    .X(_0371_));
 sky130_fd_sc_hd__nand2_1 _0821_ (.A(net439),
    .B(net711),
    .Y(_0372_));
 sky130_fd_sc_hd__o211a_1 _0822_ (.A1(net704),
    .A2(net439),
    .B1(net712),
    .C1(net475),
    .X(_0090_));
 sky130_fd_sc_hd__nor2_1 _0823_ (.A(net1051),
    .B(_0370_),
    .Y(_0373_));
 sky130_fd_sc_hd__and2_1 _0824_ (.A(net1051),
    .B(_0370_),
    .X(_0374_));
 sky130_fd_sc_hd__o21ai_1 _0825_ (.A1(net1052),
    .A2(_0374_),
    .B1(net439),
    .Y(_0375_));
 sky130_fd_sc_hd__o211a_1 _0826_ (.A1(net692),
    .A2(net439),
    .B1(net1053),
    .C1(net475),
    .X(_0091_));
 sky130_fd_sc_hd__nor2_1 _0827_ (.A(net1047),
    .B(_0374_),
    .Y(_0376_));
 sky130_fd_sc_hd__and3_1 _0828_ (.A(\wb_counter[21] ),
    .B(net1047),
    .C(_0370_),
    .X(_0377_));
 sky130_fd_sc_hd__o21ai_1 _0829_ (.A1(net1048),
    .A2(_0377_),
    .B1(net439),
    .Y(_0378_));
 sky130_fd_sc_hd__o211a_1 _0830_ (.A1(net683),
    .A2(net439),
    .B1(net1049),
    .C1(net475),
    .X(_0092_));
 sky130_fd_sc_hd__nor2_1 _0831_ (.A(net1027),
    .B(_0377_),
    .Y(_0379_));
 sky130_fd_sc_hd__and4_2 _0832_ (.A(net1051),
    .B(net1047),
    .C(net1027),
    .D(_0370_),
    .X(_0380_));
 sky130_fd_sc_hd__o21ai_1 _0833_ (.A1(net1028),
    .A2(_0380_),
    .B1(net439),
    .Y(_0381_));
 sky130_fd_sc_hd__o211a_1 _0834_ (.A1(net717),
    .A2(net439),
    .B1(net1029),
    .C1(net474),
    .X(_0093_));
 sky130_fd_sc_hd__or2_1 _0835_ (.A(net841),
    .B(_0380_),
    .X(_0382_));
 sky130_fd_sc_hd__nand2_1 _0836_ (.A(net841),
    .B(_0380_),
    .Y(_0383_));
 sky130_fd_sc_hd__a21o_1 _0837_ (.A1(_0382_),
    .A2(net842),
    .B1(_0309_),
    .X(_0384_));
 sky130_fd_sc_hd__o211a_1 _0838_ (.A1(net725),
    .A2(net439),
    .B1(_0384_),
    .C1(net474),
    .X(_0094_));
 sky130_fd_sc_hd__xnor2_1 _0839_ (.A(net356),
    .B(net842),
    .Y(_0385_));
 sky130_fd_sc_hd__or2_1 _0840_ (.A(net643),
    .B(net439),
    .X(_0386_));
 sky130_fd_sc_hd__o211a_1 _0841_ (.A1(_0309_),
    .A2(net843),
    .B1(_0386_),
    .C1(net476),
    .X(_0095_));
 sky130_fd_sc_hd__and4_2 _0842_ (.A(net841),
    .B(net356),
    .C(net673),
    .D(_0380_),
    .X(_0387_));
 sky130_fd_sc_hd__a31oi_1 _0843_ (.A1(\wb_counter[24] ),
    .A2(net356),
    .A3(_0380_),
    .B1(net673),
    .Y(_0388_));
 sky130_fd_sc_hd__o21ai_1 _0844_ (.A1(_0387_),
    .A2(net674),
    .B1(net439),
    .Y(_0389_));
 sky130_fd_sc_hd__o211a_1 _0845_ (.A1(net668),
    .A2(net439),
    .B1(net675),
    .C1(net474),
    .X(_0096_));
 sky130_fd_sc_hd__xor2_1 _0846_ (.A(net722),
    .B(_0387_),
    .X(_0390_));
 sky130_fd_sc_hd__or2_1 _0847_ (.A(net606),
    .B(net440),
    .X(_0391_));
 sky130_fd_sc_hd__o211a_1 _0848_ (.A1(_0309_),
    .A2(net723),
    .B1(_0391_),
    .C1(net474),
    .X(_0097_));
 sky130_fd_sc_hd__and3_1 _0849_ (.A(net722),
    .B(net654),
    .C(_0387_),
    .X(_0392_));
 sky130_fd_sc_hd__a21oi_1 _0850_ (.A1(\wb_counter[27] ),
    .A2(_0387_),
    .B1(net654),
    .Y(_0393_));
 sky130_fd_sc_hd__o21ai_1 _0851_ (.A1(_0392_),
    .A2(net655),
    .B1(net440),
    .Y(_0394_));
 sky130_fd_sc_hd__o211a_1 _0852_ (.A1(net652),
    .A2(net440),
    .B1(net656),
    .C1(net474),
    .X(_0098_));
 sky130_fd_sc_hd__and4_1 _0853_ (.A(net722),
    .B(net654),
    .C(net733),
    .D(_0387_),
    .X(_0395_));
 sky130_fd_sc_hd__xor2_1 _0854_ (.A(net733),
    .B(_0392_),
    .X(_0104_));
 sky130_fd_sc_hd__or2_1 _0855_ (.A(net618),
    .B(net440),
    .X(_0105_));
 sky130_fd_sc_hd__o211a_1 _0856_ (.A1(_0309_),
    .A2(net734),
    .B1(_0105_),
    .C1(net474),
    .X(_0099_));
 sky130_fd_sc_hd__xor2_1 _0857_ (.A(net832),
    .B(_0395_),
    .X(_0106_));
 sky130_fd_sc_hd__or2_1 _0858_ (.A(net620),
    .B(net440),
    .X(_0107_));
 sky130_fd_sc_hd__o211a_1 _0859_ (.A1(_0309_),
    .A2(net833),
    .B1(_0107_),
    .C1(net474),
    .X(_0100_));
 sky130_fd_sc_hd__and3b_1 _0860_ (.A_N(net849),
    .B(_0395_),
    .C(net832),
    .X(_0108_));
 sky130_fd_sc_hd__a21boi_1 _0861_ (.A1(net832),
    .A2(_0395_),
    .B1_N(net849),
    .Y(_0109_));
 sky130_fd_sc_hd__or2_1 _0862_ (.A(net662),
    .B(net440),
    .X(_0110_));
 sky130_fd_sc_hd__o311a_1 _0863_ (.A1(_0309_),
    .A2(_0108_),
    .A3(net850),
    .B1(_0110_),
    .C1(net476),
    .X(_0101_));
 sky130_fd_sc_hd__or3_1 _0864_ (.A(net845),
    .B(net872),
    .C(net857),
    .X(_0111_));
 sky130_fd_sc_hd__o211a_1 _0865_ (.A1(net847),
    .A2(net873),
    .B1(net1176),
    .C1(net475),
    .X(_0102_));
 sky130_fd_sc_hd__mux2_1 _0866_ (.A0(net556),
    .A1(net854),
    .S(net873),
    .X(_0112_));
 sky130_fd_sc_hd__or2_1 _0867_ (.A(net478),
    .B(net874),
    .X(_0103_));
 sky130_fd_sc_hd__dfxtp_1 _0868_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(net605),
    .Q(wb_feedback_delay));
 sky130_fd_sc_hd__dfxtp_2 _0869_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(net846),
    .Q(net258));
 sky130_fd_sc_hd__dfxtp_2 _0870_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(net855),
    .Q(net269));
 sky130_fd_sc_hd__dfxtp_2 _0871_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(net853),
    .Q(net280));
 sky130_fd_sc_hd__dfxtp_2 _0872_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(net701),
    .Q(net283));
 sky130_fd_sc_hd__dfxtp_2 _0873_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(net821),
    .Q(net284));
 sky130_fd_sc_hd__dfxtp_2 _0874_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(net794),
    .Q(net285));
 sky130_fd_sc_hd__dfxtp_2 _0875_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(net865),
    .Q(net286));
 sky130_fd_sc_hd__dfxtp_2 _0876_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(net667),
    .Q(net287));
 sky130_fd_sc_hd__dfxtp_2 _0877_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(net672),
    .Q(net288));
 sky130_fd_sc_hd__dfxtp_2 _0878_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(net632),
    .Q(net289));
 sky130_fd_sc_hd__dfxtp_2 _0879_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(net649),
    .Q(net259));
 sky130_fd_sc_hd__dfxtp_2 _0880_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(net651),
    .Q(net260));
 sky130_fd_sc_hd__dfxtp_2 _0881_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(net642),
    .Q(net261));
 sky130_fd_sc_hd__dfxtp_2 _0882_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(net1100),
    .Q(net262));
 sky130_fd_sc_hd__dfxtp_2 _0883_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(net630),
    .Q(net263));
 sky130_fd_sc_hd__dfxtp_2 _0884_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(net639),
    .Q(net264));
 sky130_fd_sc_hd__dfxtp_2 _0885_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(net609),
    .Q(net265));
 sky130_fd_sc_hd__dfxtp_2 _0886_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(net703),
    .Q(net266));
 sky130_fd_sc_hd__dfxtp_2 _0887_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(net682),
    .Q(net267));
 sky130_fd_sc_hd__dfxtp_2 _0888_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(net797),
    .Q(net268));
 sky130_fd_sc_hd__dfxtp_2 _0889_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(net705),
    .Q(net270));
 sky130_fd_sc_hd__dfxtp_2 _0890_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(net696),
    .Q(net271));
 sky130_fd_sc_hd__dfxtp_2 _0891_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(net691),
    .Q(net272));
 sky130_fd_sc_hd__dfxtp_2 _0892_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(net721),
    .Q(net273));
 sky130_fd_sc_hd__dfxtp_2 _0893_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(net729),
    .Q(net274));
 sky130_fd_sc_hd__dfxtp_2 _0894_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(net644),
    .Q(net275));
 sky130_fd_sc_hd__dfxtp_2 _0895_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(net669),
    .Q(net276));
 sky130_fd_sc_hd__dfxtp_2 _0896_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(net607),
    .Q(net277));
 sky130_fd_sc_hd__dfxtp_2 _0897_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(net653),
    .Q(net278));
 sky130_fd_sc_hd__dfxtp_2 _0898_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(net619),
    .Q(net279));
 sky130_fd_sc_hd__dfxtp_2 _0899_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(net621),
    .Q(net281));
 sky130_fd_sc_hd__dfxtp_2 _0900_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(net663),
    .Q(net282));
 sky130_fd_sc_hd__dfxtp_1 _0901_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(net887),
    .Q(\design_select[0] ));
 sky130_fd_sc_hd__dfxtp_1 _0902_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(net859),
    .Q(\design_select[1] ));
 sky130_fd_sc_hd__dfxtp_1 _0903_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(net883),
    .Q(\design_select[2] ));
 sky130_fd_sc_hd__dfxtp_1 _0904_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(net879),
    .Q(\design_select[3] ));
 sky130_fd_sc_hd__dfxtp_1 _0905_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(net831),
    .Q(net405));
 sky130_fd_sc_hd__dfxtp_1 _0906_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(net829),
    .Q(net416));
 sky130_fd_sc_hd__dfxtp_1 _0907_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(net827),
    .Q(net427));
 sky130_fd_sc_hd__dfxtp_1 _0908_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(net825),
    .Q(net430));
 sky130_fd_sc_hd__dfxtp_1 _0909_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(net836),
    .Q(net431));
 sky130_fd_sc_hd__dfxtp_1 _0910_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(net838),
    .Q(net432));
 sky130_fd_sc_hd__dfxtp_1 _0911_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(net840),
    .Q(net433));
 sky130_fd_sc_hd__dfxtp_1 _0912_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(net823),
    .Q(net434));
 sky130_fd_sc_hd__dfxtp_1 _0913_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(net792),
    .Q(net435));
 sky130_fd_sc_hd__dfxtp_1 _0914_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(net789),
    .Q(net436));
 sky130_fd_sc_hd__dfxtp_1 _0915_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(net813),
    .Q(net406));
 sky130_fd_sc_hd__dfxtp_1 _0916_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(net732),
    .Q(net407));
 sky130_fd_sc_hd__dfxtp_1 _0917_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(net756),
    .Q(net408));
 sky130_fd_sc_hd__dfxtp_1 _0918_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(net759),
    .Q(net409));
 sky130_fd_sc_hd__dfxtp_1 _0919_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(net810),
    .Q(net410));
 sky130_fd_sc_hd__dfxtp_1 _0920_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(net768),
    .Q(net411));
 sky130_fd_sc_hd__dfxtp_1 _0921_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(net807),
    .Q(net412));
 sky130_fd_sc_hd__dfxtp_1 _0922_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(net783),
    .Q(net413));
 sky130_fd_sc_hd__dfxtp_1 _0923_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(net750),
    .Q(net414));
 sky130_fd_sc_hd__dfxtp_1 _0924_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(net762),
    .Q(net415));
 sky130_fd_sc_hd__dfxtp_1 _0925_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(net777),
    .Q(net417));
 sky130_fd_sc_hd__dfxtp_1 _0926_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(net765),
    .Q(net418));
 sky130_fd_sc_hd__dfxtp_1 _0927_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(net780),
    .Q(net419));
 sky130_fd_sc_hd__dfxtp_1 _0928_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(net744),
    .Q(net420));
 sky130_fd_sc_hd__dfxtp_1 _0929_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(net774),
    .Q(net421));
 sky130_fd_sc_hd__dfxtp_1 _0930_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(net753),
    .Q(net422));
 sky130_fd_sc_hd__dfxtp_1 _0931_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(net786),
    .Q(net423));
 sky130_fd_sc_hd__dfxtp_1 _0932_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(net741),
    .Q(net424));
 sky130_fd_sc_hd__dfxtp_1 _0933_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(net800),
    .Q(net425));
 sky130_fd_sc_hd__dfxtp_1 _0934_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(net747),
    .Q(net426));
 sky130_fd_sc_hd__dfxtp_1 _0935_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(net771),
    .Q(net428));
 sky130_fd_sc_hd__dfxtp_1 _0936_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(net738),
    .Q(net429));
 sky130_fd_sc_hd__dfxtp_1 _0937_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(net588),
    .Q(net404));
 sky130_fd_sc_hd__dfxtp_1 _0938_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(net816),
    .Q(\wb_counter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _0939_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(net863),
    .Q(\wb_counter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _0940_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(net890),
    .Q(\wb_counter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _0941_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(net698),
    .Q(\wb_counter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _0942_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(net818),
    .Q(\wb_counter[4] ));
 sky130_fd_sc_hd__dfxtp_1 _0943_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(net804),
    .Q(\wb_counter[5] ));
 sky130_fd_sc_hd__dfxtp_1 _0944_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(net869),
    .Q(\wb_counter[6] ));
 sky130_fd_sc_hd__dfxtp_1 _0945_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(net680),
    .Q(\wb_counter[7] ));
 sky130_fd_sc_hd__dfxtp_1 _0946_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(net665),
    .Q(\wb_counter[8] ));
 sky130_fd_sc_hd__dfxtp_1 _0947_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(net636),
    .Q(\wb_counter[9] ));
 sky130_fd_sc_hd__dfxtp_1 _0948_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(net646),
    .Q(\wb_counter[10] ));
 sky130_fd_sc_hd__dfxtp_1 _0949_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(net661),
    .Q(\wb_counter[11] ));
 sky130_fd_sc_hd__dfxtp_1 _0950_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(net627),
    .Q(\wb_counter[12] ));
 sky130_fd_sc_hd__dfxtp_1 _0951_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(net625),
    .Q(\wb_counter[13] ));
 sky130_fd_sc_hd__dfxtp_1 _0952_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(net617),
    .Q(\wb_counter[14] ));
 sky130_fd_sc_hd__dfxtp_1 _0953_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(net615),
    .Q(\wb_counter[15] ));
 sky130_fd_sc_hd__dfxtp_1 _0954_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(net613),
    .Q(\wb_counter[16] ));
 sky130_fd_sc_hd__dfxtp_1 _0955_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(net709),
    .Q(\wb_counter[17] ));
 sky130_fd_sc_hd__dfxtp_1 _0956_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(net688),
    .Q(\wb_counter[18] ));
 sky130_fd_sc_hd__dfxtp_1 _0957_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(net716),
    .Q(\wb_counter[19] ));
 sky130_fd_sc_hd__dfxtp_1 _0958_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(net713),
    .Q(\wb_counter[20] ));
 sky130_fd_sc_hd__dfxtp_1 _0959_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(net693),
    .Q(\wb_counter[21] ));
 sky130_fd_sc_hd__dfxtp_1 _0960_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(net684),
    .Q(\wb_counter[22] ));
 sky130_fd_sc_hd__dfxtp_1 _0961_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(net718),
    .Q(\wb_counter[23] ));
 sky130_fd_sc_hd__dfxtp_1 _0962_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(net726),
    .Q(\wb_counter[24] ));
 sky130_fd_sc_hd__dfxtp_4 _0963_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(net844),
    .Q(net356));
 sky130_fd_sc_hd__dfxtp_1 _0964_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(net676),
    .Q(\wb_counter[26] ));
 sky130_fd_sc_hd__dfxtp_1 _0965_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(net724),
    .Q(\wb_counter[27] ));
 sky130_fd_sc_hd__dfxtp_1 _0966_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(net657),
    .Q(\wb_counter[28] ));
 sky130_fd_sc_hd__dfxtp_1 _0967_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(net735),
    .Q(\wb_counter[29] ));
 sky130_fd_sc_hd__dfxtp_1 _0968_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(net834),
    .Q(\wb_counter[30] ));
 sky130_fd_sc_hd__dfxtp_1 _0969_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(net851),
    .Q(\wb_counter[31] ));
 sky130_fd_sc_hd__dfxtp_1 _0970_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(net848),
    .Q(wb_override_act));
 sky130_fd_sc_hd__dfxtp_1 _0971_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(net875),
    .Q(wb_rst_override));
 sky130_fd_sc_hd__dfxtp_1 _0972_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(net499),
    .Q(\wbs_dat_delaybuff[0] ));
 sky130_fd_sc_hd__dfxtp_1 _0973_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(net495),
    .Q(\wbs_dat_delaybuff[1] ));
 sky130_fd_sc_hd__dfxtp_1 _0974_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(net497),
    .Q(\wbs_dat_delaybuff[2] ));
 sky130_fd_sc_hd__dfxtp_1 _0975_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(net505),
    .Q(\wbs_dat_delaybuff[3] ));
 sky130_fd_sc_hd__dfxtp_1 _0976_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(net493),
    .Q(\wbs_dat_delaybuff[4] ));
 sky130_fd_sc_hd__dfxtp_1 _0977_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(net503),
    .Q(\wbs_dat_delaybuff[5] ));
 sky130_fd_sc_hd__dfxtp_1 _0978_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(net501),
    .Q(\wbs_dat_delaybuff[6] ));
 sky130_fd_sc_hd__dfxtp_1 _0979_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(net507),
    .Q(\wbs_dat_delaybuff[7] ));
 sky130_fd_sc_hd__dfxtp_1 _0980_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(net513),
    .Q(\wbs_dat_delaybuff[8] ));
 sky130_fd_sc_hd__dfxtp_1 _0981_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(net519),
    .Q(\wbs_dat_delaybuff[9] ));
 sky130_fd_sc_hd__dfxtp_1 _0982_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(net515),
    .Q(\wbs_dat_delaybuff[10] ));
 sky130_fd_sc_hd__dfxtp_1 _0983_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(net511),
    .Q(\wbs_dat_delaybuff[11] ));
 sky130_fd_sc_hd__dfxtp_1 _0984_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(net509),
    .Q(\wbs_dat_delaybuff[12] ));
 sky130_fd_sc_hd__dfxtp_1 _0985_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(net529),
    .Q(\wbs_dat_delaybuff[13] ));
 sky130_fd_sc_hd__dfxtp_1 _0986_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(net523),
    .Q(\wbs_dat_delaybuff[14] ));
 sky130_fd_sc_hd__dfxtp_1 _0987_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(net525),
    .Q(\wbs_dat_delaybuff[15] ));
 sky130_fd_sc_hd__dfxtp_1 _0988_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(net521),
    .Q(\wbs_dat_delaybuff[16] ));
 sky130_fd_sc_hd__dfxtp_1 _0989_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(net545),
    .Q(\wbs_dat_delaybuff[17] ));
 sky130_fd_sc_hd__dfxtp_1 _0990_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(net541),
    .Q(\wbs_dat_delaybuff[18] ));
 sky130_fd_sc_hd__dfxtp_1 _0991_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(net517),
    .Q(\wbs_dat_delaybuff[19] ));
 sky130_fd_sc_hd__dfxtp_1 _0992_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(net533),
    .Q(\wbs_dat_delaybuff[20] ));
 sky130_fd_sc_hd__dfxtp_1 _0993_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(net535),
    .Q(\wbs_dat_delaybuff[21] ));
 sky130_fd_sc_hd__dfxtp_1 _0994_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(net547),
    .Q(\wbs_dat_delaybuff[22] ));
 sky130_fd_sc_hd__dfxtp_1 _0995_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(net527),
    .Q(\wbs_dat_delaybuff[23] ));
 sky130_fd_sc_hd__dfxtp_1 _0996_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(net537),
    .Q(\wbs_dat_delaybuff[24] ));
 sky130_fd_sc_hd__dfxtp_1 _0997_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(net549),
    .Q(\wbs_dat_delaybuff[25] ));
 sky130_fd_sc_hd__dfxtp_1 _0998_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(net553),
    .Q(\wbs_dat_delaybuff[26] ));
 sky130_fd_sc_hd__dfxtp_1 _0999_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(net555),
    .Q(\wbs_dat_delaybuff[27] ));
 sky130_fd_sc_hd__dfxtp_1 _1000_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(net551),
    .Q(\wbs_dat_delaybuff[28] ));
 sky130_fd_sc_hd__dfxtp_1 _1001_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(net543),
    .Q(\wbs_dat_delaybuff[29] ));
 sky130_fd_sc_hd__dfxtp_1 _1002_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(net539),
    .Q(\wbs_dat_delaybuff[30] ));
 sky130_fd_sc_hd__dfxtp_1 _1003_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(net531),
    .Q(\wbs_dat_delaybuff[31] ));
 sky130_fd_sc_hd__dfxtp_1 _1004_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(net485),
    .Q(\wbs_adr_delaybuff[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1005_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(net491),
    .Q(\wbs_adr_delaybuff[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1006_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(net489),
    .Q(\wbs_adr_delaybuff[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1007_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(net487),
    .Q(\wbs_adr_delaybuff[3] ));
 sky130_fd_sc_hd__clkbuf_1 _1013_ (.A(net568),
    .X(net373));
 sky130_fd_sc_hd__buf_1 _1014_ (.A(net575),
    .X(net384));
 sky130_fd_sc_hd__buf_1 _1015_ (.A(net561),
    .X(net395));
 sky130_fd_sc_hd__clkbuf_2 _1016_ (.A(net321),
    .X(net396));
 sky130_fd_sc_hd__clkbuf_2 _1017_ (.A(net322),
    .X(net397));
 sky130_fd_sc_hd__clkbuf_2 _1018_ (.A(net582),
    .X(net398));
 sky130_fd_sc_hd__clkbuf_2 _1019_ (.A(net324),
    .X(net399));
 sky130_fd_sc_hd__clkbuf_2 _1020_ (.A(net325),
    .X(net400));
 sky130_fd_sc_hd__clkbuf_2 _1021_ (.A(net290),
    .X(net363));
 sky130_fd_sc_hd__clkbuf_2 _1022_ (.A(net291),
    .X(net364));
 sky130_fd_sc_hd__clkbuf_2 _1023_ (.A(net292),
    .X(net365));
 sky130_fd_sc_hd__clkbuf_2 _1024_ (.A(net293),
    .X(net366));
 sky130_fd_sc_hd__clkbuf_2 _1025_ (.A(net294),
    .X(net367));
 sky130_fd_sc_hd__clkbuf_2 _1026_ (.A(net295),
    .X(net368));
 sky130_fd_sc_hd__clkbuf_2 _1027_ (.A(net296),
    .X(net369));
 sky130_fd_sc_hd__clkbuf_2 _1028_ (.A(net297),
    .X(net370));
 sky130_fd_sc_hd__clkbuf_2 _1029_ (.A(net298),
    .X(net371));
 sky130_fd_sc_hd__clkbuf_2 _1030_ (.A(net299),
    .X(net372));
 sky130_fd_sc_hd__clkbuf_2 _1031_ (.A(net301),
    .X(net374));
 sky130_fd_sc_hd__clkbuf_2 _1032_ (.A(net302),
    .X(net375));
 sky130_fd_sc_hd__clkbuf_2 _1033_ (.A(net303),
    .X(net376));
 sky130_fd_sc_hd__clkbuf_2 _1034_ (.A(net304),
    .X(net377));
 sky130_fd_sc_hd__clkbuf_2 _1035_ (.A(net305),
    .X(net378));
 sky130_fd_sc_hd__clkbuf_2 _1036_ (.A(net306),
    .X(net379));
 sky130_fd_sc_hd__clkbuf_2 _1037_ (.A(net307),
    .X(net380));
 sky130_fd_sc_hd__clkbuf_2 _1038_ (.A(net308),
    .X(net381));
 sky130_fd_sc_hd__clkbuf_2 _1039_ (.A(net309),
    .X(net382));
 sky130_fd_sc_hd__clkbuf_2 _1040_ (.A(net310),
    .X(net383));
 sky130_fd_sc_hd__clkbuf_2 _1041_ (.A(net312),
    .X(net385));
 sky130_fd_sc_hd__clkbuf_2 _1042_ (.A(net313),
    .X(net386));
 sky130_fd_sc_hd__clkbuf_2 _1043_ (.A(net314),
    .X(net387));
 sky130_fd_sc_hd__clkbuf_2 _1044_ (.A(net315),
    .X(net388));
 sky130_fd_sc_hd__clkbuf_2 _1045_ (.A(net316),
    .X(net389));
 sky130_fd_sc_hd__clkbuf_2 _1046_ (.A(net317),
    .X(net390));
 sky130_fd_sc_hd__clkbuf_2 _1047_ (.A(net318),
    .X(net391));
 sky130_fd_sc_hd__clkbuf_2 _1048_ (.A(net319),
    .X(net392));
 sky130_fd_sc_hd__clkbuf_2 _1049_ (.A(net1),
    .X(net393));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_wb_clk_i (.A(wb_clk_i),
    .X(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_0_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_10_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_11_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_12_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_13_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_14_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_15_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_1_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_2_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_3_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_4_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_5_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_6_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_7_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_8_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_9_0_wb_clk_i));
 sky130_fd_sc_hd__buf_4 fanout437 (.A(net438),
    .X(net437));
 sky130_fd_sc_hd__buf_4 fanout438 (.A(net440),
    .X(net438));
 sky130_fd_sc_hd__buf_4 fanout439 (.A(net440),
    .X(net439));
 sky130_fd_sc_hd__buf_2 fanout440 (.A(_0310_),
    .X(net440));
 sky130_fd_sc_hd__buf_4 fanout441 (.A(net442),
    .X(net441));
 sky130_fd_sc_hd__buf_4 fanout442 (.A(_0198_),
    .X(net442));
 sky130_fd_sc_hd__buf_4 fanout443 (.A(net444),
    .X(net443));
 sky130_fd_sc_hd__clkbuf_4 fanout444 (.A(_0197_),
    .X(net444));
 sky130_fd_sc_hd__buf_4 fanout445 (.A(_0260_),
    .X(net445));
 sky130_fd_sc_hd__buf_2 fanout446 (.A(_0260_),
    .X(net446));
 sky130_fd_sc_hd__clkbuf_4 fanout447 (.A(net448),
    .X(net447));
 sky130_fd_sc_hd__buf_4 fanout448 (.A(_0195_),
    .X(net448));
 sky130_fd_sc_hd__buf_4 fanout452 (.A(net453),
    .X(net452));
 sky130_fd_sc_hd__buf_4 fanout453 (.A(net454),
    .X(net453));
 sky130_fd_sc_hd__buf_4 fanout454 (.A(net565),
    .X(net454));
 sky130_fd_sc_hd__buf_4 fanout455 (.A(net456),
    .X(net455));
 sky130_fd_sc_hd__buf_4 fanout456 (.A(net565),
    .X(net456));
 sky130_fd_sc_hd__buf_8 fanout457 (.A(net458),
    .X(net457));
 sky130_fd_sc_hd__buf_8 fanout458 (.A(net459),
    .X(net458));
 sky130_fd_sc_hd__clkbuf_8 fanout459 (.A(net573),
    .X(net459));
 sky130_fd_sc_hd__buf_8 fanout460 (.A(net461),
    .X(net460));
 sky130_fd_sc_hd__buf_8 fanout461 (.A(net573),
    .X(net461));
 sky130_fd_sc_hd__buf_4 fanout462 (.A(net464),
    .X(net462));
 sky130_fd_sc_hd__buf_4 fanout463 (.A(net464),
    .X(net463));
 sky130_fd_sc_hd__buf_4 fanout464 (.A(net581),
    .X(net464));
 sky130_fd_sc_hd__buf_4 fanout465 (.A(net466),
    .X(net465));
 sky130_fd_sc_hd__buf_4 fanout466 (.A(net581),
    .X(net466));
 sky130_fd_sc_hd__buf_4 fanout467 (.A(_0237_),
    .X(net467));
 sky130_fd_sc_hd__buf_4 fanout468 (.A(_0237_),
    .X(net468));
 sky130_fd_sc_hd__buf_4 fanout469 (.A(net1081),
    .X(net469));
 sky130_fd_sc_hd__buf_4 fanout470 (.A(net1081),
    .X(net470));
 sky130_fd_sc_hd__buf_4 fanout471 (.A(net476),
    .X(net471));
 sky130_fd_sc_hd__clkbuf_4 fanout472 (.A(net476),
    .X(net472));
 sky130_fd_sc_hd__buf_4 fanout473 (.A(net476),
    .X(net473));
 sky130_fd_sc_hd__buf_4 fanout474 (.A(net475),
    .X(net474));
 sky130_fd_sc_hd__buf_4 fanout475 (.A(net476),
    .X(net475));
 sky130_fd_sc_hd__clkbuf_4 fanout476 (.A(_0113_),
    .X(net476));
 sky130_fd_sc_hd__clkbuf_8 fanout477 (.A(net218),
    .X(net477));
 sky130_fd_sc_hd__clkbuf_4 fanout478 (.A(net218),
    .X(net478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(net924),
    .X(net484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(net938),
    .X(net493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(net591),
    .X(net583));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold101 (.A(net559),
    .X(net584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(_0118_),
    .X(net585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(net601),
    .X(net586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(net603),
    .X(net587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(_0069_),
    .X(net588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(\design_select[0] ),
    .X(net589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(net579),
    .X(net590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(\design_select[1] ),
    .X(net591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(net583),
    .X(net592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(net939),
    .X(net494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(net597),
    .X(net593));
 sky130_fd_sc_hd__buf_1 hold111 (.A(net599),
    .X(net594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(net600),
    .X(net595));
 sky130_fd_sc_hd__buf_1 hold113 (.A(net602),
    .X(net596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(\design_select[2] ),
    .X(net597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(net593),
    .X(net598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(net571),
    .X(net599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(\design_select[3] ),
    .X(net600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(net595),
    .X(net601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(net586),
    .X(net602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(net941),
    .X(net495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(wb_feedback_delay),
    .X(net603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(net587),
    .X(net604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(_0000_),
    .X(net605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(net1153),
    .X(net606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(net1079),
    .X(net607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(net1137),
    .X(net608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(net1063),
    .X(net609));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold127 (.A(net1239),
    .X(net610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(_0357_),
    .X(net611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(_0358_),
    .X(net612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(net942),
    .X(net496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(_0086_),
    .X(net613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(net1142),
    .X(net614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(net1022),
    .X(net615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(net1140),
    .X(net616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(net1037),
    .X(net617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(net1155),
    .X(net618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(net1044),
    .X(net619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(net1159),
    .X(net620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(net1091),
    .X(net621));
 sky130_fd_sc_hd__buf_1 hold139 (.A(net1237),
    .X(net622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(net944),
    .X(net497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(_0347_),
    .X(net623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(_0349_),
    .X(net624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(_0083_),
    .X(net625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(net1143),
    .X(net626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(net1073),
    .X(net627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(net263),
    .X(net628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(_0213_),
    .X(net629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(_0015_),
    .X(net630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(net1141),
    .X(net631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(net1066),
    .X(net632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(net945),
    .X(net498));
 sky130_fd_sc_hd__buf_1 hold150 (.A(net1241),
    .X(net633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(_0335_),
    .X(net634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(_0337_),
    .X(net635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(_0079_),
    .X(net636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(net264),
    .X(net637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(_0214_),
    .X(net638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(_0016_),
    .X(net639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(net261),
    .X(net640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(_0211_),
    .X(net641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(_0013_),
    .X(net642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(net947),
    .X(net499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(net1161),
    .X(net643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(net1109),
    .X(net644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(net1144),
    .X(net645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(net1026),
    .X(net646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(net259),
    .X(net647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(_0209_),
    .X(net648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(_0011_),
    .X(net649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(net1145),
    .X(net650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(net1076),
    .X(net651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(net1146),
    .X(net652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(net948),
    .X(net500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(net1060),
    .X(net653));
 sky130_fd_sc_hd__buf_1 hold171 (.A(net1223),
    .X(net654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(_0393_),
    .X(net655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(_0394_),
    .X(net656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(_0098_),
    .X(net657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(\wb_counter[11] ),
    .X(net658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(_0340_),
    .X(net659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(_0343_),
    .X(net660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(_0081_),
    .X(net661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(net1164),
    .X(net662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(net950),
    .X(net501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(net1057),
    .X(net663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(net1147),
    .X(net664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(net1041),
    .X(net665));
 sky130_fd_sc_hd__buf_1 hold183 (.A(net1150),
    .X(net666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(net1103),
    .X(net667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(net1148),
    .X(net668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(net1085),
    .X(net669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(net288),
    .X(net670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(_0207_),
    .X(net671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(_0009_),
    .X(net672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(net951),
    .X(net502));
 sky130_fd_sc_hd__buf_1 hold190 (.A(net1215),
    .X(net673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold191 (.A(_0388_),
    .X(net674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(_0389_),
    .X(net675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(net1149),
    .X(net676));
 sky130_fd_sc_hd__buf_1 hold194 (.A(net1125),
    .X(net677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(_0328_),
    .X(net678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(_0331_),
    .X(net679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold197 (.A(_0077_),
    .X(net680));
 sky130_fd_sc_hd__buf_1 hold198 (.A(net1151),
    .X(net681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(net1088),
    .X(net682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(net926),
    .X(net485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(net953),
    .X(net503));
 sky130_fd_sc_hd__buf_1 hold200 (.A(net1152),
    .X(net683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(net1050),
    .X(net684));
 sky130_fd_sc_hd__buf_1 hold202 (.A(net1222),
    .X(net685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(_0363_),
    .X(net686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(_0365_),
    .X(net687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(net1187),
    .X(net688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(net272),
    .X(net689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(_0221_),
    .X(net690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(_0023_),
    .X(net691));
 sky130_fd_sc_hd__buf_1 hold209 (.A(net1136),
    .X(net692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(net954),
    .X(net504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold210 (.A(net1054),
    .X(net693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(net271),
    .X(net694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(_0220_),
    .X(net695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold213 (.A(_0022_),
    .X(net696));
 sky130_fd_sc_hd__buf_1 hold214 (.A(net1168),
    .X(net697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(net1018),
    .X(net698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(net283),
    .X(net699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold217 (.A(_0202_),
    .X(net700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold218 (.A(_0004_),
    .X(net701));
 sky130_fd_sc_hd__buf_1 hold219 (.A(net1156),
    .X(net702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(net956),
    .X(net505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(net1094),
    .X(net703));
 sky130_fd_sc_hd__buf_1 hold221 (.A(net1157),
    .X(net704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold222 (.A(net1069),
    .X(net705));
 sky130_fd_sc_hd__buf_1 hold223 (.A(net1228),
    .X(net706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(_0359_),
    .X(net707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold225 (.A(_0362_),
    .X(net708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold226 (.A(_0087_),
    .X(net709));
 sky130_fd_sc_hd__buf_1 hold227 (.A(net1230),
    .X(net710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold228 (.A(_0371_),
    .X(net711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold229 (.A(_0372_),
    .X(net712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(net981),
    .X(net506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold230 (.A(_0090_),
    .X(net713));
 sky130_fd_sc_hd__buf_1 hold231 (.A(net1160),
    .X(net714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold232 (.A(_0369_),
    .X(net715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold233 (.A(_0089_),
    .X(net716));
 sky130_fd_sc_hd__buf_1 hold234 (.A(net1158),
    .X(net717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold235 (.A(net1030),
    .X(net718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold236 (.A(net273),
    .X(net719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold237 (.A(_0222_),
    .X(net720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(_0024_),
    .X(net721));
 sky130_fd_sc_hd__buf_1 hold239 (.A(net1227),
    .X(net722));
 sky130_fd_sc_hd__buf_1 hold24 (.A(net253),
    .X(net507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold240 (.A(_0390_),
    .X(net723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(net1154),
    .X(net724));
 sky130_fd_sc_hd__buf_1 hold242 (.A(net1134),
    .X(net725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold243 (.A(net1135),
    .X(net726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold244 (.A(net274),
    .X(net727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold245 (.A(_0223_),
    .X(net728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold246 (.A(_0025_),
    .X(net729));
 sky130_fd_sc_hd__clkbuf_2 hold247 (.A(net898),
    .X(net730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold248 (.A(_0268_),
    .X(net731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold249 (.A(_0048_),
    .X(net732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(net983),
    .X(net508));
 sky130_fd_sc_hd__buf_1 hold250 (.A(net1221),
    .X(net733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold251 (.A(_0104_),
    .X(net734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold252 (.A(_0099_),
    .X(net735));
 sky130_fd_sc_hd__clkbuf_2 hold253 (.A(net891),
    .X(net736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold254 (.A(_0308_),
    .X(net737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold255 (.A(_0068_),
    .X(net738));
 sky130_fd_sc_hd__clkbuf_2 hold256 (.A(net894),
    .X(net739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold257 (.A(_0300_),
    .X(net740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold258 (.A(_0064_),
    .X(net741));
 sky130_fd_sc_hd__clkbuf_2 hold259 (.A(net912),
    .X(net742));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold26 (.A(net227),
    .X(net509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold260 (.A(_0292_),
    .X(net743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold261 (.A(_0060_),
    .X(net744));
 sky130_fd_sc_hd__clkbuf_2 hold262 (.A(net895),
    .X(net745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold263 (.A(_0304_),
    .X(net746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold264 (.A(_0066_),
    .X(net747));
 sky130_fd_sc_hd__clkbuf_2 hold265 (.A(net915),
    .X(net748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold266 (.A(_0282_),
    .X(net749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold267 (.A(_0055_),
    .X(net750));
 sky130_fd_sc_hd__clkbuf_2 hold268 (.A(net896),
    .X(net751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold269 (.A(_0296_),
    .X(net752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(net985),
    .X(net510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold270 (.A(_0062_),
    .X(net753));
 sky130_fd_sc_hd__clkbuf_2 hold271 (.A(net910),
    .X(net754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold272 (.A(_0270_),
    .X(net755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold273 (.A(_0049_),
    .X(net756));
 sky130_fd_sc_hd__clkbuf_2 hold274 (.A(net914),
    .X(net757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold275 (.A(_0272_),
    .X(net758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold276 (.A(_0050_),
    .X(net759));
 sky130_fd_sc_hd__clkbuf_2 hold277 (.A(net918),
    .X(net760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold278 (.A(_0284_),
    .X(net761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold279 (.A(_0056_),
    .X(net762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(net226),
    .X(net511));
 sky130_fd_sc_hd__clkbuf_2 hold280 (.A(net917),
    .X(net763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold281 (.A(_0288_),
    .X(net764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold282 (.A(_0058_),
    .X(net765));
 sky130_fd_sc_hd__clkbuf_2 hold283 (.A(net913),
    .X(net766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold284 (.A(_0276_),
    .X(net767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold285 (.A(_0052_),
    .X(net768));
 sky130_fd_sc_hd__clkbuf_2 hold286 (.A(net897),
    .X(net769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold287 (.A(_0306_),
    .X(net770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold288 (.A(_0067_),
    .X(net771));
 sky130_fd_sc_hd__clkbuf_2 hold289 (.A(net902),
    .X(net772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(net989),
    .X(net512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold290 (.A(_0294_),
    .X(net773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold291 (.A(_0061_),
    .X(net774));
 sky130_fd_sc_hd__clkbuf_2 hold292 (.A(net919),
    .X(net775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold293 (.A(_0286_),
    .X(net776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold294 (.A(_0057_),
    .X(net777));
 sky130_fd_sc_hd__clkbuf_2 hold295 (.A(net921),
    .X(net778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold296 (.A(_0290_),
    .X(net779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold297 (.A(_0059_),
    .X(net780));
 sky130_fd_sc_hd__clkbuf_2 hold298 (.A(net920),
    .X(net781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold299 (.A(_0280_),
    .X(net782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(net933),
    .X(net486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(net254),
    .X(net513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold300 (.A(_0054_),
    .X(net783));
 sky130_fd_sc_hd__clkbuf_2 hold301 (.A(net900),
    .X(net784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold302 (.A(_0298_),
    .X(net785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold303 (.A(_0063_),
    .X(net786));
 sky130_fd_sc_hd__clkbuf_2 hold304 (.A(net901),
    .X(net787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold305 (.A(_0264_),
    .X(net788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold306 (.A(_0046_),
    .X(net789));
 sky130_fd_sc_hd__clkbuf_2 hold307 (.A(net911),
    .X(net790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold308 (.A(_0262_),
    .X(net791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold309 (.A(_0045_),
    .X(net792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(net991),
    .X(net514));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold310 (.A(net876),
    .X(net793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold311 (.A(_0006_),
    .X(net794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold312 (.A(net268),
    .X(net795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold313 (.A(_0218_),
    .X(net796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold314 (.A(_0020_),
    .X(net797));
 sky130_fd_sc_hd__clkbuf_2 hold315 (.A(net899),
    .X(net798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold316 (.A(_0302_),
    .X(net799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold317 (.A(_0065_),
    .X(net800));
 sky130_fd_sc_hd__buf_1 hold318 (.A(net1123),
    .X(net801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold319 (.A(_0322_),
    .X(net802));
 sky130_fd_sc_hd__buf_1 hold32 (.A(net225),
    .X(net515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold320 (.A(_0324_),
    .X(net803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold321 (.A(_0075_),
    .X(net804));
 sky130_fd_sc_hd__clkbuf_2 hold322 (.A(net916),
    .X(net805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold323 (.A(_0278_),
    .X(net806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold324 (.A(_0053_),
    .X(net807));
 sky130_fd_sc_hd__clkbuf_2 hold325 (.A(net922),
    .X(net808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold326 (.A(_0274_),
    .X(net809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold327 (.A(_0051_),
    .X(net810));
 sky130_fd_sc_hd__clkbuf_2 hold328 (.A(net905),
    .X(net811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold329 (.A(_0266_),
    .X(net812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(net957),
    .X(net516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold330 (.A(_0047_),
    .X(net813));
 sky130_fd_sc_hd__clkbuf_2 hold331 (.A(net1127),
    .X(net814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold332 (.A(_0311_),
    .X(net815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold333 (.A(_0070_),
    .X(net816));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold334 (.A(net880),
    .X(net817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold335 (.A(net1217),
    .X(net818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold336 (.A(net284),
    .X(net819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold337 (.A(_0203_),
    .X(net820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold338 (.A(_0005_),
    .X(net821));
 sky130_fd_sc_hd__clkbuf_2 hold339 (.A(net892),
    .X(net822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(net959),
    .X(net517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold340 (.A(net1207),
    .X(net823));
 sky130_fd_sc_hd__clkbuf_2 hold341 (.A(net903),
    .X(net824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold342 (.A(net1198),
    .X(net825));
 sky130_fd_sc_hd__clkbuf_2 hold343 (.A(net906),
    .X(net826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold344 (.A(net1196),
    .X(net827));
 sky130_fd_sc_hd__clkbuf_2 hold345 (.A(net893),
    .X(net828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold346 (.A(net1200),
    .X(net829));
 sky130_fd_sc_hd__clkbuf_2 hold347 (.A(net908),
    .X(net830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold348 (.A(net1202),
    .X(net831));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold349 (.A(net1231),
    .X(net832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(net993),
    .X(net518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold350 (.A(_0106_),
    .X(net833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold351 (.A(_0100_),
    .X(net834));
 sky130_fd_sc_hd__clkbuf_2 hold352 (.A(net904),
    .X(net835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold353 (.A(net1189),
    .X(net836));
 sky130_fd_sc_hd__clkbuf_2 hold354 (.A(net907),
    .X(net837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold355 (.A(net1209),
    .X(net838));
 sky130_fd_sc_hd__clkbuf_2 hold356 (.A(net909),
    .X(net839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold357 (.A(net1191),
    .X(net840));
 sky130_fd_sc_hd__buf_1 hold358 (.A(net1235),
    .X(net841));
 sky130_fd_sc_hd__buf_1 hold359 (.A(_0383_),
    .X(net842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(net255),
    .X(net519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold360 (.A(_0385_),
    .X(net843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold361 (.A(net1162),
    .X(net844));
 sky130_fd_sc_hd__buf_1 hold362 (.A(net1163),
    .X(net845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold363 (.A(net1033),
    .X(net846));
 sky130_fd_sc_hd__clkbuf_2 hold364 (.A(net1167),
    .X(net847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold365 (.A(net1177),
    .X(net848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold366 (.A(\wb_counter[31] ),
    .X(net849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold367 (.A(_0109_),
    .X(net850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold368 (.A(net1165),
    .X(net851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold369 (.A(net884),
    .X(net852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(net997),
    .X(net520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold370 (.A(_0003_),
    .X(net853));
 sky130_fd_sc_hd__buf_1 hold371 (.A(net1169),
    .X(net854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold372 (.A(net1112),
    .X(net855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold373 (.A(\wbs_adr_delaybuff[2] ),
    .X(net856));
 sky130_fd_sc_hd__buf_2 hold374 (.A(net1175),
    .X(net857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold375 (.A(_0234_),
    .X(net858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold376 (.A(_0034_),
    .X(net859));
 sky130_fd_sc_hd__buf_1 hold377 (.A(net1129),
    .X(net860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold378 (.A(_0312_),
    .X(net861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold379 (.A(_0314_),
    .X(net862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(net231),
    .X(net521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold380 (.A(_0071_),
    .X(net863));
 sky130_fd_sc_hd__buf_1 hold381 (.A(net1170),
    .X(net864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold382 (.A(net1106),
    .X(net865));
 sky130_fd_sc_hd__buf_1 hold383 (.A(net1121),
    .X(net866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold384 (.A(_0326_),
    .X(net867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold385 (.A(_0327_),
    .X(net868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold386 (.A(_0076_),
    .X(net869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold387 (.A(\wbs_adr_delaybuff[3] ),
    .X(net870));
 sky130_fd_sc_hd__buf_2 hold388 (.A(_0194_),
    .X(net871));
 sky130_fd_sc_hd__buf_2 hold389 (.A(net1179),
    .X(net872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(net999),
    .X(net522));
 sky130_fd_sc_hd__clkbuf_2 hold390 (.A(_0232_),
    .X(net873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold391 (.A(_0112_),
    .X(net874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold392 (.A(_0103_),
    .X(net875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold393 (.A(net1219),
    .X(net876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold394 (.A(net793),
    .X(net877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold395 (.A(_0236_),
    .X(net878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold396 (.A(_0036_),
    .X(net879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold397 (.A(net1216),
    .X(net880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold398 (.A(net817),
    .X(net881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold399 (.A(_0235_),
    .X(net882));
 sky130_fd_sc_hd__buf_1 hold4 (.A(net935),
    .X(net487));
 sky130_fd_sc_hd__buf_1 hold40 (.A(net229),
    .X(net523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold400 (.A(_0035_),
    .X(net883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold401 (.A(\wbs_dat_delaybuff[2] ),
    .X(net884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold402 (.A(net852),
    .X(net885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold403 (.A(_0233_),
    .X(net886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold404 (.A(_0033_),
    .X(net887));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold405 (.A(net1131),
    .X(net888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold406 (.A(_0315_),
    .X(net889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold407 (.A(_0072_),
    .X(net890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold408 (.A(net1243),
    .X(net891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold409 (.A(net1206),
    .X(net892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(net1001),
    .X(net524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold410 (.A(net1199),
    .X(net893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold411 (.A(net1233),
    .X(net894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold412 (.A(net1252),
    .X(net895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold413 (.A(net1245),
    .X(net896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold414 (.A(net1236),
    .X(net897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold415 (.A(net1257),
    .X(net898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold416 (.A(net1253),
    .X(net899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold417 (.A(net1244),
    .X(net900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold418 (.A(net1249),
    .X(net901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold419 (.A(net1246),
    .X(net902));
 sky130_fd_sc_hd__buf_1 hold42 (.A(net230),
    .X(net525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold420 (.A(net1197),
    .X(net903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold421 (.A(net1188),
    .X(net904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold422 (.A(net1247),
    .X(net905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold423 (.A(net1195),
    .X(net906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold424 (.A(net1208),
    .X(net907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold425 (.A(net1201),
    .X(net908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold426 (.A(net1190),
    .X(net909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold427 (.A(net1263),
    .X(net910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold428 (.A(net1256),
    .X(net911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold429 (.A(net1258),
    .X(net912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(net960),
    .X(net526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold430 (.A(net1250),
    .X(net913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold431 (.A(net1261),
    .X(net914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold432 (.A(net1255),
    .X(net915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold433 (.A(net1254),
    .X(net916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold434 (.A(net1251),
    .X(net917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold435 (.A(net1259),
    .X(net918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold436 (.A(net1260),
    .X(net919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold437 (.A(net1262),
    .X(net920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold438 (.A(net1264),
    .X(net921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold439 (.A(net1248),
    .X(net922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(net962),
    .X(net527));
 sky130_fd_sc_hd__buf_2 hold440 (.A(net1226),
    .X(net923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold441 (.A(wbs_adr_i[2]),
    .X(net924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold442 (.A(net484),
    .X(net925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold443 (.A(net220),
    .X(net926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold444 (.A(wbs_adr_i[4]),
    .X(net927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold445 (.A(net488),
    .X(net928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold446 (.A(net222),
    .X(net929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold447 (.A(wbs_adr_i[3]),
    .X(net930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold448 (.A(net490),
    .X(net931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold449 (.A(net221),
    .X(net932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(net1003),
    .X(net528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold450 (.A(net1229),
    .X(net933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold451 (.A(net486),
    .X(net934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold452 (.A(net219),
    .X(net935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold453 (.A(wbs_dat_i[4]),
    .X(net936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold454 (.A(net492),
    .X(net937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold455 (.A(net250),
    .X(net938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold456 (.A(wbs_dat_i[1]),
    .X(net939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold457 (.A(net494),
    .X(net940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold458 (.A(net235),
    .X(net941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold459 (.A(wbs_dat_i[2]),
    .X(net942));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold46 (.A(net228),
    .X(net529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold460 (.A(net496),
    .X(net943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold461 (.A(net246),
    .X(net944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold462 (.A(wbs_dat_i[0]),
    .X(net945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold463 (.A(net498),
    .X(net946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold464 (.A(net224),
    .X(net947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold465 (.A(wbs_dat_i[6]),
    .X(net948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold466 (.A(net500),
    .X(net949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold467 (.A(net252),
    .X(net950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold468 (.A(wbs_dat_i[5]),
    .X(net951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold469 (.A(net502),
    .X(net952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(net995),
    .X(net530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold470 (.A(net251),
    .X(net953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold471 (.A(wbs_dat_i[3]),
    .X(net954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold472 (.A(net504),
    .X(net955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold473 (.A(net249),
    .X(net956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold474 (.A(wbs_dat_i[19]),
    .X(net957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold475 (.A(net516),
    .X(net958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold476 (.A(net234),
    .X(net959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold477 (.A(wbs_dat_i[23]),
    .X(net960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold478 (.A(net526),
    .X(net961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold479 (.A(net239),
    .X(net962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(net248),
    .X(net531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold480 (.A(wbs_dat_i[20]),
    .X(net963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold481 (.A(net532),
    .X(net964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold482 (.A(net236),
    .X(net965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold483 (.A(wbs_dat_i[21]),
    .X(net966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold484 (.A(net534),
    .X(net967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold485 (.A(net237),
    .X(net968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold486 (.A(wbs_dat_i[24]),
    .X(net969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold487 (.A(net536),
    .X(net970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold488 (.A(net240),
    .X(net971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold489 (.A(wbs_dat_i[18]),
    .X(net972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(net963),
    .X(net532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold490 (.A(net540),
    .X(net973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold491 (.A(net233),
    .X(net974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold492 (.A(wbs_dat_i[17]),
    .X(net975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold493 (.A(net544),
    .X(net976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold494 (.A(net232),
    .X(net977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold495 (.A(wbs_dat_i[22]),
    .X(net978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold496 (.A(net546),
    .X(net979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold497 (.A(net238),
    .X(net980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold498 (.A(net1181),
    .X(net981));
 sky130_fd_sc_hd__dlygate4sd3_1 hold499 (.A(net506),
    .X(net982));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(net927),
    .X(net488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(net965),
    .X(net533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold500 (.A(net1218),
    .X(net983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold501 (.A(net508),
    .X(net984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold502 (.A(wbs_dat_i[11]),
    .X(net985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold503 (.A(net510),
    .X(net986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold504 (.A(wbs_dat_i[25]),
    .X(net987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold505 (.A(net548),
    .X(net988));
 sky130_fd_sc_hd__dlygate4sd3_1 hold506 (.A(wbs_dat_i[8]),
    .X(net989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold507 (.A(net512),
    .X(net990));
 sky130_fd_sc_hd__dlygate4sd3_1 hold508 (.A(net1183),
    .X(net991));
 sky130_fd_sc_hd__dlygate4sd3_1 hold509 (.A(net514),
    .X(net992));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(net966),
    .X(net534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold510 (.A(wbs_dat_i[9]),
    .X(net993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold511 (.A(net518),
    .X(net994));
 sky130_fd_sc_hd__dlygate4sd3_1 hold512 (.A(wbs_dat_i[31]),
    .X(net995));
 sky130_fd_sc_hd__dlygate4sd3_1 hold513 (.A(net530),
    .X(net996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold514 (.A(wbs_dat_i[16]),
    .X(net997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold515 (.A(net520),
    .X(net998));
 sky130_fd_sc_hd__dlygate4sd3_1 hold516 (.A(net1184),
    .X(net999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold517 (.A(net522),
    .X(net1000));
 sky130_fd_sc_hd__dlygate4sd3_1 hold518 (.A(net1182),
    .X(net1001));
 sky130_fd_sc_hd__dlygate4sd3_1 hold519 (.A(net524),
    .X(net1002));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(net968),
    .X(net535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold520 (.A(net1224),
    .X(net1003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold521 (.A(net528),
    .X(net1004));
 sky130_fd_sc_hd__dlygate4sd3_1 hold522 (.A(wbs_dat_i[30]),
    .X(net1005));
 sky130_fd_sc_hd__dlygate4sd3_1 hold523 (.A(net538),
    .X(net1006));
 sky130_fd_sc_hd__dlygate4sd3_1 hold524 (.A(wbs_dat_i[29]),
    .X(net1007));
 sky130_fd_sc_hd__dlygate4sd3_1 hold525 (.A(net542),
    .X(net1008));
 sky130_fd_sc_hd__dlygate4sd3_1 hold526 (.A(wbs_dat_i[26]),
    .X(net1009));
 sky130_fd_sc_hd__dlygate4sd3_1 hold527 (.A(net552),
    .X(net1010));
 sky130_fd_sc_hd__dlygate4sd3_1 hold528 (.A(wbs_dat_i[28]),
    .X(net1011));
 sky130_fd_sc_hd__dlygate4sd3_1 hold529 (.A(net550),
    .X(net1012));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(net969),
    .X(net536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold530 (.A(wbs_dat_i[27]),
    .X(net1013));
 sky130_fd_sc_hd__dlygate4sd3_1 hold531 (.A(net554),
    .X(net1014));
 sky130_fd_sc_hd__dlygate4sd3_1 hold532 (.A(\wb_counter[3] ),
    .X(net1015));
 sky130_fd_sc_hd__dlygate4sd3_1 hold533 (.A(_0318_),
    .X(net1016));
 sky130_fd_sc_hd__dlygate4sd3_1 hold534 (.A(_0319_),
    .X(net1017));
 sky130_fd_sc_hd__dlygate4sd3_1 hold535 (.A(_0073_),
    .X(net1018));
 sky130_fd_sc_hd__dlygate4sd3_1 hold536 (.A(\wb_counter[15] ),
    .X(net1019));
 sky130_fd_sc_hd__dlygate4sd3_1 hold537 (.A(_0353_),
    .X(net1020));
 sky130_fd_sc_hd__dlygate4sd3_1 hold538 (.A(_0356_),
    .X(net1021));
 sky130_fd_sc_hd__dlygate4sd3_1 hold539 (.A(_0085_),
    .X(net1022));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(net971),
    .X(net537));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold540 (.A(net1265),
    .X(net1023));
 sky130_fd_sc_hd__dlygate4sd3_1 hold541 (.A(_0338_),
    .X(net1024));
 sky130_fd_sc_hd__dlygate4sd3_1 hold542 (.A(_0339_),
    .X(net1025));
 sky130_fd_sc_hd__dlygate4sd3_1 hold543 (.A(_0080_),
    .X(net1026));
 sky130_fd_sc_hd__dlygate4sd3_1 hold544 (.A(\wb_counter[23] ),
    .X(net1027));
 sky130_fd_sc_hd__dlygate4sd3_1 hold545 (.A(_0379_),
    .X(net1028));
 sky130_fd_sc_hd__dlygate4sd3_1 hold546 (.A(_0381_),
    .X(net1029));
 sky130_fd_sc_hd__dlygate4sd3_1 hold547 (.A(_0093_),
    .X(net1030));
 sky130_fd_sc_hd__dlygate4sd3_1 hold548 (.A(net258),
    .X(net1031));
 sky130_fd_sc_hd__dlygate4sd3_1 hold549 (.A(_0199_),
    .X(net1032));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(net1005),
    .X(net538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold550 (.A(_0001_),
    .X(net1033));
 sky130_fd_sc_hd__buf_1 hold551 (.A(net1240),
    .X(net1034));
 sky130_fd_sc_hd__dlygate4sd3_1 hold552 (.A(_0350_),
    .X(net1035));
 sky130_fd_sc_hd__dlygate4sd3_1 hold553 (.A(_0352_),
    .X(net1036));
 sky130_fd_sc_hd__dlygate4sd3_1 hold554 (.A(_0084_),
    .X(net1037));
 sky130_fd_sc_hd__buf_1 hold555 (.A(net1234),
    .X(net1038));
 sky130_fd_sc_hd__dlygate4sd3_1 hold556 (.A(_0332_),
    .X(net1039));
 sky130_fd_sc_hd__dlygate4sd3_1 hold557 (.A(_0334_),
    .X(net1040));
 sky130_fd_sc_hd__dlygate4sd3_1 hold558 (.A(_0078_),
    .X(net1041));
 sky130_fd_sc_hd__dlygate4sd3_1 hold559 (.A(net279),
    .X(net1042));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(net247),
    .X(net539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold560 (.A(_0228_),
    .X(net1043));
 sky130_fd_sc_hd__dlygate4sd3_1 hold561 (.A(_0030_),
    .X(net1044));
 sky130_fd_sc_hd__buf_1 hold562 (.A(net1220),
    .X(net1045));
 sky130_fd_sc_hd__dlygate4sd3_1 hold563 (.A(_0320_),
    .X(net1046));
 sky130_fd_sc_hd__buf_1 hold564 (.A(net1225),
    .X(net1047));
 sky130_fd_sc_hd__dlygate4sd3_1 hold565 (.A(_0376_),
    .X(net1048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold566 (.A(_0378_),
    .X(net1049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold567 (.A(_0092_),
    .X(net1050));
 sky130_fd_sc_hd__buf_1 hold568 (.A(net1232),
    .X(net1051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold569 (.A(_0373_),
    .X(net1052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(net972),
    .X(net540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold570 (.A(_0375_),
    .X(net1053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold571 (.A(_0091_),
    .X(net1054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold572 (.A(net282),
    .X(net1055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold573 (.A(_0230_),
    .X(net1056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold574 (.A(_0032_),
    .X(net1057));
 sky130_fd_sc_hd__dlygate4sd3_1 hold575 (.A(net278),
    .X(net1058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold576 (.A(_0227_),
    .X(net1059));
 sky130_fd_sc_hd__dlygate4sd3_1 hold577 (.A(_0029_),
    .X(net1060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold578 (.A(net265),
    .X(net1061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold579 (.A(_0215_),
    .X(net1062));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(net974),
    .X(net541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold580 (.A(_0017_),
    .X(net1063));
 sky130_fd_sc_hd__dlygate4sd3_1 hold581 (.A(net289),
    .X(net1064));
 sky130_fd_sc_hd__dlygate4sd3_1 hold582 (.A(_0208_),
    .X(net1065));
 sky130_fd_sc_hd__dlygate4sd3_1 hold583 (.A(_0010_),
    .X(net1066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold584 (.A(net270),
    .X(net1067));
 sky130_fd_sc_hd__dlygate4sd3_1 hold585 (.A(_0219_),
    .X(net1068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold586 (.A(_0021_),
    .X(net1069));
 sky130_fd_sc_hd__buf_1 hold587 (.A(net1242),
    .X(net1070));
 sky130_fd_sc_hd__dlygate4sd3_1 hold588 (.A(_0344_),
    .X(net1071));
 sky130_fd_sc_hd__dlygate4sd3_1 hold589 (.A(_0346_),
    .X(net1072));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(net1007),
    .X(net542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold590 (.A(_0082_),
    .X(net1073));
 sky130_fd_sc_hd__dlygate4sd3_1 hold591 (.A(net260),
    .X(net1074));
 sky130_fd_sc_hd__dlygate4sd3_1 hold592 (.A(_0210_),
    .X(net1075));
 sky130_fd_sc_hd__dlygate4sd3_1 hold593 (.A(_0012_),
    .X(net1076));
 sky130_fd_sc_hd__dlygate4sd3_1 hold594 (.A(net277),
    .X(net1077));
 sky130_fd_sc_hd__dlygate4sd3_1 hold595 (.A(_0226_),
    .X(net1078));
 sky130_fd_sc_hd__dlygate4sd3_1 hold596 (.A(_0028_),
    .X(net1079));
 sky130_fd_sc_hd__dlygate4sd3_1 hold597 (.A(\wbs_adr_delaybuff[1] ),
    .X(net1080));
 sky130_fd_sc_hd__clkbuf_2 hold598 (.A(_0192_),
    .X(net1081));
 sky130_fd_sc_hd__dlygate4sd3_1 hold599 (.A(_0248_),
    .X(net1082));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(net929),
    .X(net489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(net245),
    .X(net543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold600 (.A(net276),
    .X(net1083));
 sky130_fd_sc_hd__dlygate4sd3_1 hold601 (.A(_0225_),
    .X(net1084));
 sky130_fd_sc_hd__dlygate4sd3_1 hold602 (.A(_0027_),
    .X(net1085));
 sky130_fd_sc_hd__dlygate4sd3_1 hold603 (.A(net267),
    .X(net1086));
 sky130_fd_sc_hd__dlygate4sd3_1 hold604 (.A(_0217_),
    .X(net1087));
 sky130_fd_sc_hd__dlygate4sd3_1 hold605 (.A(_0019_),
    .X(net1088));
 sky130_fd_sc_hd__dlygate4sd3_1 hold606 (.A(net281),
    .X(net1089));
 sky130_fd_sc_hd__dlygate4sd3_1 hold607 (.A(_0229_),
    .X(net1090));
 sky130_fd_sc_hd__dlygate4sd3_1 hold608 (.A(_0031_),
    .X(net1091));
 sky130_fd_sc_hd__dlygate4sd3_1 hold609 (.A(net266),
    .X(net1092));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(net975),
    .X(net544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold610 (.A(_0216_),
    .X(net1093));
 sky130_fd_sc_hd__dlygate4sd3_1 hold611 (.A(_0018_),
    .X(net1094));
 sky130_fd_sc_hd__dlygate4sd3_1 hold612 (.A(net285),
    .X(net1095));
 sky130_fd_sc_hd__dlygate4sd3_1 hold613 (.A(_0204_),
    .X(net1096));
 sky130_fd_sc_hd__buf_1 hold614 (.A(net262),
    .X(net1097));
 sky130_fd_sc_hd__dlygate4sd3_1 hold615 (.A(_0212_),
    .X(net1098));
 sky130_fd_sc_hd__dlygate4sd3_1 hold616 (.A(_0014_),
    .X(net1099));
 sky130_fd_sc_hd__dlygate4sd3_1 hold617 (.A(net578),
    .X(net1100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold618 (.A(net287),
    .X(net1101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold619 (.A(_0206_),
    .X(net1102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(net977),
    .X(net545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold620 (.A(_0008_),
    .X(net1103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold621 (.A(net286),
    .X(net1104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold622 (.A(_0205_),
    .X(net1105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold623 (.A(_0007_),
    .X(net1106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold624 (.A(net275),
    .X(net1107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold625 (.A(_0224_),
    .X(net1108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold626 (.A(_0026_),
    .X(net1109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold627 (.A(net269),
    .X(net1110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold628 (.A(_0200_),
    .X(net1111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold629 (.A(_0002_),
    .X(net1112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(net978),
    .X(net546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold630 (.A(net280),
    .X(net1113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold631 (.A(_0201_),
    .X(net1114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold632 (.A(wb_rst_override),
    .X(net1115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold633 (.A(net556),
    .X(net1116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold634 (.A(net394),
    .X(net1117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold635 (.A(net557),
    .X(net1118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold636 (.A(\wbs_adr_delaybuff[0] ),
    .X(net1119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold637 (.A(_0251_),
    .X(net1120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold638 (.A(\wb_counter[6] ),
    .X(net1121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold639 (.A(_0256_),
    .X(net1122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(net980),
    .X(net547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold640 (.A(\wb_counter[5] ),
    .X(net1123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold641 (.A(_0254_),
    .X(net1124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold642 (.A(\wb_counter[7] ),
    .X(net1125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold643 (.A(_0258_),
    .X(net1126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold644 (.A(\wb_counter[0] ),
    .X(net1127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold645 (.A(_0239_),
    .X(net1128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold646 (.A(\wb_counter[1] ),
    .X(net1129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold647 (.A(_0242_),
    .X(net1130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold648 (.A(\wb_counter[2] ),
    .X(net1131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold649 (.A(net888),
    .X(net1132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(net987),
    .X(net548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold650 (.A(_0245_),
    .X(net1133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold651 (.A(net1193),
    .X(net1134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold652 (.A(_0094_),
    .X(net1135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold653 (.A(net1185),
    .X(net1136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold654 (.A(\wbs_dat_delaybuff[16] ),
    .X(net1137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold655 (.A(net608),
    .X(net1138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold656 (.A(\wbs_dat_delaybuff[13] ),
    .X(net1139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold657 (.A(\wbs_dat_delaybuff[14] ),
    .X(net1140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold658 (.A(\wbs_dat_delaybuff[9] ),
    .X(net1141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold659 (.A(\wbs_dat_delaybuff[15] ),
    .X(net1142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(net241),
    .X(net549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold660 (.A(\wbs_dat_delaybuff[12] ),
    .X(net1143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold661 (.A(\wbs_dat_delaybuff[10] ),
    .X(net1144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold662 (.A(\wbs_dat_delaybuff[11] ),
    .X(net1145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold663 (.A(\wbs_dat_delaybuff[28] ),
    .X(net1146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold664 (.A(\wbs_dat_delaybuff[8] ),
    .X(net1147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold665 (.A(\wbs_dat_delaybuff[26] ),
    .X(net1148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold666 (.A(_0096_),
    .X(net1149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold667 (.A(net1192),
    .X(net1150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold668 (.A(net1186),
    .X(net1151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold669 (.A(net1213),
    .X(net1152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(net1011),
    .X(net550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold670 (.A(\wbs_dat_delaybuff[27] ),
    .X(net1153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold671 (.A(_0097_),
    .X(net1154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold672 (.A(\wbs_dat_delaybuff[29] ),
    .X(net1155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold673 (.A(net1204),
    .X(net1156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold674 (.A(net1194),
    .X(net1157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold675 (.A(net1205),
    .X(net1158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold676 (.A(\wbs_dat_delaybuff[30] ),
    .X(net1159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold677 (.A(net1203),
    .X(net1160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold678 (.A(\wbs_dat_delaybuff[25] ),
    .X(net1161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold679 (.A(_0095_),
    .X(net1162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(net244),
    .X(net551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold680 (.A(net1212),
    .X(net1163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold681 (.A(\wbs_dat_delaybuff[31] ),
    .X(net1164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold682 (.A(_0101_),
    .X(net1165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold683 (.A(\wb_counter[19] ),
    .X(net1166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold684 (.A(wb_override_act),
    .X(net1167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold685 (.A(net1214),
    .X(net1168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold686 (.A(net1210),
    .X(net1169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold687 (.A(net1211),
    .X(net1170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold688 (.A(wbs_cyc_i),
    .X(net1171));
 sky130_fd_sc_hd__buf_1 hold689 (.A(_0191_),
    .X(net1172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(net1009),
    .X(net552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold690 (.A(net356),
    .X(net1173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold691 (.A(\wbs_adr_delaybuff[0] ),
    .X(net1174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold692 (.A(_0231_),
    .X(net1175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold693 (.A(_0111_),
    .X(net1176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold694 (.A(_0102_),
    .X(net1177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold695 (.A(wbs_we_i),
    .X(net1178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold696 (.A(_0196_),
    .X(net1179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold697 (.A(net872),
    .X(net1180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold698 (.A(wbs_dat_i[7]),
    .X(net1181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold699 (.A(wbs_dat_i[15]),
    .X(net1182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(net930),
    .X(net490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(net242),
    .X(net553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold700 (.A(wbs_dat_i[10]),
    .X(net1183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold701 (.A(wbs_dat_i[14]),
    .X(net1184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold702 (.A(\wbs_dat_delaybuff[21] ),
    .X(net1185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold703 (.A(\wbs_dat_delaybuff[18] ),
    .X(net1186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold704 (.A(_0088_),
    .X(net1187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold705 (.A(net431),
    .X(net1188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold706 (.A(_0041_),
    .X(net1189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold707 (.A(net433),
    .X(net1190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold708 (.A(_0043_),
    .X(net1191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold709 (.A(\wbs_dat_delaybuff[7] ),
    .X(net1192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(net1013),
    .X(net554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold710 (.A(\wbs_dat_delaybuff[24] ),
    .X(net1193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold711 (.A(\wbs_dat_delaybuff[20] ),
    .X(net1194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold712 (.A(net427),
    .X(net1195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold713 (.A(_0039_),
    .X(net1196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold714 (.A(net430),
    .X(net1197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold715 (.A(_0040_),
    .X(net1198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold716 (.A(net416),
    .X(net1199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold717 (.A(_0038_),
    .X(net1200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold718 (.A(net405),
    .X(net1201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold719 (.A(_0037_),
    .X(net1202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(net243),
    .X(net555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold720 (.A(\wbs_dat_delaybuff[19] ),
    .X(net1203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold721 (.A(\wbs_dat_delaybuff[17] ),
    .X(net1204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold722 (.A(\wbs_dat_delaybuff[23] ),
    .X(net1205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold723 (.A(net434),
    .X(net1206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold724 (.A(_0044_),
    .X(net1207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold725 (.A(net432),
    .X(net1208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold726 (.A(_0042_),
    .X(net1209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold727 (.A(\wbs_dat_delaybuff[1] ),
    .X(net1210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold728 (.A(\wbs_dat_delaybuff[6] ),
    .X(net1211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold729 (.A(\wbs_dat_delaybuff[0] ),
    .X(net1212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(net1115),
    .X(net556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold730 (.A(\wbs_dat_delaybuff[22] ),
    .X(net1213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold731 (.A(\wbs_dat_delaybuff[3] ),
    .X(net1214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold732 (.A(\wb_counter[26] ),
    .X(net1215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold733 (.A(\wbs_dat_delaybuff[4] ),
    .X(net1216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold734 (.A(_0074_),
    .X(net1217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold735 (.A(wbs_dat_i[12]),
    .X(net1218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold736 (.A(\wbs_dat_delaybuff[5] ),
    .X(net1219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold737 (.A(\wb_counter[4] ),
    .X(net1220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold738 (.A(\wb_counter[29] ),
    .X(net1221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold739 (.A(\wb_counter[18] ),
    .X(net1222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(net1117),
    .X(net557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold740 (.A(\wb_counter[28] ),
    .X(net1223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold741 (.A(wbs_dat_i[13]),
    .X(net1224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold742 (.A(\wb_counter[22] ),
    .X(net1225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold743 (.A(net404),
    .X(net1226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold744 (.A(\wb_counter[27] ),
    .X(net1227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold745 (.A(\wb_counter[17] ),
    .X(net1228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold746 (.A(wbs_adr_i[20]),
    .X(net1229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold747 (.A(\wb_counter[20] ),
    .X(net1230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold748 (.A(\wb_counter[30] ),
    .X(net1231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold749 (.A(\wb_counter[21] ),
    .X(net1232));
 sky130_fd_sc_hd__buf_12 hold75 (.A(net558),
    .X(la_data_out[39]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold750 (.A(net424),
    .X(net1233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold751 (.A(\wb_counter[8] ),
    .X(net1234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold752 (.A(\wb_counter[24] ),
    .X(net1235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold753 (.A(net428),
    .X(net1236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold754 (.A(\wb_counter[13] ),
    .X(net1237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold755 (.A(_0271_),
    .X(net1238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold756 (.A(\wb_counter[16] ),
    .X(net1239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold757 (.A(\wb_counter[14] ),
    .X(net1240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold758 (.A(\wb_counter[9] ),
    .X(net1241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold759 (.A(\wb_counter[12] ),
    .X(net1242));
 sky130_fd_sc_hd__buf_2 hold76 (.A(net592),
    .X(net559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold760 (.A(net429),
    .X(net1243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold761 (.A(net423),
    .X(net1244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold762 (.A(net422),
    .X(net1245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold763 (.A(net421),
    .X(net1246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold764 (.A(net406),
    .X(net1247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold765 (.A(net410),
    .X(net1248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold766 (.A(net436),
    .X(net1249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold767 (.A(net411),
    .X(net1250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold768 (.A(net418),
    .X(net1251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold769 (.A(net426),
    .X(net1252));
 sky130_fd_sc_hd__buf_2 hold77 (.A(net585),
    .X(net560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold770 (.A(net425),
    .X(net1253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold771 (.A(net412),
    .X(net1254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold772 (.A(net414),
    .X(net1255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold773 (.A(net435),
    .X(net1256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold774 (.A(net407),
    .X(net1257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold775 (.A(net420),
    .X(net1258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold776 (.A(net415),
    .X(net1259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold777 (.A(net417),
    .X(net1260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold778 (.A(net409),
    .X(net1261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold779 (.A(net413),
    .X(net1262));
 sky130_fd_sc_hd__buf_1 hold78 (.A(net320),
    .X(net561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold780 (.A(net408),
    .X(net1263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold781 (.A(net419),
    .X(net1264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold782 (.A(\wb_counter[10] ),
    .X(net1265));
 sky130_fd_sc_hd__buf_1 hold79 (.A(net395),
    .X(net562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(net932),
    .X(net491));
 sky130_fd_sc_hd__buf_12 hold80 (.A(net563),
    .X(la_data_out[4]));
 sky130_fd_sc_hd__buf_2 hold81 (.A(net590),
    .X(net564));
 sky130_fd_sc_hd__buf_2 hold82 (.A(_0117_),
    .X(net565));
 sky130_fd_sc_hd__buf_2 hold83 (.A(net454),
    .X(net566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(_0182_),
    .X(net567));
 sky130_fd_sc_hd__buf_1 hold85 (.A(net300),
    .X(net568));
 sky130_fd_sc_hd__buf_1 hold86 (.A(net373),
    .X(net569));
 sky130_fd_sc_hd__buf_12 hold87 (.A(net570),
    .X(la_data_out[1]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(net598),
    .X(net571));
 sky130_fd_sc_hd__clkbuf_2 hold89 (.A(_0114_),
    .X(net572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(net936),
    .X(net492));
 sky130_fd_sc_hd__clkbuf_2 hold90 (.A(_0116_),
    .X(net573));
 sky130_fd_sc_hd__clkbuf_2 hold91 (.A(net459),
    .X(net574));
 sky130_fd_sc_hd__buf_1 hold92 (.A(net311),
    .X(net575));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold93 (.A(net384),
    .X(net576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(net1139),
    .X(net577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(net1099),
    .X(net578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(net589),
    .X(net579));
 sky130_fd_sc_hd__clkbuf_2 hold97 (.A(net564),
    .X(net580));
 sky130_fd_sc_hd__buf_2 hold98 (.A(_0115_),
    .X(net581));
 sky130_fd_sc_hd__buf_1 hold99 (.A(net323),
    .X(net582));
 sky130_fd_sc_hd__clkbuf_8 input1 (.A(io_in_0),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(io_oeb_scrapcpu[17]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_2 input100 (.A(io_oeb_z80[33]),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_2 input101 (.A(io_oeb_z80[34]),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_2 input102 (.A(io_oeb_z80[35]),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_2 input103 (.A(io_oeb_z80[3]),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_2 input104 (.A(io_oeb_z80[4]),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_2 input105 (.A(io_oeb_z80[5]),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_2 input106 (.A(io_oeb_z80[6]),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_2 input107 (.A(io_oeb_z80[7]),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_2 input108 (.A(io_oeb_z80[8]),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_2 input109 (.A(io_oeb_z80[9]),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_2 input11 (.A(io_oeb_scrapcpu[18]),
    .X(net11));
 sky130_fd_sc_hd__buf_2 input110 (.A(io_out_scrapcpu[0]),
    .X(net110));
 sky130_fd_sc_hd__buf_2 input111 (.A(io_out_scrapcpu[10]),
    .X(net111));
 sky130_fd_sc_hd__buf_2 input112 (.A(io_out_scrapcpu[11]),
    .X(net112));
 sky130_fd_sc_hd__buf_2 input113 (.A(io_out_scrapcpu[12]),
    .X(net113));
 sky130_fd_sc_hd__buf_2 input114 (.A(io_out_scrapcpu[13]),
    .X(net114));
 sky130_fd_sc_hd__buf_2 input115 (.A(io_out_scrapcpu[14]),
    .X(net115));
 sky130_fd_sc_hd__buf_2 input116 (.A(io_out_scrapcpu[15]),
    .X(net116));
 sky130_fd_sc_hd__buf_2 input117 (.A(io_out_scrapcpu[16]),
    .X(net117));
 sky130_fd_sc_hd__buf_2 input118 (.A(io_out_scrapcpu[17]),
    .X(net118));
 sky130_fd_sc_hd__buf_2 input119 (.A(io_out_scrapcpu[18]),
    .X(net119));
 sky130_fd_sc_hd__clkbuf_2 input12 (.A(io_oeb_scrapcpu[19]),
    .X(net12));
 sky130_fd_sc_hd__buf_2 input120 (.A(io_out_scrapcpu[19]),
    .X(net120));
 sky130_fd_sc_hd__buf_2 input121 (.A(io_out_scrapcpu[1]),
    .X(net121));
 sky130_fd_sc_hd__buf_2 input122 (.A(io_out_scrapcpu[20]),
    .X(net122));
 sky130_fd_sc_hd__buf_2 input123 (.A(io_out_scrapcpu[21]),
    .X(net123));
 sky130_fd_sc_hd__buf_2 input124 (.A(io_out_scrapcpu[22]),
    .X(net124));
 sky130_fd_sc_hd__buf_2 input125 (.A(io_out_scrapcpu[23]),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_2 input126 (.A(io_out_scrapcpu[24]),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_2 input127 (.A(io_out_scrapcpu[25]),
    .X(net127));
 sky130_fd_sc_hd__clkbuf_2 input128 (.A(io_out_scrapcpu[26]),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_2 input129 (.A(io_out_scrapcpu[27]),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_2 input13 (.A(io_oeb_scrapcpu[1]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_2 input130 (.A(io_out_scrapcpu[28]),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_2 input131 (.A(io_out_scrapcpu[29]),
    .X(net131));
 sky130_fd_sc_hd__buf_2 input132 (.A(io_out_scrapcpu[2]),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_2 input133 (.A(io_out_scrapcpu[30]),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_2 input134 (.A(io_out_scrapcpu[31]),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_2 input135 (.A(io_out_scrapcpu[32]),
    .X(net135));
 sky130_fd_sc_hd__clkbuf_2 input136 (.A(io_out_scrapcpu[33]),
    .X(net136));
 sky130_fd_sc_hd__clkbuf_2 input137 (.A(io_out_scrapcpu[34]),
    .X(net137));
 sky130_fd_sc_hd__clkbuf_2 input138 (.A(io_out_scrapcpu[35]),
    .X(net138));
 sky130_fd_sc_hd__buf_2 input139 (.A(io_out_scrapcpu[3]),
    .X(net139));
 sky130_fd_sc_hd__clkbuf_2 input14 (.A(io_oeb_scrapcpu[20]),
    .X(net14));
 sky130_fd_sc_hd__buf_2 input140 (.A(io_out_scrapcpu[4]),
    .X(net140));
 sky130_fd_sc_hd__clkbuf_2 input141 (.A(io_out_scrapcpu[5]),
    .X(net141));
 sky130_fd_sc_hd__buf_2 input142 (.A(io_out_scrapcpu[6]),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_2 input143 (.A(io_out_scrapcpu[7]),
    .X(net143));
 sky130_fd_sc_hd__clkbuf_2 input144 (.A(io_out_scrapcpu[8]),
    .X(net144));
 sky130_fd_sc_hd__clkbuf_2 input145 (.A(io_out_scrapcpu[9]),
    .X(net145));
 sky130_fd_sc_hd__buf_4 input146 (.A(io_out_vliw[0]),
    .X(net146));
 sky130_fd_sc_hd__buf_4 input147 (.A(io_out_vliw[10]),
    .X(net147));
 sky130_fd_sc_hd__buf_4 input148 (.A(io_out_vliw[11]),
    .X(net148));
 sky130_fd_sc_hd__buf_4 input149 (.A(io_out_vliw[12]),
    .X(net149));
 sky130_fd_sc_hd__clkbuf_2 input15 (.A(io_oeb_scrapcpu[21]),
    .X(net15));
 sky130_fd_sc_hd__buf_4 input150 (.A(io_out_vliw[13]),
    .X(net150));
 sky130_fd_sc_hd__buf_4 input151 (.A(io_out_vliw[14]),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_4 input152 (.A(io_out_vliw[15]),
    .X(net152));
 sky130_fd_sc_hd__clkbuf_4 input153 (.A(io_out_vliw[16]),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_4 input154 (.A(io_out_vliw[17]),
    .X(net154));
 sky130_fd_sc_hd__clkbuf_4 input155 (.A(io_out_vliw[18]),
    .X(net155));
 sky130_fd_sc_hd__clkbuf_4 input156 (.A(io_out_vliw[19]),
    .X(net156));
 sky130_fd_sc_hd__buf_4 input157 (.A(io_out_vliw[1]),
    .X(net157));
 sky130_fd_sc_hd__clkbuf_4 input158 (.A(io_out_vliw[20]),
    .X(net158));
 sky130_fd_sc_hd__clkbuf_4 input159 (.A(io_out_vliw[21]),
    .X(net159));
 sky130_fd_sc_hd__clkbuf_2 input16 (.A(io_oeb_scrapcpu[22]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_4 input160 (.A(io_out_vliw[22]),
    .X(net160));
 sky130_fd_sc_hd__buf_2 input161 (.A(io_out_vliw[23]),
    .X(net161));
 sky130_fd_sc_hd__buf_2 input162 (.A(io_out_vliw[24]),
    .X(net162));
 sky130_fd_sc_hd__buf_2 input163 (.A(io_out_vliw[25]),
    .X(net163));
 sky130_fd_sc_hd__buf_2 input164 (.A(io_out_vliw[26]),
    .X(net164));
 sky130_fd_sc_hd__buf_2 input165 (.A(io_out_vliw[27]),
    .X(net165));
 sky130_fd_sc_hd__buf_2 input166 (.A(io_out_vliw[28]),
    .X(net166));
 sky130_fd_sc_hd__buf_2 input167 (.A(io_out_vliw[29]),
    .X(net167));
 sky130_fd_sc_hd__buf_4 input168 (.A(io_out_vliw[2]),
    .X(net168));
 sky130_fd_sc_hd__buf_2 input169 (.A(io_out_vliw[30]),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_2 input17 (.A(io_oeb_scrapcpu[23]),
    .X(net17));
 sky130_fd_sc_hd__buf_2 input170 (.A(io_out_vliw[31]),
    .X(net170));
 sky130_fd_sc_hd__buf_2 input171 (.A(io_out_vliw[32]),
    .X(net171));
 sky130_fd_sc_hd__buf_2 input172 (.A(io_out_vliw[33]),
    .X(net172));
 sky130_fd_sc_hd__buf_2 input173 (.A(io_out_vliw[34]),
    .X(net173));
 sky130_fd_sc_hd__clkbuf_2 input174 (.A(io_out_vliw[35]),
    .X(net174));
 sky130_fd_sc_hd__buf_4 input175 (.A(io_out_vliw[3]),
    .X(net175));
 sky130_fd_sc_hd__buf_4 input176 (.A(io_out_vliw[4]),
    .X(net176));
 sky130_fd_sc_hd__buf_4 input177 (.A(io_out_vliw[5]),
    .X(net177));
 sky130_fd_sc_hd__buf_4 input178 (.A(io_out_vliw[6]),
    .X(net178));
 sky130_fd_sc_hd__buf_4 input179 (.A(io_out_vliw[7]),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_2 input18 (.A(io_oeb_scrapcpu[24]),
    .X(net18));
 sky130_fd_sc_hd__buf_4 input180 (.A(io_out_vliw[8]),
    .X(net180));
 sky130_fd_sc_hd__buf_4 input181 (.A(io_out_vliw[9]),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_1 input182 (.A(io_out_z80[0]),
    .X(net182));
 sky130_fd_sc_hd__clkbuf_1 input183 (.A(io_out_z80[10]),
    .X(net183));
 sky130_fd_sc_hd__clkbuf_1 input184 (.A(io_out_z80[11]),
    .X(net184));
 sky130_fd_sc_hd__clkbuf_1 input185 (.A(io_out_z80[12]),
    .X(net185));
 sky130_fd_sc_hd__clkbuf_1 input186 (.A(io_out_z80[13]),
    .X(net186));
 sky130_fd_sc_hd__clkbuf_1 input187 (.A(io_out_z80[14]),
    .X(net187));
 sky130_fd_sc_hd__clkbuf_1 input188 (.A(io_out_z80[15]),
    .X(net188));
 sky130_fd_sc_hd__clkbuf_1 input189 (.A(io_out_z80[16]),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_2 input19 (.A(io_oeb_scrapcpu[25]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input190 (.A(io_out_z80[17]),
    .X(net190));
 sky130_fd_sc_hd__clkbuf_1 input191 (.A(io_out_z80[18]),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_1 input192 (.A(io_out_z80[19]),
    .X(net192));
 sky130_fd_sc_hd__clkbuf_1 input193 (.A(io_out_z80[1]),
    .X(net193));
 sky130_fd_sc_hd__clkbuf_1 input194 (.A(io_out_z80[20]),
    .X(net194));
 sky130_fd_sc_hd__clkbuf_1 input195 (.A(io_out_z80[21]),
    .X(net195));
 sky130_fd_sc_hd__clkbuf_1 input196 (.A(io_out_z80[22]),
    .X(net196));
 sky130_fd_sc_hd__clkbuf_1 input197 (.A(io_out_z80[23]),
    .X(net197));
 sky130_fd_sc_hd__clkbuf_1 input198 (.A(io_out_z80[24]),
    .X(net198));
 sky130_fd_sc_hd__clkbuf_1 input199 (.A(io_out_z80[25]),
    .X(net199));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(io_oeb_scrapcpu[0]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_2 input20 (.A(io_oeb_scrapcpu[26]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input200 (.A(io_out_z80[26]),
    .X(net200));
 sky130_fd_sc_hd__clkbuf_1 input201 (.A(io_out_z80[27]),
    .X(net201));
 sky130_fd_sc_hd__clkbuf_1 input202 (.A(io_out_z80[28]),
    .X(net202));
 sky130_fd_sc_hd__clkbuf_1 input203 (.A(io_out_z80[29]),
    .X(net203));
 sky130_fd_sc_hd__clkbuf_1 input204 (.A(io_out_z80[2]),
    .X(net204));
 sky130_fd_sc_hd__clkbuf_1 input205 (.A(io_out_z80[30]),
    .X(net205));
 sky130_fd_sc_hd__clkbuf_1 input206 (.A(io_out_z80[31]),
    .X(net206));
 sky130_fd_sc_hd__clkbuf_1 input207 (.A(io_out_z80[32]),
    .X(net207));
 sky130_fd_sc_hd__clkbuf_1 input208 (.A(io_out_z80[33]),
    .X(net208));
 sky130_fd_sc_hd__clkbuf_1 input209 (.A(io_out_z80[34]),
    .X(net209));
 sky130_fd_sc_hd__clkbuf_2 input21 (.A(io_oeb_scrapcpu[27]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input210 (.A(io_out_z80[35]),
    .X(net210));
 sky130_fd_sc_hd__clkbuf_1 input211 (.A(io_out_z80[3]),
    .X(net211));
 sky130_fd_sc_hd__clkbuf_1 input212 (.A(io_out_z80[4]),
    .X(net212));
 sky130_fd_sc_hd__clkbuf_1 input213 (.A(io_out_z80[5]),
    .X(net213));
 sky130_fd_sc_hd__clkbuf_1 input214 (.A(io_out_z80[6]),
    .X(net214));
 sky130_fd_sc_hd__clkbuf_1 input215 (.A(io_out_z80[7]),
    .X(net215));
 sky130_fd_sc_hd__clkbuf_1 input216 (.A(io_out_z80[8]),
    .X(net216));
 sky130_fd_sc_hd__clkbuf_1 input217 (.A(io_out_z80[9]),
    .X(net217));
 sky130_fd_sc_hd__dlymetal6s2s_1 input218 (.A(wb_rst_i),
    .X(net218));
 sky130_fd_sc_hd__buf_1 input219 (.A(net934),
    .X(net219));
 sky130_fd_sc_hd__clkbuf_2 input22 (.A(io_oeb_scrapcpu[28]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input220 (.A(net925),
    .X(net220));
 sky130_fd_sc_hd__clkbuf_1 input221 (.A(net931),
    .X(net221));
 sky130_fd_sc_hd__clkbuf_1 input222 (.A(net928),
    .X(net222));
 sky130_fd_sc_hd__clkbuf_1 input223 (.A(net1171),
    .X(net223));
 sky130_fd_sc_hd__clkbuf_1 input224 (.A(net946),
    .X(net224));
 sky130_fd_sc_hd__clkbuf_2 input225 (.A(net992),
    .X(net225));
 sky130_fd_sc_hd__clkbuf_2 input226 (.A(net986),
    .X(net226));
 sky130_fd_sc_hd__clkbuf_2 input227 (.A(net984),
    .X(net227));
 sky130_fd_sc_hd__clkbuf_2 input228 (.A(net1004),
    .X(net228));
 sky130_fd_sc_hd__buf_1 input229 (.A(net1000),
    .X(net229));
 sky130_fd_sc_hd__clkbuf_2 input23 (.A(io_oeb_scrapcpu[29]),
    .X(net23));
 sky130_fd_sc_hd__buf_1 input230 (.A(net1002),
    .X(net230));
 sky130_fd_sc_hd__clkbuf_2 input231 (.A(net998),
    .X(net231));
 sky130_fd_sc_hd__clkbuf_1 input232 (.A(net976),
    .X(net232));
 sky130_fd_sc_hd__clkbuf_1 input233 (.A(net973),
    .X(net233));
 sky130_fd_sc_hd__clkbuf_1 input234 (.A(net958),
    .X(net234));
 sky130_fd_sc_hd__clkbuf_1 input235 (.A(net940),
    .X(net235));
 sky130_fd_sc_hd__clkbuf_1 input236 (.A(net964),
    .X(net236));
 sky130_fd_sc_hd__clkbuf_1 input237 (.A(net967),
    .X(net237));
 sky130_fd_sc_hd__clkbuf_1 input238 (.A(net979),
    .X(net238));
 sky130_fd_sc_hd__clkbuf_1 input239 (.A(net961),
    .X(net239));
 sky130_fd_sc_hd__clkbuf_2 input24 (.A(io_oeb_scrapcpu[2]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input240 (.A(net970),
    .X(net240));
 sky130_fd_sc_hd__buf_1 input241 (.A(net988),
    .X(net241));
 sky130_fd_sc_hd__buf_1 input242 (.A(net1010),
    .X(net242));
 sky130_fd_sc_hd__buf_1 input243 (.A(net1014),
    .X(net243));
 sky130_fd_sc_hd__buf_1 input244 (.A(net1012),
    .X(net244));
 sky130_fd_sc_hd__buf_1 input245 (.A(net1008),
    .X(net245));
 sky130_fd_sc_hd__clkbuf_1 input246 (.A(net943),
    .X(net246));
 sky130_fd_sc_hd__buf_1 input247 (.A(net1006),
    .X(net247));
 sky130_fd_sc_hd__buf_1 input248 (.A(net996),
    .X(net248));
 sky130_fd_sc_hd__clkbuf_1 input249 (.A(net955),
    .X(net249));
 sky130_fd_sc_hd__clkbuf_2 input25 (.A(io_oeb_scrapcpu[30]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input250 (.A(net937),
    .X(net250));
 sky130_fd_sc_hd__clkbuf_1 input251 (.A(net952),
    .X(net251));
 sky130_fd_sc_hd__clkbuf_1 input252 (.A(net949),
    .X(net252));
 sky130_fd_sc_hd__clkbuf_2 input253 (.A(net982),
    .X(net253));
 sky130_fd_sc_hd__clkbuf_2 input254 (.A(net990),
    .X(net254));
 sky130_fd_sc_hd__clkbuf_2 input255 (.A(net994),
    .X(net255));
 sky130_fd_sc_hd__clkbuf_1 input256 (.A(wbs_stb_i),
    .X(net256));
 sky130_fd_sc_hd__buf_2 input257 (.A(net1178),
    .X(net257));
 sky130_fd_sc_hd__clkbuf_2 input26 (.A(io_oeb_scrapcpu[31]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_2 input27 (.A(io_oeb_scrapcpu[32]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_2 input28 (.A(io_oeb_scrapcpu[33]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_2 input29 (.A(io_oeb_scrapcpu[34]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_2 input3 (.A(io_oeb_scrapcpu[10]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_2 input30 (.A(io_oeb_scrapcpu[35]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_2 input31 (.A(io_oeb_scrapcpu[3]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_2 input32 (.A(io_oeb_scrapcpu[4]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_2 input33 (.A(io_oeb_scrapcpu[5]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_2 input34 (.A(io_oeb_scrapcpu[6]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_2 input35 (.A(io_oeb_scrapcpu[7]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_2 input36 (.A(io_oeb_scrapcpu[8]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_2 input37 (.A(io_oeb_scrapcpu[9]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 input38 (.A(io_oeb_vliw[0]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(io_oeb_vliw[10]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_2 input4 (.A(io_oeb_scrapcpu[11]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(io_oeb_vliw[11]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 input41 (.A(io_oeb_vliw[12]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 input42 (.A(io_oeb_vliw[13]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 input43 (.A(io_oeb_vliw[14]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(io_oeb_vliw[15]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(io_oeb_vliw[16]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 input46 (.A(io_oeb_vliw[17]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_1 input47 (.A(io_oeb_vliw[18]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 input48 (.A(io_oeb_vliw[19]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_1 input49 (.A(io_oeb_vliw[1]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_2 input5 (.A(io_oeb_scrapcpu[12]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input50 (.A(io_oeb_vliw[20]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 input51 (.A(io_oeb_vliw[21]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_1 input52 (.A(io_oeb_vliw[22]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 input53 (.A(io_oeb_vliw[23]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 input54 (.A(io_oeb_vliw[24]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_1 input55 (.A(io_oeb_vliw[25]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_1 input56 (.A(io_oeb_vliw[26]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_1 input57 (.A(io_oeb_vliw[27]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_1 input58 (.A(io_oeb_vliw[28]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 input59 (.A(io_oeb_vliw[29]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_2 input6 (.A(io_oeb_scrapcpu[13]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input60 (.A(io_oeb_vliw[2]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_1 input61 (.A(io_oeb_vliw[30]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 input62 (.A(io_oeb_vliw[31]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_1 input63 (.A(io_oeb_vliw[32]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_1 input64 (.A(io_oeb_vliw[33]),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_1 input65 (.A(io_oeb_vliw[34]),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_1 input66 (.A(io_oeb_vliw[35]),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_1 input67 (.A(io_oeb_vliw[3]),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_1 input68 (.A(io_oeb_vliw[4]),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_1 input69 (.A(io_oeb_vliw[5]),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_2 input7 (.A(io_oeb_scrapcpu[14]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input70 (.A(io_oeb_vliw[6]),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_1 input71 (.A(io_oeb_vliw[7]),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_1 input72 (.A(io_oeb_vliw[8]),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_1 input73 (.A(io_oeb_vliw[9]),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_2 input74 (.A(io_oeb_z80[0]),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_2 input75 (.A(io_oeb_z80[10]),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_2 input76 (.A(io_oeb_z80[11]),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_2 input77 (.A(io_oeb_z80[12]),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_2 input78 (.A(io_oeb_z80[13]),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_2 input79 (.A(io_oeb_z80[14]),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_2 input8 (.A(io_oeb_scrapcpu[15]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_2 input80 (.A(io_oeb_z80[15]),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_2 input81 (.A(io_oeb_z80[16]),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_2 input82 (.A(io_oeb_z80[17]),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_2 input83 (.A(io_oeb_z80[18]),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_2 input84 (.A(io_oeb_z80[19]),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_2 input85 (.A(io_oeb_z80[1]),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_2 input86 (.A(io_oeb_z80[20]),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_2 input87 (.A(io_oeb_z80[21]),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_2 input88 (.A(io_oeb_z80[22]),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_2 input89 (.A(io_oeb_z80[23]),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_2 input9 (.A(io_oeb_scrapcpu[16]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_2 input90 (.A(io_oeb_z80[24]),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_2 input91 (.A(io_oeb_z80[25]),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_2 input92 (.A(io_oeb_z80[26]),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_2 input93 (.A(io_oeb_z80[27]),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_2 input94 (.A(io_oeb_z80[28]),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_2 input95 (.A(io_oeb_z80[29]),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_2 input96 (.A(io_oeb_z80[2]),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_2 input97 (.A(io_oeb_z80[30]),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_2 input98 (.A(io_oeb_z80[31]),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_2 input99 (.A(io_oeb_z80[32]),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_8 max_cap449 (.A(net450),
    .X(net449));
 sky130_fd_sc_hd__clkbuf_8 max_cap450 (.A(net451),
    .X(net450));
 sky130_fd_sc_hd__clkbuf_8 max_cap451 (.A(net560),
    .X(net451));
 sky130_fd_sc_hd__conb_1 multiplexer_479 (.LO(net479));
 sky130_fd_sc_hd__conb_1 multiplexer_480 (.LO(net480));
 sky130_fd_sc_hd__conb_1 multiplexer_481 (.LO(net481));
 sky130_fd_sc_hd__conb_1 multiplexer_482 (.HI(net482));
 sky130_fd_sc_hd__conb_1 multiplexer_483 (.HI(net483));
 sky130_fd_sc_hd__buf_12 output258 (.A(net258),
    .X(custom_settings[0]));
 sky130_fd_sc_hd__buf_12 output259 (.A(net259),
    .X(custom_settings[10]));
 sky130_fd_sc_hd__buf_12 output260 (.A(net260),
    .X(custom_settings[11]));
 sky130_fd_sc_hd__buf_12 output261 (.A(net261),
    .X(custom_settings[12]));
 sky130_fd_sc_hd__buf_12 output262 (.A(net262),
    .X(custom_settings[13]));
 sky130_fd_sc_hd__buf_12 output263 (.A(net263),
    .X(custom_settings[14]));
 sky130_fd_sc_hd__buf_12 output264 (.A(net264),
    .X(custom_settings[15]));
 sky130_fd_sc_hd__buf_12 output265 (.A(net265),
    .X(custom_settings[16]));
 sky130_fd_sc_hd__buf_12 output266 (.A(net266),
    .X(custom_settings[17]));
 sky130_fd_sc_hd__buf_12 output267 (.A(net267),
    .X(custom_settings[18]));
 sky130_fd_sc_hd__buf_12 output268 (.A(net268),
    .X(custom_settings[19]));
 sky130_fd_sc_hd__buf_12 output269 (.A(net269),
    .X(custom_settings[1]));
 sky130_fd_sc_hd__buf_12 output270 (.A(net270),
    .X(custom_settings[20]));
 sky130_fd_sc_hd__buf_12 output271 (.A(net271),
    .X(custom_settings[21]));
 sky130_fd_sc_hd__buf_12 output272 (.A(net272),
    .X(custom_settings[22]));
 sky130_fd_sc_hd__buf_12 output273 (.A(net273),
    .X(custom_settings[23]));
 sky130_fd_sc_hd__buf_12 output274 (.A(net274),
    .X(custom_settings[24]));
 sky130_fd_sc_hd__buf_12 output275 (.A(net275),
    .X(custom_settings[25]));
 sky130_fd_sc_hd__buf_12 output276 (.A(net276),
    .X(custom_settings[26]));
 sky130_fd_sc_hd__buf_12 output277 (.A(net277),
    .X(custom_settings[27]));
 sky130_fd_sc_hd__buf_12 output278 (.A(net278),
    .X(custom_settings[28]));
 sky130_fd_sc_hd__buf_12 output279 (.A(net279),
    .X(custom_settings[29]));
 sky130_fd_sc_hd__buf_12 output280 (.A(net280),
    .X(custom_settings[2]));
 sky130_fd_sc_hd__buf_12 output281 (.A(net281),
    .X(custom_settings[30]));
 sky130_fd_sc_hd__buf_12 output282 (.A(net282),
    .X(custom_settings[31]));
 sky130_fd_sc_hd__buf_12 output283 (.A(net283),
    .X(custom_settings[3]));
 sky130_fd_sc_hd__buf_12 output284 (.A(net284),
    .X(custom_settings[4]));
 sky130_fd_sc_hd__buf_12 output285 (.A(net285),
    .X(custom_settings[5]));
 sky130_fd_sc_hd__buf_12 output286 (.A(net286),
    .X(custom_settings[6]));
 sky130_fd_sc_hd__buf_12 output287 (.A(net287),
    .X(custom_settings[7]));
 sky130_fd_sc_hd__buf_12 output288 (.A(net288),
    .X(custom_settings[8]));
 sky130_fd_sc_hd__buf_12 output289 (.A(net289),
    .X(custom_settings[9]));
 sky130_fd_sc_hd__buf_12 output290 (.A(net290),
    .X(io_oeb[10]));
 sky130_fd_sc_hd__buf_12 output291 (.A(net291),
    .X(io_oeb[11]));
 sky130_fd_sc_hd__buf_12 output292 (.A(net292),
    .X(io_oeb[12]));
 sky130_fd_sc_hd__buf_12 output293 (.A(net293),
    .X(io_oeb[13]));
 sky130_fd_sc_hd__buf_12 output294 (.A(net294),
    .X(io_oeb[14]));
 sky130_fd_sc_hd__buf_12 output295 (.A(net295),
    .X(io_oeb[15]));
 sky130_fd_sc_hd__buf_12 output296 (.A(net296),
    .X(io_oeb[16]));
 sky130_fd_sc_hd__buf_12 output297 (.A(net297),
    .X(io_oeb[17]));
 sky130_fd_sc_hd__buf_12 output298 (.A(net298),
    .X(io_oeb[18]));
 sky130_fd_sc_hd__buf_12 output299 (.A(net299),
    .X(io_oeb[19]));
 sky130_fd_sc_hd__buf_12 output300 (.A(net300),
    .X(io_oeb[1]));
 sky130_fd_sc_hd__buf_12 output301 (.A(net301),
    .X(io_oeb[20]));
 sky130_fd_sc_hd__buf_12 output302 (.A(net302),
    .X(io_oeb[21]));
 sky130_fd_sc_hd__buf_12 output303 (.A(net303),
    .X(io_oeb[22]));
 sky130_fd_sc_hd__buf_12 output304 (.A(net304),
    .X(io_oeb[23]));
 sky130_fd_sc_hd__buf_12 output305 (.A(net305),
    .X(io_oeb[24]));
 sky130_fd_sc_hd__buf_12 output306 (.A(net306),
    .X(io_oeb[25]));
 sky130_fd_sc_hd__buf_12 output307 (.A(net307),
    .X(io_oeb[26]));
 sky130_fd_sc_hd__buf_12 output308 (.A(net308),
    .X(io_oeb[27]));
 sky130_fd_sc_hd__buf_12 output309 (.A(net309),
    .X(io_oeb[28]));
 sky130_fd_sc_hd__buf_12 output310 (.A(net310),
    .X(io_oeb[29]));
 sky130_fd_sc_hd__buf_12 output311 (.A(net311),
    .X(io_oeb[2]));
 sky130_fd_sc_hd__buf_12 output312 (.A(net312),
    .X(io_oeb[30]));
 sky130_fd_sc_hd__buf_12 output313 (.A(net313),
    .X(io_oeb[31]));
 sky130_fd_sc_hd__buf_12 output314 (.A(net314),
    .X(io_oeb[32]));
 sky130_fd_sc_hd__buf_12 output315 (.A(net315),
    .X(io_oeb[33]));
 sky130_fd_sc_hd__buf_12 output316 (.A(net316),
    .X(io_oeb[34]));
 sky130_fd_sc_hd__buf_12 output317 (.A(net317),
    .X(io_oeb[35]));
 sky130_fd_sc_hd__buf_12 output318 (.A(net318),
    .X(io_oeb[36]));
 sky130_fd_sc_hd__buf_12 output319 (.A(net319),
    .X(io_oeb[37]));
 sky130_fd_sc_hd__buf_12 output320 (.A(net320),
    .X(io_oeb[4]));
 sky130_fd_sc_hd__buf_12 output321 (.A(net321),
    .X(io_oeb[5]));
 sky130_fd_sc_hd__buf_12 output322 (.A(net322),
    .X(io_oeb[6]));
 sky130_fd_sc_hd__buf_12 output323 (.A(net323),
    .X(io_oeb[7]));
 sky130_fd_sc_hd__buf_12 output324 (.A(net324),
    .X(io_oeb[8]));
 sky130_fd_sc_hd__buf_12 output325 (.A(net325),
    .X(io_oeb[9]));
 sky130_fd_sc_hd__buf_12 output326 (.A(net326),
    .X(io_out[10]));
 sky130_fd_sc_hd__buf_12 output327 (.A(net327),
    .X(io_out[11]));
 sky130_fd_sc_hd__buf_12 output328 (.A(net328),
    .X(io_out[12]));
 sky130_fd_sc_hd__buf_12 output329 (.A(net329),
    .X(io_out[13]));
 sky130_fd_sc_hd__buf_12 output330 (.A(net330),
    .X(io_out[14]));
 sky130_fd_sc_hd__buf_12 output331 (.A(net331),
    .X(io_out[15]));
 sky130_fd_sc_hd__buf_12 output332 (.A(net332),
    .X(io_out[16]));
 sky130_fd_sc_hd__buf_12 output333 (.A(net333),
    .X(io_out[17]));
 sky130_fd_sc_hd__buf_12 output334 (.A(net334),
    .X(io_out[18]));
 sky130_fd_sc_hd__buf_12 output335 (.A(net335),
    .X(io_out[19]));
 sky130_fd_sc_hd__buf_12 output336 (.A(net336),
    .X(io_out[1]));
 sky130_fd_sc_hd__buf_12 output337 (.A(net337),
    .X(io_out[20]));
 sky130_fd_sc_hd__buf_12 output338 (.A(net338),
    .X(io_out[21]));
 sky130_fd_sc_hd__buf_12 output339 (.A(net339),
    .X(io_out[22]));
 sky130_fd_sc_hd__buf_12 output340 (.A(net340),
    .X(io_out[23]));
 sky130_fd_sc_hd__buf_12 output341 (.A(net341),
    .X(io_out[24]));
 sky130_fd_sc_hd__buf_12 output342 (.A(net342),
    .X(io_out[25]));
 sky130_fd_sc_hd__buf_12 output343 (.A(net343),
    .X(io_out[26]));
 sky130_fd_sc_hd__buf_12 output344 (.A(net344),
    .X(io_out[27]));
 sky130_fd_sc_hd__buf_12 output345 (.A(net345),
    .X(io_out[28]));
 sky130_fd_sc_hd__buf_12 output346 (.A(net346),
    .X(io_out[29]));
 sky130_fd_sc_hd__buf_12 output347 (.A(net347),
    .X(io_out[2]));
 sky130_fd_sc_hd__buf_12 output348 (.A(net348),
    .X(io_out[30]));
 sky130_fd_sc_hd__buf_12 output349 (.A(net349),
    .X(io_out[31]));
 sky130_fd_sc_hd__buf_12 output350 (.A(net350),
    .X(io_out[32]));
 sky130_fd_sc_hd__buf_12 output351 (.A(net351),
    .X(io_out[33]));
 sky130_fd_sc_hd__buf_12 output352 (.A(net352),
    .X(io_out[34]));
 sky130_fd_sc_hd__buf_12 output353 (.A(net353),
    .X(io_out[35]));
 sky130_fd_sc_hd__buf_12 output354 (.A(net354),
    .X(io_out[36]));
 sky130_fd_sc_hd__buf_12 output355 (.A(net355),
    .X(io_out[37]));
 sky130_fd_sc_hd__buf_12 output356 (.A(net356),
    .X(io_out[3]));
 sky130_fd_sc_hd__buf_12 output357 (.A(net357),
    .X(io_out[4]));
 sky130_fd_sc_hd__buf_12 output358 (.A(net358),
    .X(io_out[5]));
 sky130_fd_sc_hd__buf_12 output359 (.A(net359),
    .X(io_out[6]));
 sky130_fd_sc_hd__buf_12 output360 (.A(net360),
    .X(io_out[7]));
 sky130_fd_sc_hd__buf_12 output361 (.A(net361),
    .X(io_out[8]));
 sky130_fd_sc_hd__buf_12 output362 (.A(net362),
    .X(io_out[9]));
 sky130_fd_sc_hd__buf_12 output363 (.A(net363),
    .X(la_data_out[10]));
 sky130_fd_sc_hd__buf_12 output364 (.A(net364),
    .X(la_data_out[11]));
 sky130_fd_sc_hd__buf_12 output365 (.A(net365),
    .X(la_data_out[12]));
 sky130_fd_sc_hd__buf_12 output366 (.A(net366),
    .X(la_data_out[13]));
 sky130_fd_sc_hd__buf_12 output367 (.A(net367),
    .X(la_data_out[14]));
 sky130_fd_sc_hd__buf_12 output368 (.A(net368),
    .X(la_data_out[15]));
 sky130_fd_sc_hd__buf_12 output369 (.A(net369),
    .X(la_data_out[16]));
 sky130_fd_sc_hd__buf_12 output370 (.A(net370),
    .X(la_data_out[17]));
 sky130_fd_sc_hd__buf_12 output371 (.A(net371),
    .X(la_data_out[18]));
 sky130_fd_sc_hd__buf_12 output372 (.A(net372),
    .X(la_data_out[19]));
 sky130_fd_sc_hd__buf_6 output373 (.A(net569),
    .X(net570));
 sky130_fd_sc_hd__buf_12 output374 (.A(net374),
    .X(la_data_out[20]));
 sky130_fd_sc_hd__buf_12 output375 (.A(net375),
    .X(la_data_out[21]));
 sky130_fd_sc_hd__buf_12 output376 (.A(net376),
    .X(la_data_out[22]));
 sky130_fd_sc_hd__buf_12 output377 (.A(net377),
    .X(la_data_out[23]));
 sky130_fd_sc_hd__buf_12 output378 (.A(net378),
    .X(la_data_out[24]));
 sky130_fd_sc_hd__buf_12 output379 (.A(net379),
    .X(la_data_out[25]));
 sky130_fd_sc_hd__buf_12 output380 (.A(net380),
    .X(la_data_out[26]));
 sky130_fd_sc_hd__buf_12 output381 (.A(net381),
    .X(la_data_out[27]));
 sky130_fd_sc_hd__buf_12 output382 (.A(net382),
    .X(la_data_out[28]));
 sky130_fd_sc_hd__buf_12 output383 (.A(net383),
    .X(la_data_out[29]));
 sky130_fd_sc_hd__buf_12 output384 (.A(net576),
    .X(la_data_out[2]));
 sky130_fd_sc_hd__buf_12 output385 (.A(net385),
    .X(la_data_out[30]));
 sky130_fd_sc_hd__buf_12 output386 (.A(net386),
    .X(la_data_out[31]));
 sky130_fd_sc_hd__buf_12 output387 (.A(net387),
    .X(la_data_out[32]));
 sky130_fd_sc_hd__buf_12 output388 (.A(net388),
    .X(la_data_out[33]));
 sky130_fd_sc_hd__buf_12 output389 (.A(net389),
    .X(la_data_out[34]));
 sky130_fd_sc_hd__buf_12 output390 (.A(net390),
    .X(la_data_out[35]));
 sky130_fd_sc_hd__buf_12 output391 (.A(net391),
    .X(la_data_out[36]));
 sky130_fd_sc_hd__buf_12 output392 (.A(net392),
    .X(la_data_out[37]));
 sky130_fd_sc_hd__buf_12 output393 (.A(net393),
    .X(la_data_out[38]));
 sky130_fd_sc_hd__buf_6 output394 (.A(net1118),
    .X(net558));
 sky130_fd_sc_hd__buf_6 output395 (.A(net562),
    .X(net563));
 sky130_fd_sc_hd__buf_12 output396 (.A(net396),
    .X(la_data_out[5]));
 sky130_fd_sc_hd__buf_12 output397 (.A(net397),
    .X(la_data_out[6]));
 sky130_fd_sc_hd__buf_12 output398 (.A(net398),
    .X(la_data_out[7]));
 sky130_fd_sc_hd__buf_12 output399 (.A(net399),
    .X(la_data_out[8]));
 sky130_fd_sc_hd__buf_12 output400 (.A(net400),
    .X(la_data_out[9]));
 sky130_fd_sc_hd__buf_12 output401 (.A(net401),
    .X(rst_scrapcpu));
 sky130_fd_sc_hd__buf_12 output402 (.A(net402),
    .X(rst_vliw));
 sky130_fd_sc_hd__buf_12 output403 (.A(net403),
    .X(rst_z80));
 sky130_fd_sc_hd__buf_12 output404 (.A(net923),
    .X(wbs_ack_o));
 sky130_fd_sc_hd__buf_12 output405 (.A(net830),
    .X(wbs_dat_o[0]));
 sky130_fd_sc_hd__buf_12 output406 (.A(net811),
    .X(wbs_dat_o[10]));
 sky130_fd_sc_hd__buf_12 output407 (.A(net730),
    .X(wbs_dat_o[11]));
 sky130_fd_sc_hd__buf_12 output408 (.A(net754),
    .X(wbs_dat_o[12]));
 sky130_fd_sc_hd__buf_12 output409 (.A(net757),
    .X(wbs_dat_o[13]));
 sky130_fd_sc_hd__buf_12 output410 (.A(net808),
    .X(wbs_dat_o[14]));
 sky130_fd_sc_hd__buf_12 output411 (.A(net766),
    .X(wbs_dat_o[15]));
 sky130_fd_sc_hd__buf_12 output412 (.A(net805),
    .X(wbs_dat_o[16]));
 sky130_fd_sc_hd__buf_12 output413 (.A(net781),
    .X(wbs_dat_o[17]));
 sky130_fd_sc_hd__buf_12 output414 (.A(net748),
    .X(wbs_dat_o[18]));
 sky130_fd_sc_hd__buf_12 output415 (.A(net760),
    .X(wbs_dat_o[19]));
 sky130_fd_sc_hd__buf_12 output416 (.A(net828),
    .X(wbs_dat_o[1]));
 sky130_fd_sc_hd__buf_12 output417 (.A(net775),
    .X(wbs_dat_o[20]));
 sky130_fd_sc_hd__buf_12 output418 (.A(net763),
    .X(wbs_dat_o[21]));
 sky130_fd_sc_hd__buf_12 output419 (.A(net778),
    .X(wbs_dat_o[22]));
 sky130_fd_sc_hd__buf_12 output420 (.A(net742),
    .X(wbs_dat_o[23]));
 sky130_fd_sc_hd__buf_12 output421 (.A(net772),
    .X(wbs_dat_o[24]));
 sky130_fd_sc_hd__buf_12 output422 (.A(net751),
    .X(wbs_dat_o[25]));
 sky130_fd_sc_hd__buf_12 output423 (.A(net784),
    .X(wbs_dat_o[26]));
 sky130_fd_sc_hd__buf_12 output424 (.A(net739),
    .X(wbs_dat_o[27]));
 sky130_fd_sc_hd__buf_12 output425 (.A(net798),
    .X(wbs_dat_o[28]));
 sky130_fd_sc_hd__buf_12 output426 (.A(net745),
    .X(wbs_dat_o[29]));
 sky130_fd_sc_hd__buf_12 output427 (.A(net826),
    .X(wbs_dat_o[2]));
 sky130_fd_sc_hd__buf_12 output428 (.A(net769),
    .X(wbs_dat_o[30]));
 sky130_fd_sc_hd__buf_12 output429 (.A(net736),
    .X(wbs_dat_o[31]));
 sky130_fd_sc_hd__buf_12 output430 (.A(net824),
    .X(wbs_dat_o[3]));
 sky130_fd_sc_hd__buf_12 output431 (.A(net835),
    .X(wbs_dat_o[4]));
 sky130_fd_sc_hd__buf_12 output432 (.A(net837),
    .X(wbs_dat_o[5]));
 sky130_fd_sc_hd__buf_12 output433 (.A(net839),
    .X(wbs_dat_o[6]));
 sky130_fd_sc_hd__buf_12 output434 (.A(net822),
    .X(wbs_dat_o[7]));
 sky130_fd_sc_hd__buf_12 output435 (.A(net790),
    .X(wbs_dat_o[8]));
 sky130_fd_sc_hd__buf_12 output436 (.A(net787),
    .X(wbs_dat_o[9]));
 assign io_oeb[0] = net482;
 assign io_oeb[3] = net479;
 assign io_out[0] = net480;
 assign la_data_out[0] = net483;
 assign la_data_out[3] = net481;
endmodule

