VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO vliw
  CLASS BLOCK ;
  FOREIGN vliw ;
  ORIGIN 0.000 0.000 ;
  SIZE 2200.000 BY 650.000 ;
  PIN cache_PC[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 36.890 646.000 37.170 650.000 ;
    END
  END cache_PC[0]
  PIN cache_PC[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 87.490 646.000 87.770 650.000 ;
    END
  END cache_PC[10]
  PIN cache_PC[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 92.550 646.000 92.830 650.000 ;
    END
  END cache_PC[11]
  PIN cache_PC[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 97.610 646.000 97.890 650.000 ;
    END
  END cache_PC[12]
  PIN cache_PC[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 102.670 646.000 102.950 650.000 ;
    END
  END cache_PC[13]
  PIN cache_PC[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 107.730 646.000 108.010 650.000 ;
    END
  END cache_PC[14]
  PIN cache_PC[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 112.790 646.000 113.070 650.000 ;
    END
  END cache_PC[15]
  PIN cache_PC[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 117.850 646.000 118.130 650.000 ;
    END
  END cache_PC[16]
  PIN cache_PC[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 122.910 646.000 123.190 650.000 ;
    END
  END cache_PC[17]
  PIN cache_PC[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 127.970 646.000 128.250 650.000 ;
    END
  END cache_PC[18]
  PIN cache_PC[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 133.030 646.000 133.310 650.000 ;
    END
  END cache_PC[19]
  PIN cache_PC[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 41.950 646.000 42.230 650.000 ;
    END
  END cache_PC[1]
  PIN cache_PC[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 138.090 646.000 138.370 650.000 ;
    END
  END cache_PC[20]
  PIN cache_PC[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 143.150 646.000 143.430 650.000 ;
    END
  END cache_PC[21]
  PIN cache_PC[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 148.210 646.000 148.490 650.000 ;
    END
  END cache_PC[22]
  PIN cache_PC[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 153.270 646.000 153.550 650.000 ;
    END
  END cache_PC[23]
  PIN cache_PC[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 158.330 646.000 158.610 650.000 ;
    END
  END cache_PC[24]
  PIN cache_PC[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 163.390 646.000 163.670 650.000 ;
    END
  END cache_PC[25]
  PIN cache_PC[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 168.450 646.000 168.730 650.000 ;
    END
  END cache_PC[26]
  PIN cache_PC[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 173.510 646.000 173.790 650.000 ;
    END
  END cache_PC[27]
  PIN cache_PC[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 47.010 646.000 47.290 650.000 ;
    END
  END cache_PC[2]
  PIN cache_PC[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 52.070 646.000 52.350 650.000 ;
    END
  END cache_PC[3]
  PIN cache_PC[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 57.130 646.000 57.410 650.000 ;
    END
  END cache_PC[4]
  PIN cache_PC[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 62.190 646.000 62.470 650.000 ;
    END
  END cache_PC[5]
  PIN cache_PC[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 67.250 646.000 67.530 650.000 ;
    END
  END cache_PC[6]
  PIN cache_PC[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 72.310 646.000 72.590 650.000 ;
    END
  END cache_PC[7]
  PIN cache_PC[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 77.370 646.000 77.650 650.000 ;
    END
  END cache_PC[8]
  PIN cache_PC[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 82.430 646.000 82.710 650.000 ;
    END
  END cache_PC[9]
  PIN cache_entry[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 178.570 646.000 178.850 650.000 ;
    END
  END cache_entry[0]
  PIN cache_entry[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 684.570 646.000 684.850 650.000 ;
    END
  END cache_entry[100]
  PIN cache_entry[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 689.630 646.000 689.910 650.000 ;
    END
  END cache_entry[101]
  PIN cache_entry[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 694.690 646.000 694.970 650.000 ;
    END
  END cache_entry[102]
  PIN cache_entry[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 699.750 646.000 700.030 650.000 ;
    END
  END cache_entry[103]
  PIN cache_entry[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 704.810 646.000 705.090 650.000 ;
    END
  END cache_entry[104]
  PIN cache_entry[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 709.870 646.000 710.150 650.000 ;
    END
  END cache_entry[105]
  PIN cache_entry[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 714.930 646.000 715.210 650.000 ;
    END
  END cache_entry[106]
  PIN cache_entry[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 719.990 646.000 720.270 650.000 ;
    END
  END cache_entry[107]
  PIN cache_entry[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 725.050 646.000 725.330 650.000 ;
    END
  END cache_entry[108]
  PIN cache_entry[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 730.110 646.000 730.390 650.000 ;
    END
  END cache_entry[109]
  PIN cache_entry[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 229.170 646.000 229.450 650.000 ;
    END
  END cache_entry[10]
  PIN cache_entry[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 3.912300 ;
    PORT
      LAYER met2 ;
        RECT 735.170 646.000 735.450 650.000 ;
    END
  END cache_entry[110]
  PIN cache_entry[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 740.230 646.000 740.510 650.000 ;
    END
  END cache_entry[111]
  PIN cache_entry[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 745.290 646.000 745.570 650.000 ;
    END
  END cache_entry[112]
  PIN cache_entry[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 750.350 646.000 750.630 650.000 ;
    END
  END cache_entry[113]
  PIN cache_entry[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 755.410 646.000 755.690 650.000 ;
    END
  END cache_entry[114]
  PIN cache_entry[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 760.470 646.000 760.750 650.000 ;
    END
  END cache_entry[115]
  PIN cache_entry[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 765.530 646.000 765.810 650.000 ;
    END
  END cache_entry[116]
  PIN cache_entry[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 770.590 646.000 770.870 650.000 ;
    END
  END cache_entry[117]
  PIN cache_entry[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 775.650 646.000 775.930 650.000 ;
    END
  END cache_entry[118]
  PIN cache_entry[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 780.710 646.000 780.990 650.000 ;
    END
  END cache_entry[119]
  PIN cache_entry[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 234.230 646.000 234.510 650.000 ;
    END
  END cache_entry[11]
  PIN cache_entry[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 785.770 646.000 786.050 650.000 ;
    END
  END cache_entry[120]
  PIN cache_entry[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 790.830 646.000 791.110 650.000 ;
    END
  END cache_entry[121]
  PIN cache_entry[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 795.890 646.000 796.170 650.000 ;
    END
  END cache_entry[122]
  PIN cache_entry[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 800.950 646.000 801.230 650.000 ;
    END
  END cache_entry[123]
  PIN cache_entry[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 806.010 646.000 806.290 650.000 ;
    END
  END cache_entry[124]
  PIN cache_entry[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 811.070 646.000 811.350 650.000 ;
    END
  END cache_entry[125]
  PIN cache_entry[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 816.130 646.000 816.410 650.000 ;
    END
  END cache_entry[126]
  PIN cache_entry[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 821.190 646.000 821.470 650.000 ;
    END
  END cache_entry[127]
  PIN cache_entry[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 239.290 646.000 239.570 650.000 ;
    END
  END cache_entry[12]
  PIN cache_entry[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 244.350 646.000 244.630 650.000 ;
    END
  END cache_entry[13]
  PIN cache_entry[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 249.410 646.000 249.690 650.000 ;
    END
  END cache_entry[14]
  PIN cache_entry[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 254.470 646.000 254.750 650.000 ;
    END
  END cache_entry[15]
  PIN cache_entry[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 259.530 646.000 259.810 650.000 ;
    END
  END cache_entry[16]
  PIN cache_entry[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 264.590 646.000 264.870 650.000 ;
    END
  END cache_entry[17]
  PIN cache_entry[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 269.650 646.000 269.930 650.000 ;
    END
  END cache_entry[18]
  PIN cache_entry[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 274.710 646.000 274.990 650.000 ;
    END
  END cache_entry[19]
  PIN cache_entry[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 183.630 646.000 183.910 650.000 ;
    END
  END cache_entry[1]
  PIN cache_entry[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 279.770 646.000 280.050 650.000 ;
    END
  END cache_entry[20]
  PIN cache_entry[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 284.830 646.000 285.110 650.000 ;
    END
  END cache_entry[21]
  PIN cache_entry[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 289.890 646.000 290.170 650.000 ;
    END
  END cache_entry[22]
  PIN cache_entry[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 294.950 646.000 295.230 650.000 ;
    END
  END cache_entry[23]
  PIN cache_entry[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 300.010 646.000 300.290 650.000 ;
    END
  END cache_entry[24]
  PIN cache_entry[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 305.070 646.000 305.350 650.000 ;
    END
  END cache_entry[25]
  PIN cache_entry[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 310.130 646.000 310.410 650.000 ;
    END
  END cache_entry[26]
  PIN cache_entry[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 315.190 646.000 315.470 650.000 ;
    END
  END cache_entry[27]
  PIN cache_entry[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 320.250 646.000 320.530 650.000 ;
    END
  END cache_entry[28]
  PIN cache_entry[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 325.310 646.000 325.590 650.000 ;
    END
  END cache_entry[29]
  PIN cache_entry[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met2 ;
        RECT 188.690 646.000 188.970 650.000 ;
    END
  END cache_entry[2]
  PIN cache_entry[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 330.370 646.000 330.650 650.000 ;
    END
  END cache_entry[30]
  PIN cache_entry[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 335.430 646.000 335.710 650.000 ;
    END
  END cache_entry[31]
  PIN cache_entry[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 340.490 646.000 340.770 650.000 ;
    END
  END cache_entry[32]
  PIN cache_entry[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 345.550 646.000 345.830 650.000 ;
    END
  END cache_entry[33]
  PIN cache_entry[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 350.610 646.000 350.890 650.000 ;
    END
  END cache_entry[34]
  PIN cache_entry[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 355.670 646.000 355.950 650.000 ;
    END
  END cache_entry[35]
  PIN cache_entry[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 360.730 646.000 361.010 650.000 ;
    END
  END cache_entry[36]
  PIN cache_entry[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 365.790 646.000 366.070 650.000 ;
    END
  END cache_entry[37]
  PIN cache_entry[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 370.850 646.000 371.130 650.000 ;
    END
  END cache_entry[38]
  PIN cache_entry[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 375.910 646.000 376.190 650.000 ;
    END
  END cache_entry[39]
  PIN cache_entry[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 193.750 646.000 194.030 650.000 ;
    END
  END cache_entry[3]
  PIN cache_entry[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 380.970 646.000 381.250 650.000 ;
    END
  END cache_entry[40]
  PIN cache_entry[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 386.030 646.000 386.310 650.000 ;
    END
  END cache_entry[41]
  PIN cache_entry[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 391.090 646.000 391.370 650.000 ;
    END
  END cache_entry[42]
  PIN cache_entry[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 396.150 646.000 396.430 650.000 ;
    END
  END cache_entry[43]
  PIN cache_entry[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 401.210 646.000 401.490 650.000 ;
    END
  END cache_entry[44]
  PIN cache_entry[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 406.270 646.000 406.550 650.000 ;
    END
  END cache_entry[45]
  PIN cache_entry[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 411.330 646.000 411.610 650.000 ;
    END
  END cache_entry[46]
  PIN cache_entry[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 416.390 646.000 416.670 650.000 ;
    END
  END cache_entry[47]
  PIN cache_entry[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 421.450 646.000 421.730 650.000 ;
    END
  END cache_entry[48]
  PIN cache_entry[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 426.510 646.000 426.790 650.000 ;
    END
  END cache_entry[49]
  PIN cache_entry[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 198.810 646.000 199.090 650.000 ;
    END
  END cache_entry[4]
  PIN cache_entry[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 431.570 646.000 431.850 650.000 ;
    END
  END cache_entry[50]
  PIN cache_entry[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 436.630 646.000 436.910 650.000 ;
    END
  END cache_entry[51]
  PIN cache_entry[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 441.690 646.000 441.970 650.000 ;
    END
  END cache_entry[52]
  PIN cache_entry[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 446.750 646.000 447.030 650.000 ;
    END
  END cache_entry[53]
  PIN cache_entry[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 451.810 646.000 452.090 650.000 ;
    END
  END cache_entry[54]
  PIN cache_entry[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 456.870 646.000 457.150 650.000 ;
    END
  END cache_entry[55]
  PIN cache_entry[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 461.930 646.000 462.210 650.000 ;
    END
  END cache_entry[56]
  PIN cache_entry[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 466.990 646.000 467.270 650.000 ;
    END
  END cache_entry[57]
  PIN cache_entry[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 472.050 646.000 472.330 650.000 ;
    END
  END cache_entry[58]
  PIN cache_entry[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 477.110 646.000 477.390 650.000 ;
    END
  END cache_entry[59]
  PIN cache_entry[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 203.870 646.000 204.150 650.000 ;
    END
  END cache_entry[5]
  PIN cache_entry[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 482.170 646.000 482.450 650.000 ;
    END
  END cache_entry[60]
  PIN cache_entry[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 487.230 646.000 487.510 650.000 ;
    END
  END cache_entry[61]
  PIN cache_entry[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 492.290 646.000 492.570 650.000 ;
    END
  END cache_entry[62]
  PIN cache_entry[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 497.350 646.000 497.630 650.000 ;
    END
  END cache_entry[63]
  PIN cache_entry[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 502.410 646.000 502.690 650.000 ;
    END
  END cache_entry[64]
  PIN cache_entry[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 507.470 646.000 507.750 650.000 ;
    END
  END cache_entry[65]
  PIN cache_entry[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 512.530 646.000 512.810 650.000 ;
    END
  END cache_entry[66]
  PIN cache_entry[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 517.590 646.000 517.870 650.000 ;
    END
  END cache_entry[67]
  PIN cache_entry[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 522.650 646.000 522.930 650.000 ;
    END
  END cache_entry[68]
  PIN cache_entry[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 527.710 646.000 527.990 650.000 ;
    END
  END cache_entry[69]
  PIN cache_entry[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 208.930 646.000 209.210 650.000 ;
    END
  END cache_entry[6]
  PIN cache_entry[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 532.770 646.000 533.050 650.000 ;
    END
  END cache_entry[70]
  PIN cache_entry[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 537.830 646.000 538.110 650.000 ;
    END
  END cache_entry[71]
  PIN cache_entry[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 542.890 646.000 543.170 650.000 ;
    END
  END cache_entry[72]
  PIN cache_entry[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 547.950 646.000 548.230 650.000 ;
    END
  END cache_entry[73]
  PIN cache_entry[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 553.010 646.000 553.290 650.000 ;
    END
  END cache_entry[74]
  PIN cache_entry[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 558.070 646.000 558.350 650.000 ;
    END
  END cache_entry[75]
  PIN cache_entry[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 563.130 646.000 563.410 650.000 ;
    END
  END cache_entry[76]
  PIN cache_entry[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 568.190 646.000 568.470 650.000 ;
    END
  END cache_entry[77]
  PIN cache_entry[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 573.250 646.000 573.530 650.000 ;
    END
  END cache_entry[78]
  PIN cache_entry[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 578.310 646.000 578.590 650.000 ;
    END
  END cache_entry[79]
  PIN cache_entry[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 213.990 646.000 214.270 650.000 ;
    END
  END cache_entry[7]
  PIN cache_entry[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 583.370 646.000 583.650 650.000 ;
    END
  END cache_entry[80]
  PIN cache_entry[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 588.430 646.000 588.710 650.000 ;
    END
  END cache_entry[81]
  PIN cache_entry[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 593.490 646.000 593.770 650.000 ;
    END
  END cache_entry[82]
  PIN cache_entry[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 598.550 646.000 598.830 650.000 ;
    END
  END cache_entry[83]
  PIN cache_entry[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 603.610 646.000 603.890 650.000 ;
    END
  END cache_entry[84]
  PIN cache_entry[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 608.670 646.000 608.950 650.000 ;
    END
  END cache_entry[85]
  PIN cache_entry[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 613.730 646.000 614.010 650.000 ;
    END
  END cache_entry[86]
  PIN cache_entry[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 618.790 646.000 619.070 650.000 ;
    END
  END cache_entry[87]
  PIN cache_entry[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 623.850 646.000 624.130 650.000 ;
    END
  END cache_entry[88]
  PIN cache_entry[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 628.910 646.000 629.190 650.000 ;
    END
  END cache_entry[89]
  PIN cache_entry[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 2.173500 ;
    PORT
      LAYER met2 ;
        RECT 219.050 646.000 219.330 650.000 ;
    END
  END cache_entry[8]
  PIN cache_entry[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 633.970 646.000 634.250 650.000 ;
    END
  END cache_entry[90]
  PIN cache_entry[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 639.030 646.000 639.310 650.000 ;
    END
  END cache_entry[91]
  PIN cache_entry[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 644.090 646.000 644.370 650.000 ;
    END
  END cache_entry[92]
  PIN cache_entry[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 649.150 646.000 649.430 650.000 ;
    END
  END cache_entry[93]
  PIN cache_entry[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 654.210 646.000 654.490 650.000 ;
    END
  END cache_entry[94]
  PIN cache_entry[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 659.270 646.000 659.550 650.000 ;
    END
  END cache_entry[95]
  PIN cache_entry[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 664.330 646.000 664.610 650.000 ;
    END
  END cache_entry[96]
  PIN cache_entry[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 669.390 646.000 669.670 650.000 ;
    END
  END cache_entry[97]
  PIN cache_entry[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 674.450 646.000 674.730 650.000 ;
    END
  END cache_entry[98]
  PIN cache_entry[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 679.510 646.000 679.790 650.000 ;
    END
  END cache_entry[99]
  PIN cache_entry[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 224.110 646.000 224.390 650.000 ;
    END
  END cache_entry[9]
  PIN cache_entry_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 165.960 2200.000 166.560 ;
    END
  END cache_entry_valid
  PIN cache_hit
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.363500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 161.880 2200.000 162.480 ;
    END
  END cache_hit
  PIN cache_invalidate
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 163.240 2200.000 163.840 ;
    END
  END cache_invalidate
  PIN cache_new_entry[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.363500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END cache_new_entry[0]
  PIN cache_new_entry[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.737000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 915.950 0.000 916.230 4.000 ;
    END
  END cache_new_entry[100]
  PIN cache_new_entry[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.737000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 924.690 0.000 924.970 4.000 ;
    END
  END cache_new_entry[101]
  PIN cache_new_entry[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.737000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 933.430 0.000 933.710 4.000 ;
    END
  END cache_new_entry[102]
  PIN cache_new_entry[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.737000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 942.170 0.000 942.450 4.000 ;
    END
  END cache_new_entry[103]
  PIN cache_new_entry[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.737000 ;
    ANTENNADIFFAREA 1.325700 ;
    PORT
      LAYER met2 ;
        RECT 950.910 0.000 951.190 4.000 ;
    END
  END cache_new_entry[104]
  PIN cache_new_entry[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.737000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 959.650 0.000 959.930 4.000 ;
    END
  END cache_new_entry[105]
  PIN cache_new_entry[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.737000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 968.390 0.000 968.670 4.000 ;
    END
  END cache_new_entry[106]
  PIN cache_new_entry[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.737000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 977.130 0.000 977.410 4.000 ;
    END
  END cache_new_entry[107]
  PIN cache_new_entry[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.737000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 985.870 0.000 986.150 4.000 ;
    END
  END cache_new_entry[108]
  PIN cache_new_entry[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.737000 ;
    ANTENNADIFFAREA 1.325700 ;
    PORT
      LAYER met2 ;
        RECT 994.610 0.000 994.890 4.000 ;
    END
  END cache_new_entry[109]
  PIN cache_new_entry[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.732500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 129.350 0.000 129.630 4.000 ;
    END
  END cache_new_entry[10]
  PIN cache_new_entry[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.621000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1003.350 0.000 1003.630 4.000 ;
    END
  END cache_new_entry[110]
  PIN cache_new_entry[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.994500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1012.090 0.000 1012.370 4.000 ;
    END
  END cache_new_entry[111]
  PIN cache_new_entry[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1020.830 0.000 1021.110 4.000 ;
    END
  END cache_new_entry[112]
  PIN cache_new_entry[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1029.570 0.000 1029.850 4.000 ;
    END
  END cache_new_entry[113]
  PIN cache_new_entry[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1038.310 0.000 1038.590 4.000 ;
    END
  END cache_new_entry[114]
  PIN cache_new_entry[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1047.050 0.000 1047.330 4.000 ;
    END
  END cache_new_entry[115]
  PIN cache_new_entry[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1055.790 0.000 1056.070 4.000 ;
    END
  END cache_new_entry[116]
  PIN cache_new_entry[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1064.530 0.000 1064.810 4.000 ;
    END
  END cache_new_entry[117]
  PIN cache_new_entry[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1073.270 0.000 1073.550 4.000 ;
    END
  END cache_new_entry[118]
  PIN cache_new_entry[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1082.010 0.000 1082.290 4.000 ;
    END
  END cache_new_entry[119]
  PIN cache_new_entry[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.732500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 138.090 0.000 138.370 4.000 ;
    END
  END cache_new_entry[11]
  PIN cache_new_entry[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1090.750 0.000 1091.030 4.000 ;
    END
  END cache_new_entry[120]
  PIN cache_new_entry[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1099.490 0.000 1099.770 4.000 ;
    END
  END cache_new_entry[121]
  PIN cache_new_entry[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1108.230 0.000 1108.510 4.000 ;
    END
  END cache_new_entry[122]
  PIN cache_new_entry[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1116.970 0.000 1117.250 4.000 ;
    END
  END cache_new_entry[123]
  PIN cache_new_entry[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1125.710 0.000 1125.990 4.000 ;
    END
  END cache_new_entry[124]
  PIN cache_new_entry[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1134.450 0.000 1134.730 4.000 ;
    END
  END cache_new_entry[125]
  PIN cache_new_entry[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1143.190 0.000 1143.470 4.000 ;
    END
  END cache_new_entry[126]
  PIN cache_new_entry[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1151.930 0.000 1152.210 4.000 ;
    END
  END cache_new_entry[127]
  PIN cache_new_entry[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.732500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 146.830 0.000 147.110 4.000 ;
    END
  END cache_new_entry[12]
  PIN cache_new_entry[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.732500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 155.570 0.000 155.850 4.000 ;
    END
  END cache_new_entry[13]
  PIN cache_new_entry[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 4.000 ;
    END
  END cache_new_entry[14]
  PIN cache_new_entry[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.673500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 173.050 0.000 173.330 4.000 ;
    END
  END cache_new_entry[15]
  PIN cache_new_entry[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.186500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 181.790 0.000 182.070 4.000 ;
    END
  END cache_new_entry[16]
  PIN cache_new_entry[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 190.530 0.000 190.810 4.000 ;
    END
  END cache_new_entry[17]
  PIN cache_new_entry[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.186500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 199.270 0.000 199.550 4.000 ;
    END
  END cache_new_entry[18]
  PIN cache_new_entry[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.732500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 208.010 0.000 208.290 4.000 ;
    END
  END cache_new_entry[19]
  PIN cache_new_entry[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.203000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 50.690 0.000 50.970 4.000 ;
    END
  END cache_new_entry[1]
  PIN cache_new_entry[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.732500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 216.750 0.000 217.030 4.000 ;
    END
  END cache_new_entry[20]
  PIN cache_new_entry[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.732500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 4.000 ;
    END
  END cache_new_entry[21]
  PIN cache_new_entry[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.732500 ;
    ANTENNADIFFAREA 1.325700 ;
    PORT
      LAYER met2 ;
        RECT 234.230 0.000 234.510 4.000 ;
    END
  END cache_new_entry[22]
  PIN cache_new_entry[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.732500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 242.970 0.000 243.250 4.000 ;
    END
  END cache_new_entry[23]
  PIN cache_new_entry[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.611000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 251.710 0.000 251.990 4.000 ;
    END
  END cache_new_entry[24]
  PIN cache_new_entry[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.611000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 260.450 0.000 260.730 4.000 ;
    END
  END cache_new_entry[25]
  PIN cache_new_entry[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 269.190 0.000 269.470 4.000 ;
    END
  END cache_new_entry[26]
  PIN cache_new_entry[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.203000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 277.930 0.000 278.210 4.000 ;
    END
  END cache_new_entry[27]
  PIN cache_new_entry[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.611000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 286.670 0.000 286.950 4.000 ;
    END
  END cache_new_entry[28]
  PIN cache_new_entry[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.611000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 295.410 0.000 295.690 4.000 ;
    END
  END cache_new_entry[29]
  PIN cache_new_entry[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.203000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 59.430 0.000 59.710 4.000 ;
    END
  END cache_new_entry[2]
  PIN cache_new_entry[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.203000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 304.150 0.000 304.430 4.000 ;
    END
  END cache_new_entry[30]
  PIN cache_new_entry[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.065000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 312.890 0.000 313.170 4.000 ;
    END
  END cache_new_entry[31]
  PIN cache_new_entry[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.149000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 321.630 0.000 321.910 4.000 ;
    END
  END cache_new_entry[32]
  PIN cache_new_entry[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.149000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 330.370 0.000 330.650 4.000 ;
    END
  END cache_new_entry[33]
  PIN cache_new_entry[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.011000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 339.110 0.000 339.390 4.000 ;
    END
  END cache_new_entry[34]
  PIN cache_new_entry[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.203000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 347.850 0.000 348.130 4.000 ;
    END
  END cache_new_entry[35]
  PIN cache_new_entry[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.203000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 356.590 0.000 356.870 4.000 ;
    END
  END cache_new_entry[36]
  PIN cache_new_entry[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.203000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 365.330 0.000 365.610 4.000 ;
    END
  END cache_new_entry[37]
  PIN cache_new_entry[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.203000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 374.070 0.000 374.350 4.000 ;
    END
  END cache_new_entry[38]
  PIN cache_new_entry[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.065000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 382.810 0.000 383.090 4.000 ;
    END
  END cache_new_entry[39]
  PIN cache_new_entry[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.149000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 68.170 0.000 68.450 4.000 ;
    END
  END cache_new_entry[3]
  PIN cache_new_entry[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.203000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 391.550 0.000 391.830 4.000 ;
    END
  END cache_new_entry[40]
  PIN cache_new_entry[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.203000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 400.290 0.000 400.570 4.000 ;
    END
  END cache_new_entry[41]
  PIN cache_new_entry[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.203000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 409.030 0.000 409.310 4.000 ;
    END
  END cache_new_entry[42]
  PIN cache_new_entry[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.203000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 417.770 0.000 418.050 4.000 ;
    END
  END cache_new_entry[43]
  PIN cache_new_entry[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.203000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 426.510 0.000 426.790 4.000 ;
    END
  END cache_new_entry[44]
  PIN cache_new_entry[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.203000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 435.250 0.000 435.530 4.000 ;
    END
  END cache_new_entry[45]
  PIN cache_new_entry[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.186500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 443.990 0.000 444.270 4.000 ;
    END
  END cache_new_entry[46]
  PIN cache_new_entry[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.203000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 452.730 0.000 453.010 4.000 ;
    END
  END cache_new_entry[47]
  PIN cache_new_entry[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.732500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 461.470 0.000 461.750 4.000 ;
    END
  END cache_new_entry[48]
  PIN cache_new_entry[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 470.210 0.000 470.490 4.000 ;
    END
  END cache_new_entry[49]
  PIN cache_new_entry[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.203000 ;
    ANTENNADIFFAREA 1.325700 ;
    PORT
      LAYER met2 ;
        RECT 76.910 0.000 77.190 4.000 ;
    END
  END cache_new_entry[4]
  PIN cache_new_entry[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.203000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 478.950 0.000 479.230 4.000 ;
    END
  END cache_new_entry[50]
  PIN cache_new_entry[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.203000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 487.690 0.000 487.970 4.000 ;
    END
  END cache_new_entry[51]
  PIN cache_new_entry[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 496.430 0.000 496.710 4.000 ;
    END
  END cache_new_entry[52]
  PIN cache_new_entry[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 505.170 0.000 505.450 4.000 ;
    END
  END cache_new_entry[53]
  PIN cache_new_entry[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.473000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 513.910 0.000 514.190 4.000 ;
    END
  END cache_new_entry[54]
  PIN cache_new_entry[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 522.650 0.000 522.930 4.000 ;
    END
  END cache_new_entry[55]
  PIN cache_new_entry[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.186500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 531.390 0.000 531.670 4.000 ;
    END
  END cache_new_entry[56]
  PIN cache_new_entry[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.186500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 540.130 0.000 540.410 4.000 ;
    END
  END cache_new_entry[57]
  PIN cache_new_entry[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.186500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 548.870 0.000 549.150 4.000 ;
    END
  END cache_new_entry[58]
  PIN cache_new_entry[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 557.610 0.000 557.890 4.000 ;
    END
  END cache_new_entry[59]
  PIN cache_new_entry[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.363500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 85.650 0.000 85.930 4.000 ;
    END
  END cache_new_entry[5]
  PIN cache_new_entry[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.203000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 566.350 0.000 566.630 4.000 ;
    END
  END cache_new_entry[60]
  PIN cache_new_entry[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.611000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 575.090 0.000 575.370 4.000 ;
    END
  END cache_new_entry[61]
  PIN cache_new_entry[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.203000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 583.830 0.000 584.110 4.000 ;
    END
  END cache_new_entry[62]
  PIN cache_new_entry[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.186500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 592.570 0.000 592.850 4.000 ;
    END
  END cache_new_entry[63]
  PIN cache_new_entry[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 601.310 0.000 601.590 4.000 ;
    END
  END cache_new_entry[64]
  PIN cache_new_entry[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.363500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 610.050 0.000 610.330 4.000 ;
    END
  END cache_new_entry[65]
  PIN cache_new_entry[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.363500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 618.790 0.000 619.070 4.000 ;
    END
  END cache_new_entry[66]
  PIN cache_new_entry[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 627.530 0.000 627.810 4.000 ;
    END
  END cache_new_entry[67]
  PIN cache_new_entry[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.363500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 636.270 0.000 636.550 4.000 ;
    END
  END cache_new_entry[68]
  PIN cache_new_entry[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.732500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 645.010 0.000 645.290 4.000 ;
    END
  END cache_new_entry[69]
  PIN cache_new_entry[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.149000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 94.390 0.000 94.670 4.000 ;
    END
  END cache_new_entry[6]
  PIN cache_new_entry[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.363500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 653.750 0.000 654.030 4.000 ;
    END
  END cache_new_entry[70]
  PIN cache_new_entry[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.363500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 662.490 0.000 662.770 4.000 ;
    END
  END cache_new_entry[71]
  PIN cache_new_entry[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.363500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 671.230 0.000 671.510 4.000 ;
    END
  END cache_new_entry[72]
  PIN cache_new_entry[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.363500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 679.970 0.000 680.250 4.000 ;
    END
  END cache_new_entry[73]
  PIN cache_new_entry[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.363500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 688.710 0.000 688.990 4.000 ;
    END
  END cache_new_entry[74]
  PIN cache_new_entry[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.363500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 697.450 0.000 697.730 4.000 ;
    END
  END cache_new_entry[75]
  PIN cache_new_entry[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 706.190 0.000 706.470 4.000 ;
    END
  END cache_new_entry[76]
  PIN cache_new_entry[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.363500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 714.930 0.000 715.210 4.000 ;
    END
  END cache_new_entry[77]
  PIN cache_new_entry[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.363500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 723.670 0.000 723.950 4.000 ;
    END
  END cache_new_entry[78]
  PIN cache_new_entry[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.363500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 732.410 0.000 732.690 4.000 ;
    END
  END cache_new_entry[79]
  PIN cache_new_entry[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.149000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END cache_new_entry[7]
  PIN cache_new_entry[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.455000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 741.150 0.000 741.430 4.000 ;
    END
  END cache_new_entry[80]
  PIN cache_new_entry[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 749.890 0.000 750.170 4.000 ;
    END
  END cache_new_entry[81]
  PIN cache_new_entry[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 758.630 0.000 758.910 4.000 ;
    END
  END cache_new_entry[82]
  PIN cache_new_entry[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 767.370 0.000 767.650 4.000 ;
    END
  END cache_new_entry[83]
  PIN cache_new_entry[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 776.110 0.000 776.390 4.000 ;
    END
  END cache_new_entry[84]
  PIN cache_new_entry[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.455000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 784.850 0.000 785.130 4.000 ;
    END
  END cache_new_entry[85]
  PIN cache_new_entry[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 793.590 0.000 793.870 4.000 ;
    END
  END cache_new_entry[86]
  PIN cache_new_entry[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 802.330 0.000 802.610 4.000 ;
    END
  END cache_new_entry[87]
  PIN cache_new_entry[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 811.070 0.000 811.350 4.000 ;
    END
  END cache_new_entry[88]
  PIN cache_new_entry[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 819.810 0.000 820.090 4.000 ;
    END
  END cache_new_entry[89]
  PIN cache_new_entry[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.732500 ;
    ANTENNADIFFAREA 1.760400 ;
    PORT
      LAYER met2 ;
        RECT 111.870 0.000 112.150 4.000 ;
    END
  END cache_new_entry[8]
  PIN cache_new_entry[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 828.550 0.000 828.830 4.000 ;
    END
  END cache_new_entry[90]
  PIN cache_new_entry[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 837.290 0.000 837.570 4.000 ;
    END
  END cache_new_entry[91]
  PIN cache_new_entry[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 846.030 0.000 846.310 4.000 ;
    END
  END cache_new_entry[92]
  PIN cache_new_entry[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 854.770 0.000 855.050 4.000 ;
    END
  END cache_new_entry[93]
  PIN cache_new_entry[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 863.510 0.000 863.790 4.000 ;
    END
  END cache_new_entry[94]
  PIN cache_new_entry[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 872.250 0.000 872.530 4.000 ;
    END
  END cache_new_entry[95]
  PIN cache_new_entry[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.737000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 880.990 0.000 881.270 4.000 ;
    END
  END cache_new_entry[96]
  PIN cache_new_entry[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.737000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 889.730 0.000 890.010 4.000 ;
    END
  END cache_new_entry[97]
  PIN cache_new_entry[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.737000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 898.470 0.000 898.750 4.000 ;
    END
  END cache_new_entry[98]
  PIN cache_new_entry[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.737000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 907.210 0.000 907.490 4.000 ;
    END
  END cache_new_entry[99]
  PIN cache_new_entry[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.732500 ;
    ANTENNADIFFAREA 1.325700 ;
    PORT
      LAYER met2 ;
        RECT 120.610 0.000 120.890 4.000 ;
    END
  END cache_new_entry[9]
  PIN cache_rst
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 164.600 2200.000 165.200 ;
    END
  END cache_rst
  PIN curr_PC[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.049000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 831.310 646.000 831.590 650.000 ;
    END
  END curr_PC[0]
  PIN curr_PC[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.852500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 881.910 646.000 882.190 650.000 ;
    END
  END curr_PC[10]
  PIN curr_PC[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.357500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 886.970 646.000 887.250 650.000 ;
    END
  END curr_PC[11]
  PIN curr_PC[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.431000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 892.030 646.000 892.310 650.000 ;
    END
  END curr_PC[12]
  PIN curr_PC[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.357500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 897.090 646.000 897.370 650.000 ;
    END
  END curr_PC[13]
  PIN curr_PC[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.855500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 902.150 646.000 902.430 650.000 ;
    END
  END curr_PC[14]
  PIN curr_PC[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.821000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 907.210 646.000 907.490 650.000 ;
    END
  END curr_PC[15]
  PIN curr_PC[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 912.270 646.000 912.550 650.000 ;
    END
  END curr_PC[16]
  PIN curr_PC[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.435500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 917.330 646.000 917.610 650.000 ;
    END
  END curr_PC[17]
  PIN curr_PC[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.483500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 922.390 646.000 922.670 650.000 ;
    END
  END curr_PC[18]
  PIN curr_PC[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.200000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 927.450 646.000 927.730 650.000 ;
    END
  END curr_PC[19]
  PIN curr_PC[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.049000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 836.370 646.000 836.650 650.000 ;
    END
  END curr_PC[1]
  PIN curr_PC[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.738500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 932.510 646.000 932.790 650.000 ;
    END
  END curr_PC[20]
  PIN curr_PC[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.326000 ;
    ANTENNADIFFAREA 1.760400 ;
    PORT
      LAYER met2 ;
        RECT 937.570 646.000 937.850 650.000 ;
    END
  END curr_PC[21]
  PIN curr_PC[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.113000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 942.630 646.000 942.910 650.000 ;
    END
  END curr_PC[22]
  PIN curr_PC[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.355000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 947.690 646.000 947.970 650.000 ;
    END
  END curr_PC[23]
  PIN curr_PC[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.365000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 952.750 646.000 953.030 650.000 ;
    END
  END curr_PC[24]
  PIN curr_PC[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.113000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 957.810 646.000 958.090 650.000 ;
    END
  END curr_PC[25]
  PIN curr_PC[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.239000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 962.870 646.000 963.150 650.000 ;
    END
  END curr_PC[26]
  PIN curr_PC[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.360500 ;
    ANTENNADIFFAREA 1.325700 ;
    PORT
      LAYER met2 ;
        RECT 967.930 646.000 968.210 650.000 ;
    END
  END curr_PC[27]
  PIN curr_PC[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.365000 ;
    ANTENNADIFFAREA 3.933900 ;
    PORT
      LAYER met2 ;
        RECT 841.430 646.000 841.710 650.000 ;
    END
  END curr_PC[2]
  PIN curr_PC[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.236000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 846.490 646.000 846.770 650.000 ;
    END
  END curr_PC[3]
  PIN curr_PC[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.857000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 851.550 646.000 851.830 650.000 ;
    END
  END curr_PC[4]
  PIN curr_PC[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.570500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 856.610 646.000 856.890 650.000 ;
    END
  END curr_PC[5]
  PIN curr_PC[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.357500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 861.670 646.000 861.950 650.000 ;
    END
  END curr_PC[6]
  PIN curr_PC[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.272000 ;
    ANTENNADIFFAREA 2.629800 ;
    PORT
      LAYER met2 ;
        RECT 866.730 646.000 867.010 650.000 ;
    END
  END curr_PC[7]
  PIN curr_PC[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.923000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 871.790 646.000 872.070 650.000 ;
    END
  END curr_PC[8]
  PIN curr_PC[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.675500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 876.850 646.000 877.130 650.000 ;
    END
  END curr_PC[9]
  PIN custom_settings[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 2122.070 0.000 2122.350 4.000 ;
    END
  END custom_settings[0]
  PIN custom_settings[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 2130.810 0.000 2131.090 4.000 ;
    END
  END custom_settings[1]
  PIN custom_settings[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.719500 ;
    PORT
      LAYER met2 ;
        RECT 2139.550 0.000 2139.830 4.000 ;
    END
  END custom_settings[2]
  PIN custom_settings[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.719500 ;
    PORT
      LAYER met2 ;
        RECT 2148.290 0.000 2148.570 4.000 ;
    END
  END custom_settings[3]
  PIN custom_settings[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 2157.030 0.000 2157.310 4.000 ;
    END
  END custom_settings[4]
  PIN dest_idx0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.469500 ;
    PORT
      LAYER met2 ;
        RECT 1195.630 646.000 1195.910 650.000 ;
    END
  END dest_idx0[0]
  PIN dest_idx0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.222000 ;
    PORT
      LAYER met2 ;
        RECT 1200.690 646.000 1200.970 650.000 ;
    END
  END dest_idx0[1]
  PIN dest_idx0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.372500 ;
    PORT
      LAYER met2 ;
        RECT 1205.750 646.000 1206.030 650.000 ;
    END
  END dest_idx0[2]
  PIN dest_idx0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.372500 ;
    PORT
      LAYER met2 ;
        RECT 1210.810 646.000 1211.090 650.000 ;
    END
  END dest_idx0[3]
  PIN dest_idx0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.372500 ;
    PORT
      LAYER met2 ;
        RECT 1215.870 646.000 1216.150 650.000 ;
    END
  END dest_idx0[4]
  PIN dest_idx1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.605500 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 227.160 2200.000 227.760 ;
    END
  END dest_idx1[0]
  PIN dest_idx1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.605500 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 228.520 2200.000 229.120 ;
    END
  END dest_idx1[1]
  PIN dest_idx1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.372500 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 229.880 2200.000 230.480 ;
    END
  END dest_idx1[2]
  PIN dest_idx1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.372500 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 231.240 2200.000 231.840 ;
    END
  END dest_idx1[3]
  PIN dest_idx1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.372500 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 232.600 2200.000 233.200 ;
    END
  END dest_idx1[4]
  PIN dest_idx2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.621000 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.800 4.000 124.400 ;
    END
  END dest_idx2[0]
  PIN dest_idx2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.520 4.000 127.120 ;
    END
  END dest_idx2[1]
  PIN dest_idx2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.621000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END dest_idx2[2]
  PIN dest_idx2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.621000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.960 4.000 132.560 ;
    END
  END dest_idx2[3]
  PIN dest_idx2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.621000 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.680 4.000 135.280 ;
    END
  END dest_idx2[4]
  PIN dest_mask0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met2 ;
        RECT 1185.510 646.000 1185.790 650.000 ;
    END
  END dest_mask0[0]
  PIN dest_mask0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1190.570 646.000 1190.850 650.000 ;
    END
  END dest_mask0[1]
  PIN dest_mask1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 224.440 2200.000 225.040 ;
    END
  END dest_mask1[0]
  PIN dest_mask1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 225.800 2200.000 226.400 ;
    END
  END dest_mask1[1]
  PIN dest_mask2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.360 4.000 118.960 ;
    END
  END dest_mask2[0]
  PIN dest_mask2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 5.651100 ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.080 4.000 121.680 ;
    END
  END dest_mask2[1]
  PIN dest_pred0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.499500 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met2 ;
        RECT 1236.110 646.000 1236.390 650.000 ;
    END
  END dest_pred0[0]
  PIN dest_pred0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.877500 ;
    ANTENNADIFFAREA 2.608200 ;
    PORT
      LAYER met2 ;
        RECT 1241.170 646.000 1241.450 650.000 ;
    END
  END dest_pred0[1]
  PIN dest_pred0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.877500 ;
    ANTENNADIFFAREA 2.608200 ;
    PORT
      LAYER met2 ;
        RECT 1246.230 646.000 1246.510 650.000 ;
    END
  END dest_pred0[2]
  PIN dest_pred1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.499500 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 238.040 2200.000 238.640 ;
    END
  END dest_pred1[0]
  PIN dest_pred1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.368000 ;
    ANTENNADIFFAREA 2.173500 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 239.400 2200.000 240.000 ;
    END
  END dest_pred1[1]
  PIN dest_pred1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.246500 ;
    ANTENNADIFFAREA 2.608200 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 240.760 2200.000 241.360 ;
    END
  END dest_pred1[2]
  PIN dest_pred2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.499500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.560 4.000 146.160 ;
    END
  END dest_pred2[0]
  PIN dest_pred2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.120500 ;
    ANTENNADIFFAREA 2.173500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.280 4.000 148.880 ;
    END
  END dest_pred2[1]
  PIN dest_pred2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.877500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.000 4.000 151.600 ;
    END
  END dest_pred2[2]
  PIN dest_pred_val0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.003500 ;
    ANTENNADIFFAREA 3.042900 ;
    PORT
      LAYER met2 ;
        RECT 1251.290 646.000 1251.570 650.000 ;
    END
  END dest_pred_val0
  PIN dest_pred_val1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.747000 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 242.120 2200.000 242.720 ;
    END
  END dest_pred_val1
  PIN dest_pred_val2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.125000 ;
    ANTENNADIFFAREA 5.651100 ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.720 4.000 154.320 ;
    END
  END dest_pred_val2
  PIN dest_val0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1023.590 646.000 1023.870 650.000 ;
    END
  END dest_val0[0]
  PIN dest_val0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1074.190 646.000 1074.470 650.000 ;
    END
  END dest_val0[10]
  PIN dest_val0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.673500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1079.250 646.000 1079.530 650.000 ;
    END
  END dest_val0[11]
  PIN dest_val0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1084.310 646.000 1084.590 650.000 ;
    END
  END dest_val0[12]
  PIN dest_val0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 1089.370 646.000 1089.650 650.000 ;
    END
  END dest_val0[13]
  PIN dest_val0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1094.430 646.000 1094.710 650.000 ;
    END
  END dest_val0[14]
  PIN dest_val0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 1099.490 646.000 1099.770 650.000 ;
    END
  END dest_val0[15]
  PIN dest_val0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met2 ;
        RECT 1104.550 646.000 1104.830 650.000 ;
    END
  END dest_val0[16]
  PIN dest_val0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.673500 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met2 ;
        RECT 1109.610 646.000 1109.890 650.000 ;
    END
  END dest_val0[17]
  PIN dest_val0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.921000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1114.670 646.000 1114.950 650.000 ;
    END
  END dest_val0[18]
  PIN dest_val0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1119.730 646.000 1120.010 650.000 ;
    END
  END dest_val0[19]
  PIN dest_val0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1028.650 646.000 1028.930 650.000 ;
    END
  END dest_val0[1]
  PIN dest_val0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1124.790 646.000 1125.070 650.000 ;
    END
  END dest_val0[20]
  PIN dest_val0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.921000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1129.850 646.000 1130.130 650.000 ;
    END
  END dest_val0[21]
  PIN dest_val0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 1134.910 646.000 1135.190 650.000 ;
    END
  END dest_val0[22]
  PIN dest_val0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 1139.970 646.000 1140.250 650.000 ;
    END
  END dest_val0[23]
  PIN dest_val0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 1145.030 646.000 1145.310 650.000 ;
    END
  END dest_val0[24]
  PIN dest_val0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 1150.090 646.000 1150.370 650.000 ;
    END
  END dest_val0[25]
  PIN dest_val0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 1155.150 646.000 1155.430 650.000 ;
    END
  END dest_val0[26]
  PIN dest_val0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 1160.210 646.000 1160.490 650.000 ;
    END
  END dest_val0[27]
  PIN dest_val0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.921000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1165.270 646.000 1165.550 650.000 ;
    END
  END dest_val0[28]
  PIN dest_val0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1170.330 646.000 1170.610 650.000 ;
    END
  END dest_val0[29]
  PIN dest_val0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1033.710 646.000 1033.990 650.000 ;
    END
  END dest_val0[2]
  PIN dest_val0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 1175.390 646.000 1175.670 650.000 ;
    END
  END dest_val0[30]
  PIN dest_val0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 1180.450 646.000 1180.730 650.000 ;
    END
  END dest_val0[31]
  PIN dest_val0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1038.770 646.000 1039.050 650.000 ;
    END
  END dest_val0[3]
  PIN dest_val0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1043.830 646.000 1044.110 650.000 ;
    END
  END dest_val0[4]
  PIN dest_val0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1048.890 646.000 1049.170 650.000 ;
    END
  END dest_val0[5]
  PIN dest_val0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1053.950 646.000 1054.230 650.000 ;
    END
  END dest_val0[6]
  PIN dest_val0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1059.010 646.000 1059.290 650.000 ;
    END
  END dest_val0[7]
  PIN dest_val0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1064.070 646.000 1064.350 650.000 ;
    END
  END dest_val0[8]
  PIN dest_val0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1069.130 646.000 1069.410 650.000 ;
    END
  END dest_val0[9]
  PIN dest_val1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 180.920 2200.000 181.520 ;
    END
  END dest_val1[0]
  PIN dest_val1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 194.520 2200.000 195.120 ;
    END
  END dest_val1[10]
  PIN dest_val1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 195.880 2200.000 196.480 ;
    END
  END dest_val1[11]
  PIN dest_val1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 197.240 2200.000 197.840 ;
    END
  END dest_val1[12]
  PIN dest_val1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.460500 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 198.600 2200.000 199.200 ;
    END
  END dest_val1[13]
  PIN dest_val1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 199.960 2200.000 200.560 ;
    END
  END dest_val1[14]
  PIN dest_val1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.460500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 201.320 2200.000 201.920 ;
    END
  END dest_val1[15]
  PIN dest_val1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.673500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 202.680 2200.000 203.280 ;
    END
  END dest_val1[16]
  PIN dest_val1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.708000 ;
    ANTENNADIFFAREA 2.608200 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 204.040 2200.000 204.640 ;
    END
  END dest_val1[17]
  PIN dest_val1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 205.400 2200.000 206.000 ;
    END
  END dest_val1[18]
  PIN dest_val1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 206.760 2200.000 207.360 ;
    END
  END dest_val1[19]
  PIN dest_val1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 182.280 2200.000 182.880 ;
    END
  END dest_val1[1]
  PIN dest_val1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.639000 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 208.120 2200.000 208.720 ;
    END
  END dest_val1[20]
  PIN dest_val1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 209.480 2200.000 210.080 ;
    END
  END dest_val1[21]
  PIN dest_val1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 210.840 2200.000 211.440 ;
    END
  END dest_val1[22]
  PIN dest_val1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 212.200 2200.000 212.800 ;
    END
  END dest_val1[23]
  PIN dest_val1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 213.560 2200.000 214.160 ;
    END
  END dest_val1[24]
  PIN dest_val1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 214.920 2200.000 215.520 ;
    END
  END dest_val1[25]
  PIN dest_val1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.673500 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 216.280 2200.000 216.880 ;
    END
  END dest_val1[26]
  PIN dest_val1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 217.640 2200.000 218.240 ;
    END
  END dest_val1[27]
  PIN dest_val1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 219.000 2200.000 219.600 ;
    END
  END dest_val1[28]
  PIN dest_val1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.673500 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 220.360 2200.000 220.960 ;
    END
  END dest_val1[29]
  PIN dest_val1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 183.640 2200.000 184.240 ;
    END
  END dest_val1[2]
  PIN dest_val1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.673500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 221.720 2200.000 222.320 ;
    END
  END dest_val1[30]
  PIN dest_val1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 223.080 2200.000 223.680 ;
    END
  END dest_val1[31]
  PIN dest_val1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 185.000 2200.000 185.600 ;
    END
  END dest_val1[3]
  PIN dest_val1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 186.360 2200.000 186.960 ;
    END
  END dest_val1[4]
  PIN dest_val1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 187.720 2200.000 188.320 ;
    END
  END dest_val1[5]
  PIN dest_val1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 189.080 2200.000 189.680 ;
    END
  END dest_val1[6]
  PIN dest_val1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 190.440 2200.000 191.040 ;
    END
  END dest_val1[7]
  PIN dest_val1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 191.800 2200.000 192.400 ;
    END
  END dest_val1[8]
  PIN dest_val1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.639000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 193.160 2200.000 193.760 ;
    END
  END dest_val1[9]
  PIN dest_val2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.485000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.320 4.000 31.920 ;
    END
  END dest_val2[0]
  PIN dest_val2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 58.520 4.000 59.120 ;
    END
  END dest_val2[10]
  PIN dest_val2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END dest_val2[11]
  PIN dest_val2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.960 4.000 64.560 ;
    END
  END dest_val2[12]
  PIN dest_val2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.680 4.000 67.280 ;
    END
  END dest_val2[13]
  PIN dest_val2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.400 4.000 70.000 ;
    END
  END dest_val2[14]
  PIN dest_val2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.120 4.000 72.720 ;
    END
  END dest_val2[15]
  PIN dest_val2[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.485000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END dest_val2[16]
  PIN dest_val2[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 77.560 4.000 78.160 ;
    END
  END dest_val2[17]
  PIN dest_val2[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.485000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.280 4.000 80.880 ;
    END
  END dest_val2[18]
  PIN dest_val2[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 4.000 83.600 ;
    END
  END dest_val2[19]
  PIN dest_val2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.485000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END dest_val2[1]
  PIN dest_val2[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.485000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.720 4.000 86.320 ;
    END
  END dest_val2[20]
  PIN dest_val2[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.485000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END dest_val2[21]
  PIN dest_val2[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.485000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.160 4.000 91.760 ;
    END
  END dest_val2[22]
  PIN dest_val2[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.880 4.000 94.480 ;
    END
  END dest_val2[23]
  PIN dest_val2[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.485000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.600 4.000 97.200 ;
    END
  END dest_val2[24]
  PIN dest_val2[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.485000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 99.320 4.000 99.920 ;
    END
  END dest_val2[25]
  PIN dest_val2[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.485000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END dest_val2[26]
  PIN dest_val2[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.485000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.760 4.000 105.360 ;
    END
  END dest_val2[27]
  PIN dest_val2[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.485000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 107.480 4.000 108.080 ;
    END
  END dest_val2[28]
  PIN dest_val2[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.485000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.200 4.000 110.800 ;
    END
  END dest_val2[29]
  PIN dest_val2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.760 4.000 37.360 ;
    END
  END dest_val2[2]
  PIN dest_val2[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.485000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.920 4.000 113.520 ;
    END
  END dest_val2[30]
  PIN dest_val2[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.485000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END dest_val2[31]
  PIN dest_val2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.485000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 4.000 40.080 ;
    END
  END dest_val2[3]
  PIN dest_val2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.485000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.200 4.000 42.800 ;
    END
  END dest_val2[4]
  PIN dest_val2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.920 4.000 45.520 ;
    END
  END dest_val2[5]
  PIN dest_val2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END dest_val2[6]
  PIN dest_val2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.485000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.360 4.000 50.960 ;
    END
  END dest_val2[7]
  PIN dest_val2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.080 4.000 53.680 ;
    END
  END dest_val2[8]
  PIN dest_val2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 4.000 56.400 ;
    END
  END dest_val2[9]
  PIN eu0_busy
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1615.610 646.000 1615.890 650.000 ;
    END
  END eu0_busy
  PIN eu0_instruction[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1620.670 646.000 1620.950 650.000 ;
    END
  END eu0_instruction[0]
  PIN eu0_instruction[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 10.454400 ;
    PORT
      LAYER met2 ;
        RECT 1671.270 646.000 1671.550 650.000 ;
    END
  END eu0_instruction[10]
  PIN eu0_instruction[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1676.330 646.000 1676.610 650.000 ;
    END
  END eu0_instruction[11]
  PIN eu0_instruction[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 10.454400 ;
    PORT
      LAYER met2 ;
        RECT 1681.390 646.000 1681.670 650.000 ;
    END
  END eu0_instruction[12]
  PIN eu0_instruction[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1686.450 646.000 1686.730 650.000 ;
    END
  END eu0_instruction[13]
  PIN eu0_instruction[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1691.510 646.000 1691.790 650.000 ;
    END
  END eu0_instruction[14]
  PIN eu0_instruction[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1696.570 646.000 1696.850 650.000 ;
    END
  END eu0_instruction[15]
  PIN eu0_instruction[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1701.630 646.000 1701.910 650.000 ;
    END
  END eu0_instruction[16]
  PIN eu0_instruction[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1706.690 646.000 1706.970 650.000 ;
    END
  END eu0_instruction[17]
  PIN eu0_instruction[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1711.750 646.000 1712.030 650.000 ;
    END
  END eu0_instruction[18]
  PIN eu0_instruction[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1716.810 646.000 1717.090 650.000 ;
    END
  END eu0_instruction[19]
  PIN eu0_instruction[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 10.454400 ;
    PORT
      LAYER met2 ;
        RECT 1625.730 646.000 1626.010 650.000 ;
    END
  END eu0_instruction[1]
  PIN eu0_instruction[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1721.870 646.000 1722.150 650.000 ;
    END
  END eu0_instruction[20]
  PIN eu0_instruction[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1726.930 646.000 1727.210 650.000 ;
    END
  END eu0_instruction[21]
  PIN eu0_instruction[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1731.990 646.000 1732.270 650.000 ;
    END
  END eu0_instruction[22]
  PIN eu0_instruction[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1737.050 646.000 1737.330 650.000 ;
    END
  END eu0_instruction[23]
  PIN eu0_instruction[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1742.110 646.000 1742.390 650.000 ;
    END
  END eu0_instruction[24]
  PIN eu0_instruction[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1747.170 646.000 1747.450 650.000 ;
    END
  END eu0_instruction[25]
  PIN eu0_instruction[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1752.230 646.000 1752.510 650.000 ;
    END
  END eu0_instruction[26]
  PIN eu0_instruction[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1757.290 646.000 1757.570 650.000 ;
    END
  END eu0_instruction[27]
  PIN eu0_instruction[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1762.350 646.000 1762.630 650.000 ;
    END
  END eu0_instruction[28]
  PIN eu0_instruction[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1767.410 646.000 1767.690 650.000 ;
    END
  END eu0_instruction[29]
  PIN eu0_instruction[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 10.454400 ;
    PORT
      LAYER met2 ;
        RECT 1630.790 646.000 1631.070 650.000 ;
    END
  END eu0_instruction[2]
  PIN eu0_instruction[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1772.470 646.000 1772.750 650.000 ;
    END
  END eu0_instruction[30]
  PIN eu0_instruction[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1777.530 646.000 1777.810 650.000 ;
    END
  END eu0_instruction[31]
  PIN eu0_instruction[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1782.590 646.000 1782.870 650.000 ;
    END
  END eu0_instruction[32]
  PIN eu0_instruction[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1787.650 646.000 1787.930 650.000 ;
    END
  END eu0_instruction[33]
  PIN eu0_instruction[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1792.710 646.000 1792.990 650.000 ;
    END
  END eu0_instruction[34]
  PIN eu0_instruction[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1797.770 646.000 1798.050 650.000 ;
    END
  END eu0_instruction[35]
  PIN eu0_instruction[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1802.830 646.000 1803.110 650.000 ;
    END
  END eu0_instruction[36]
  PIN eu0_instruction[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1807.890 646.000 1808.170 650.000 ;
    END
  END eu0_instruction[37]
  PIN eu0_instruction[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1812.950 646.000 1813.230 650.000 ;
    END
  END eu0_instruction[38]
  PIN eu0_instruction[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1818.010 646.000 1818.290 650.000 ;
    END
  END eu0_instruction[39]
  PIN eu0_instruction[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 10.454400 ;
    PORT
      LAYER met2 ;
        RECT 1635.850 646.000 1636.130 650.000 ;
    END
  END eu0_instruction[3]
  PIN eu0_instruction[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1823.070 646.000 1823.350 650.000 ;
    END
  END eu0_instruction[40]
  PIN eu0_instruction[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1828.130 646.000 1828.410 650.000 ;
    END
  END eu0_instruction[41]
  PIN eu0_instruction[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 15.670799 ;
    PORT
      LAYER met2 ;
        RECT 1640.910 646.000 1641.190 650.000 ;
    END
  END eu0_instruction[4]
  PIN eu0_instruction[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 10.454400 ;
    PORT
      LAYER met2 ;
        RECT 1645.970 646.000 1646.250 650.000 ;
    END
  END eu0_instruction[5]
  PIN eu0_instruction[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 10.454400 ;
    PORT
      LAYER met2 ;
        RECT 1651.030 646.000 1651.310 650.000 ;
    END
  END eu0_instruction[6]
  PIN eu0_instruction[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 10.454400 ;
    PORT
      LAYER met2 ;
        RECT 1656.090 646.000 1656.370 650.000 ;
    END
  END eu0_instruction[7]
  PIN eu0_instruction[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 20.887199 ;
    PORT
      LAYER met2 ;
        RECT 1661.150 646.000 1661.430 650.000 ;
    END
  END eu0_instruction[8]
  PIN eu0_instruction[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 20.887199 ;
    PORT
      LAYER met2 ;
        RECT 1666.210 646.000 1666.490 650.000 ;
    END
  END eu0_instruction[9]
  PIN eu1_busy
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 340.040 2200.000 340.640 ;
    END
  END eu1_busy
  PIN eu1_instruction[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 341.400 2200.000 342.000 ;
    END
  END eu1_instruction[0]
  PIN eu1_instruction[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 355.000 2200.000 355.600 ;
    END
  END eu1_instruction[10]
  PIN eu1_instruction[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 356.360 2200.000 356.960 ;
    END
  END eu1_instruction[11]
  PIN eu1_instruction[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 357.720 2200.000 358.320 ;
    END
  END eu1_instruction[12]
  PIN eu1_instruction[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 359.080 2200.000 359.680 ;
    END
  END eu1_instruction[13]
  PIN eu1_instruction[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 360.440 2200.000 361.040 ;
    END
  END eu1_instruction[14]
  PIN eu1_instruction[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 361.800 2200.000 362.400 ;
    END
  END eu1_instruction[15]
  PIN eu1_instruction[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 363.160 2200.000 363.760 ;
    END
  END eu1_instruction[16]
  PIN eu1_instruction[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 364.520 2200.000 365.120 ;
    END
  END eu1_instruction[17]
  PIN eu1_instruction[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 365.880 2200.000 366.480 ;
    END
  END eu1_instruction[18]
  PIN eu1_instruction[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 367.240 2200.000 367.840 ;
    END
  END eu1_instruction[19]
  PIN eu1_instruction[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 342.760 2200.000 343.360 ;
    END
  END eu1_instruction[1]
  PIN eu1_instruction[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 368.600 2200.000 369.200 ;
    END
  END eu1_instruction[20]
  PIN eu1_instruction[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 369.960 2200.000 370.560 ;
    END
  END eu1_instruction[21]
  PIN eu1_instruction[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 371.320 2200.000 371.920 ;
    END
  END eu1_instruction[22]
  PIN eu1_instruction[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 372.680 2200.000 373.280 ;
    END
  END eu1_instruction[23]
  PIN eu1_instruction[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 374.040 2200.000 374.640 ;
    END
  END eu1_instruction[24]
  PIN eu1_instruction[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 375.400 2200.000 376.000 ;
    END
  END eu1_instruction[25]
  PIN eu1_instruction[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 376.760 2200.000 377.360 ;
    END
  END eu1_instruction[26]
  PIN eu1_instruction[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 378.120 2200.000 378.720 ;
    END
  END eu1_instruction[27]
  PIN eu1_instruction[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 379.480 2200.000 380.080 ;
    END
  END eu1_instruction[28]
  PIN eu1_instruction[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 380.840 2200.000 381.440 ;
    END
  END eu1_instruction[29]
  PIN eu1_instruction[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 344.120 2200.000 344.720 ;
    END
  END eu1_instruction[2]
  PIN eu1_instruction[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 382.200 2200.000 382.800 ;
    END
  END eu1_instruction[30]
  PIN eu1_instruction[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 383.560 2200.000 384.160 ;
    END
  END eu1_instruction[31]
  PIN eu1_instruction[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 384.920 2200.000 385.520 ;
    END
  END eu1_instruction[32]
  PIN eu1_instruction[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 386.280 2200.000 386.880 ;
    END
  END eu1_instruction[33]
  PIN eu1_instruction[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 387.640 2200.000 388.240 ;
    END
  END eu1_instruction[34]
  PIN eu1_instruction[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 389.000 2200.000 389.600 ;
    END
  END eu1_instruction[35]
  PIN eu1_instruction[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 390.360 2200.000 390.960 ;
    END
  END eu1_instruction[36]
  PIN eu1_instruction[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 391.720 2200.000 392.320 ;
    END
  END eu1_instruction[37]
  PIN eu1_instruction[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 393.080 2200.000 393.680 ;
    END
  END eu1_instruction[38]
  PIN eu1_instruction[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 394.440 2200.000 395.040 ;
    END
  END eu1_instruction[39]
  PIN eu1_instruction[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 345.480 2200.000 346.080 ;
    END
  END eu1_instruction[3]
  PIN eu1_instruction[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 395.800 2200.000 396.400 ;
    END
  END eu1_instruction[40]
  PIN eu1_instruction[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 397.160 2200.000 397.760 ;
    END
  END eu1_instruction[41]
  PIN eu1_instruction[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 346.840 2200.000 347.440 ;
    END
  END eu1_instruction[4]
  PIN eu1_instruction[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 348.200 2200.000 348.800 ;
    END
  END eu1_instruction[5]
  PIN eu1_instruction[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 349.560 2200.000 350.160 ;
    END
  END eu1_instruction[6]
  PIN eu1_instruction[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 350.920 2200.000 351.520 ;
    END
  END eu1_instruction[7]
  PIN eu1_instruction[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 352.280 2200.000 352.880 ;
    END
  END eu1_instruction[8]
  PIN eu1_instruction[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 353.640 2200.000 354.240 ;
    END
  END eu1_instruction[9]
  PIN eu2_busy
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 0.000 349.560 4.000 350.160 ;
    END
  END eu2_busy
  PIN eu2_instruction[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 352.280 4.000 352.880 ;
    END
  END eu2_instruction[0]
  PIN eu2_instruction[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 379.480 4.000 380.080 ;
    END
  END eu2_instruction[10]
  PIN eu2_instruction[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 382.200 4.000 382.800 ;
    END
  END eu2_instruction[11]
  PIN eu2_instruction[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.920 4.000 385.520 ;
    END
  END eu2_instruction[12]
  PIN eu2_instruction[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 387.640 4.000 388.240 ;
    END
  END eu2_instruction[13]
  PIN eu2_instruction[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 390.360 4.000 390.960 ;
    END
  END eu2_instruction[14]
  PIN eu2_instruction[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 393.080 4.000 393.680 ;
    END
  END eu2_instruction[15]
  PIN eu2_instruction[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 395.800 4.000 396.400 ;
    END
  END eu2_instruction[16]
  PIN eu2_instruction[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 398.520 4.000 399.120 ;
    END
  END eu2_instruction[17]
  PIN eu2_instruction[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 401.240 4.000 401.840 ;
    END
  END eu2_instruction[18]
  PIN eu2_instruction[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 403.960 4.000 404.560 ;
    END
  END eu2_instruction[19]
  PIN eu2_instruction[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 355.000 4.000 355.600 ;
    END
  END eu2_instruction[1]
  PIN eu2_instruction[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 406.680 4.000 407.280 ;
    END
  END eu2_instruction[20]
  PIN eu2_instruction[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 409.400 4.000 410.000 ;
    END
  END eu2_instruction[21]
  PIN eu2_instruction[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 412.120 4.000 412.720 ;
    END
  END eu2_instruction[22]
  PIN eu2_instruction[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 414.840 4.000 415.440 ;
    END
  END eu2_instruction[23]
  PIN eu2_instruction[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 417.560 4.000 418.160 ;
    END
  END eu2_instruction[24]
  PIN eu2_instruction[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 420.280 4.000 420.880 ;
    END
  END eu2_instruction[25]
  PIN eu2_instruction[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 423.000 4.000 423.600 ;
    END
  END eu2_instruction[26]
  PIN eu2_instruction[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 425.720 4.000 426.320 ;
    END
  END eu2_instruction[27]
  PIN eu2_instruction[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 428.440 4.000 429.040 ;
    END
  END eu2_instruction[28]
  PIN eu2_instruction[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 431.160 4.000 431.760 ;
    END
  END eu2_instruction[29]
  PIN eu2_instruction[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.720 4.000 358.320 ;
    END
  END eu2_instruction[2]
  PIN eu2_instruction[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 433.880 4.000 434.480 ;
    END
  END eu2_instruction[30]
  PIN eu2_instruction[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 436.600 4.000 437.200 ;
    END
  END eu2_instruction[31]
  PIN eu2_instruction[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 439.320 4.000 439.920 ;
    END
  END eu2_instruction[32]
  PIN eu2_instruction[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 442.040 4.000 442.640 ;
    END
  END eu2_instruction[33]
  PIN eu2_instruction[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 444.760 4.000 445.360 ;
    END
  END eu2_instruction[34]
  PIN eu2_instruction[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 447.480 4.000 448.080 ;
    END
  END eu2_instruction[35]
  PIN eu2_instruction[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 450.200 4.000 450.800 ;
    END
  END eu2_instruction[36]
  PIN eu2_instruction[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 452.920 4.000 453.520 ;
    END
  END eu2_instruction[37]
  PIN eu2_instruction[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 455.640 4.000 456.240 ;
    END
  END eu2_instruction[38]
  PIN eu2_instruction[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 458.360 4.000 458.960 ;
    END
  END eu2_instruction[39]
  PIN eu2_instruction[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 360.440 4.000 361.040 ;
    END
  END eu2_instruction[3]
  PIN eu2_instruction[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 461.080 4.000 461.680 ;
    END
  END eu2_instruction[40]
  PIN eu2_instruction[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 463.800 4.000 464.400 ;
    END
  END eu2_instruction[41]
  PIN eu2_instruction[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.160 4.000 363.760 ;
    END
  END eu2_instruction[4]
  PIN eu2_instruction[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 365.880 4.000 366.480 ;
    END
  END eu2_instruction[5]
  PIN eu2_instruction[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 368.600 4.000 369.200 ;
    END
  END eu2_instruction[6]
  PIN eu2_instruction[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 371.320 4.000 371.920 ;
    END
  END eu2_instruction[7]
  PIN eu2_instruction[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.040 4.000 374.640 ;
    END
  END eu2_instruction[8]
  PIN eu2_instruction[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 376.760 4.000 377.360 ;
    END
  END eu2_instruction[9]
  PIN int_return0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 2162.090 646.000 2162.370 650.000 ;
    END
  END int_return0
  PIN int_return1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 486.920 2200.000 487.520 ;
    END
  END int_return1
  PIN int_return2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 643.320 4.000 643.920 ;
    END
  END int_return2
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 1160.670 0.000 1160.950 4.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.106000 ;
    ANTENNADIFFAREA 2.608200 ;
    PORT
      LAYER met2 ;
        RECT 1248.070 0.000 1248.350 4.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.106000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1256.810 0.000 1257.090 4.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.106000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1265.550 0.000 1265.830 4.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.106000 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met2 ;
        RECT 1274.290 0.000 1274.570 4.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.106000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1283.030 0.000 1283.310 4.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.353500 ;
    ANTENNADIFFAREA 2.173500 ;
    PORT
      LAYER met2 ;
        RECT 1291.770 0.000 1292.050 4.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.353500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1300.510 0.000 1300.790 4.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.848500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1309.250 0.000 1309.530 4.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.727000 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met2 ;
        RECT 1317.990 0.000 1318.270 4.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1326.730 0.000 1327.010 4.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1169.410 0.000 1169.690 4.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1335.470 0.000 1335.750 4.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1344.210 0.000 1344.490 4.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1352.950 0.000 1353.230 4.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1361.690 0.000 1361.970 4.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1370.430 0.000 1370.710 4.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1379.170 0.000 1379.450 4.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER met2 ;
        RECT 1387.910 0.000 1388.190 4.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1396.650 0.000 1396.930 4.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1405.390 0.000 1405.670 4.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 1414.130 0.000 1414.410 4.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 1178.150 0.000 1178.430 4.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 1422.870 0.000 1423.150 4.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.621000 ;
    PORT
      LAYER met2 ;
        RECT 1431.610 0.000 1431.890 4.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 1440.350 0.000 1440.630 4.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 1449.090 0.000 1449.370 4.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 1457.830 0.000 1458.110 4.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 1466.570 0.000 1466.850 4.000 ;
    END
  END io_in[35]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.106000 ;
    PORT
      LAYER met2 ;
        RECT 1186.890 0.000 1187.170 4.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.980000 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met2 ;
        RECT 1195.630 0.000 1195.910 4.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.227500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1204.370 0.000 1204.650 4.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.980000 ;
    ANTENNADIFFAREA 2.173500 ;
    PORT
      LAYER met2 ;
        RECT 1213.110 0.000 1213.390 4.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.227500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1221.850 0.000 1222.130 4.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.227500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1230.590 0.000 1230.870 4.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.227500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1239.330 0.000 1239.610 4.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.484000 ;
    PORT
      LAYER met2 ;
        RECT 1475.310 0.000 1475.590 4.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1562.710 0.000 1562.990 4.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1571.450 0.000 1571.730 4.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1580.190 0.000 1580.470 4.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1588.930 0.000 1589.210 4.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1597.670 0.000 1597.950 4.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1606.410 0.000 1606.690 4.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1615.150 0.000 1615.430 4.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1623.890 0.000 1624.170 4.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 13.860000 ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1632.630 0.000 1632.910 4.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1641.370 0.000 1641.650 4.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1484.050 0.000 1484.330 4.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1650.110 0.000 1650.390 4.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1658.850 0.000 1659.130 4.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1667.590 0.000 1667.870 4.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1676.330 0.000 1676.610 4.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1685.070 0.000 1685.350 4.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1693.810 0.000 1694.090 4.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1702.550 0.000 1702.830 4.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1711.290 0.000 1711.570 4.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1720.030 0.000 1720.310 4.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1728.770 0.000 1729.050 4.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.484000 ;
    PORT
      LAYER met2 ;
        RECT 1492.790 0.000 1493.070 4.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1737.510 0.000 1737.790 4.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1746.250 0.000 1746.530 4.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1754.990 0.000 1755.270 4.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1763.730 0.000 1764.010 4.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1772.470 0.000 1772.750 4.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1781.210 0.000 1781.490 4.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1501.530 0.000 1501.810 4.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1510.270 0.000 1510.550 4.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1519.010 0.000 1519.290 4.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1527.750 0.000 1528.030 4.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1536.490 0.000 1536.770 4.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1545.230 0.000 1545.510 4.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1553.970 0.000 1554.250 4.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1789.950 0.000 1790.230 4.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1877.350 0.000 1877.630 4.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1886.090 0.000 1886.370 4.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1894.830 0.000 1895.110 4.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1903.570 0.000 1903.850 4.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1912.310 0.000 1912.590 4.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1921.050 0.000 1921.330 4.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1929.790 0.000 1930.070 4.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1938.530 0.000 1938.810 4.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.484000 ;
    PORT
      LAYER met2 ;
        RECT 1947.270 0.000 1947.550 4.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1956.010 0.000 1956.290 4.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1798.690 0.000 1798.970 4.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1964.750 0.000 1965.030 4.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1973.490 0.000 1973.770 4.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1982.230 0.000 1982.510 4.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1990.970 0.000 1991.250 4.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.462000 ;
    PORT
      LAYER met2 ;
        RECT 1999.710 0.000 1999.990 4.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 2008.450 0.000 2008.730 4.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2017.190 0.000 2017.470 4.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 2025.930 0.000 2026.210 4.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 2034.670 0.000 2034.950 4.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2043.410 0.000 2043.690 4.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1807.430 0.000 1807.710 4.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 2052.150 0.000 2052.430 4.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 2060.890 0.000 2061.170 4.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 3.499200 ;
    PORT
      LAYER met2 ;
        RECT 2069.630 0.000 2069.910 4.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 2078.370 0.000 2078.650 4.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 2087.110 0.000 2087.390 4.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 2095.850 0.000 2096.130 4.000 ;
    END
  END io_out[35]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1816.170 0.000 1816.450 4.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1824.910 0.000 1825.190 4.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1833.650 0.000 1833.930 4.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1842.390 0.000 1842.670 4.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1851.130 0.000 1851.410 4.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1859.870 0.000 1860.150 4.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1868.610 0.000 1868.890 4.000 ;
    END
  END io_out[9]
  PIN is_load0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1418.270 646.000 1418.550 650.000 ;
    END
  END is_load0
  PIN is_load1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.621000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 287.000 2200.000 287.600 ;
    END
  END is_load1
  PIN is_load2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.621000 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 0.000 243.480 4.000 244.080 ;
    END
  END is_load2
  PIN is_store0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.621000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1423.330 646.000 1423.610 650.000 ;
    END
  END is_store0
  PIN is_store1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 288.360 2200.000 288.960 ;
    END
  END is_store1
  PIN is_store2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 246.200 4.000 246.800 ;
    END
  END is_store2
  PIN loadstore_address0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1256.350 646.000 1256.630 650.000 ;
    END
  END loadstore_address0[0]
  PIN loadstore_address0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1306.950 646.000 1307.230 650.000 ;
    END
  END loadstore_address0[10]
  PIN loadstore_address0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1312.010 646.000 1312.290 650.000 ;
    END
  END loadstore_address0[11]
  PIN loadstore_address0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1317.070 646.000 1317.350 650.000 ;
    END
  END loadstore_address0[12]
  PIN loadstore_address0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1322.130 646.000 1322.410 650.000 ;
    END
  END loadstore_address0[13]
  PIN loadstore_address0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1327.190 646.000 1327.470 650.000 ;
    END
  END loadstore_address0[14]
  PIN loadstore_address0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1332.250 646.000 1332.530 650.000 ;
    END
  END loadstore_address0[15]
  PIN loadstore_address0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1337.310 646.000 1337.590 650.000 ;
    END
  END loadstore_address0[16]
  PIN loadstore_address0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1342.370 646.000 1342.650 650.000 ;
    END
  END loadstore_address0[17]
  PIN loadstore_address0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1347.430 646.000 1347.710 650.000 ;
    END
  END loadstore_address0[18]
  PIN loadstore_address0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1352.490 646.000 1352.770 650.000 ;
    END
  END loadstore_address0[19]
  PIN loadstore_address0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1261.410 646.000 1261.690 650.000 ;
    END
  END loadstore_address0[1]
  PIN loadstore_address0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1357.550 646.000 1357.830 650.000 ;
    END
  END loadstore_address0[20]
  PIN loadstore_address0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1362.610 646.000 1362.890 650.000 ;
    END
  END loadstore_address0[21]
  PIN loadstore_address0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1367.670 646.000 1367.950 650.000 ;
    END
  END loadstore_address0[22]
  PIN loadstore_address0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1372.730 646.000 1373.010 650.000 ;
    END
  END loadstore_address0[23]
  PIN loadstore_address0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1377.790 646.000 1378.070 650.000 ;
    END
  END loadstore_address0[24]
  PIN loadstore_address0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1382.850 646.000 1383.130 650.000 ;
    END
  END loadstore_address0[25]
  PIN loadstore_address0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1387.910 646.000 1388.190 650.000 ;
    END
  END loadstore_address0[26]
  PIN loadstore_address0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1392.970 646.000 1393.250 650.000 ;
    END
  END loadstore_address0[27]
  PIN loadstore_address0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1398.030 646.000 1398.310 650.000 ;
    END
  END loadstore_address0[28]
  PIN loadstore_address0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1403.090 646.000 1403.370 650.000 ;
    END
  END loadstore_address0[29]
  PIN loadstore_address0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1266.470 646.000 1266.750 650.000 ;
    END
  END loadstore_address0[2]
  PIN loadstore_address0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1408.150 646.000 1408.430 650.000 ;
    END
  END loadstore_address0[30]
  PIN loadstore_address0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1413.210 646.000 1413.490 650.000 ;
    END
  END loadstore_address0[31]
  PIN loadstore_address0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1271.530 646.000 1271.810 650.000 ;
    END
  END loadstore_address0[3]
  PIN loadstore_address0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1276.590 646.000 1276.870 650.000 ;
    END
  END loadstore_address0[4]
  PIN loadstore_address0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1281.650 646.000 1281.930 650.000 ;
    END
  END loadstore_address0[5]
  PIN loadstore_address0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1286.710 646.000 1286.990 650.000 ;
    END
  END loadstore_address0[6]
  PIN loadstore_address0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1291.770 646.000 1292.050 650.000 ;
    END
  END loadstore_address0[7]
  PIN loadstore_address0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1296.830 646.000 1297.110 650.000 ;
    END
  END loadstore_address0[8]
  PIN loadstore_address0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1301.890 646.000 1302.170 650.000 ;
    END
  END loadstore_address0[9]
  PIN loadstore_address1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 243.480 2200.000 244.080 ;
    END
  END loadstore_address1[0]
  PIN loadstore_address1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 257.080 2200.000 257.680 ;
    END
  END loadstore_address1[10]
  PIN loadstore_address1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 258.440 2200.000 259.040 ;
    END
  END loadstore_address1[11]
  PIN loadstore_address1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 259.800 2200.000 260.400 ;
    END
  END loadstore_address1[12]
  PIN loadstore_address1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 261.160 2200.000 261.760 ;
    END
  END loadstore_address1[13]
  PIN loadstore_address1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 7.389900 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 262.520 2200.000 263.120 ;
    END
  END loadstore_address1[14]
  PIN loadstore_address1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 263.880 2200.000 264.480 ;
    END
  END loadstore_address1[15]
  PIN loadstore_address1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 265.240 2200.000 265.840 ;
    END
  END loadstore_address1[16]
  PIN loadstore_address1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 266.600 2200.000 267.200 ;
    END
  END loadstore_address1[17]
  PIN loadstore_address1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 267.960 2200.000 268.560 ;
    END
  END loadstore_address1[18]
  PIN loadstore_address1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 269.320 2200.000 269.920 ;
    END
  END loadstore_address1[19]
  PIN loadstore_address1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 244.840 2200.000 245.440 ;
    END
  END loadstore_address1[1]
  PIN loadstore_address1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 3.912300 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 270.680 2200.000 271.280 ;
    END
  END loadstore_address1[20]
  PIN loadstore_address1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 5.216400 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 272.040 2200.000 272.640 ;
    END
  END loadstore_address1[21]
  PIN loadstore_address1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 7.389900 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 273.400 2200.000 274.000 ;
    END
  END loadstore_address1[22]
  PIN loadstore_address1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 2.173500 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 274.760 2200.000 275.360 ;
    END
  END loadstore_address1[23]
  PIN loadstore_address1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 276.120 2200.000 276.720 ;
    END
  END loadstore_address1[24]
  PIN loadstore_address1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 277.480 2200.000 278.080 ;
    END
  END loadstore_address1[25]
  PIN loadstore_address1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 278.840 2200.000 279.440 ;
    END
  END loadstore_address1[26]
  PIN loadstore_address1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 8.694000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 280.200 2200.000 280.800 ;
    END
  END loadstore_address1[27]
  PIN loadstore_address1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 281.560 2200.000 282.160 ;
    END
  END loadstore_address1[28]
  PIN loadstore_address1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 282.920 2200.000 283.520 ;
    END
  END loadstore_address1[29]
  PIN loadstore_address1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 2.173500 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 246.200 2200.000 246.800 ;
    END
  END loadstore_address1[2]
  PIN loadstore_address1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 284.280 2200.000 284.880 ;
    END
  END loadstore_address1[30]
  PIN loadstore_address1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 285.640 2200.000 286.240 ;
    END
  END loadstore_address1[31]
  PIN loadstore_address1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 5.216400 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 247.560 2200.000 248.160 ;
    END
  END loadstore_address1[3]
  PIN loadstore_address1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 248.920 2200.000 249.520 ;
    END
  END loadstore_address1[4]
  PIN loadstore_address1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 250.280 2200.000 250.880 ;
    END
  END loadstore_address1[5]
  PIN loadstore_address1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 251.640 2200.000 252.240 ;
    END
  END loadstore_address1[6]
  PIN loadstore_address1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 5.216400 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 253.000 2200.000 253.600 ;
    END
  END loadstore_address1[7]
  PIN loadstore_address1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 8.694000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 254.360 2200.000 254.960 ;
    END
  END loadstore_address1[8]
  PIN loadstore_address1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 255.720 2200.000 256.320 ;
    END
  END loadstore_address1[9]
  PIN loadstore_address2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END loadstore_address2[0]
  PIN loadstore_address2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END loadstore_address2[10]
  PIN loadstore_address2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 186.360 4.000 186.960 ;
    END
  END loadstore_address2[11]
  PIN loadstore_address2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 9.998099 ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.080 4.000 189.680 ;
    END
  END loadstore_address2[12]
  PIN loadstore_address2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.800 4.000 192.400 ;
    END
  END loadstore_address2[13]
  PIN loadstore_address2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 14.345099 ;
    PORT
      LAYER met3 ;
        RECT 0.000 194.520 4.000 195.120 ;
    END
  END loadstore_address2[14]
  PIN loadstore_address2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.240 4.000 197.840 ;
    END
  END loadstore_address2[15]
  PIN loadstore_address2[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 20.865599 ;
    PORT
      LAYER met3 ;
        RECT 0.000 199.960 4.000 200.560 ;
    END
  END loadstore_address2[16]
  PIN loadstore_address2[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 15.214499 ;
    PORT
      LAYER met3 ;
        RECT 0.000 202.680 4.000 203.280 ;
    END
  END loadstore_address2[17]
  PIN loadstore_address2[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 22.604399 ;
    PORT
      LAYER met3 ;
        RECT 0.000 205.400 4.000 206.000 ;
    END
  END loadstore_address2[18]
  PIN loadstore_address2[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 9.998099 ;
    PORT
      LAYER met3 ;
        RECT 0.000 208.120 4.000 208.720 ;
    END
  END loadstore_address2[19]
  PIN loadstore_address2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 9.998099 ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.160 4.000 159.760 ;
    END
  END loadstore_address2[1]
  PIN loadstore_address2[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.840 4.000 211.440 ;
    END
  END loadstore_address2[20]
  PIN loadstore_address2[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 213.560 4.000 214.160 ;
    END
  END loadstore_address2[21]
  PIN loadstore_address2[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 19.126799 ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.280 4.000 216.880 ;
    END
  END loadstore_address2[22]
  PIN loadstore_address2[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 9.998099 ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.000 4.000 219.600 ;
    END
  END loadstore_address2[23]
  PIN loadstore_address2[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.720 4.000 222.320 ;
    END
  END loadstore_address2[24]
  PIN loadstore_address2[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.440 4.000 225.040 ;
    END
  END loadstore_address2[25]
  PIN loadstore_address2[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.160 4.000 227.760 ;
    END
  END loadstore_address2[26]
  PIN loadstore_address2[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.880 4.000 230.480 ;
    END
  END loadstore_address2[27]
  PIN loadstore_address2[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 232.600 4.000 233.200 ;
    END
  END loadstore_address2[28]
  PIN loadstore_address2[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 16.518600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 235.320 4.000 235.920 ;
    END
  END loadstore_address2[29]
  PIN loadstore_address2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.880 4.000 162.480 ;
    END
  END loadstore_address2[2]
  PIN loadstore_address2[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 6.085800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.040 4.000 238.640 ;
    END
  END loadstore_address2[30]
  PIN loadstore_address2[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 19.561499 ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.760 4.000 241.360 ;
    END
  END loadstore_address2[31]
  PIN loadstore_address2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 164.600 4.000 165.200 ;
    END
  END loadstore_address2[3]
  PIN loadstore_address2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 167.320 4.000 167.920 ;
    END
  END loadstore_address2[4]
  PIN loadstore_address2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END loadstore_address2[5]
  PIN loadstore_address2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.760 4.000 173.360 ;
    END
  END loadstore_address2[6]
  PIN loadstore_address2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 175.480 4.000 176.080 ;
    END
  END loadstore_address2[7]
  PIN loadstore_address2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.200 4.000 178.800 ;
    END
  END loadstore_address2[8]
  PIN loadstore_address2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.920 4.000 181.520 ;
    END
  END loadstore_address2[9]
  PIN loadstore_dest0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 3.477600 ;
    PORT
      LAYER met2 ;
        RECT 1443.570 646.000 1443.850 650.000 ;
    END
  END loadstore_dest0[0]
  PIN loadstore_dest0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met2 ;
        RECT 1448.630 646.000 1448.910 650.000 ;
    END
  END loadstore_dest0[1]
  PIN loadstore_dest0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met2 ;
        RECT 1453.690 646.000 1453.970 650.000 ;
    END
  END loadstore_dest0[2]
  PIN loadstore_dest0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met2 ;
        RECT 1458.750 646.000 1459.030 650.000 ;
    END
  END loadstore_dest0[3]
  PIN loadstore_dest0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met2 ;
        RECT 1463.810 646.000 1464.090 650.000 ;
    END
  END loadstore_dest0[4]
  PIN loadstore_dest1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.237500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 293.800 2200.000 294.400 ;
    END
  END loadstore_dest1[0]
  PIN loadstore_dest1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.237500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 295.160 2200.000 295.760 ;
    END
  END loadstore_dest1[1]
  PIN loadstore_dest1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.485000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 296.520 2200.000 297.120 ;
    END
  END loadstore_dest1[2]
  PIN loadstore_dest1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.485000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 297.880 2200.000 298.480 ;
    END
  END loadstore_dest1[3]
  PIN loadstore_dest1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.485000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 299.240 2200.000 299.840 ;
    END
  END loadstore_dest1[4]
  PIN loadstore_dest2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.237500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 257.080 4.000 257.680 ;
    END
  END loadstore_dest2[0]
  PIN loadstore_dest2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.237500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.800 4.000 260.400 ;
    END
  END loadstore_dest2[1]
  PIN loadstore_dest2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.485000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 262.520 4.000 263.120 ;
    END
  END loadstore_dest2[2]
  PIN loadstore_dest2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.485000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.240 4.000 265.840 ;
    END
  END loadstore_dest2[3]
  PIN loadstore_dest2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.485000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 267.960 4.000 268.560 ;
    END
  END loadstore_dest2[4]
  PIN loadstore_size0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1433.450 646.000 1433.730 650.000 ;
    END
  END loadstore_size0[0]
  PIN loadstore_size0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1438.510 646.000 1438.790 650.000 ;
    END
  END loadstore_size0[1]
  PIN loadstore_size1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 291.080 2200.000 291.680 ;
    END
  END loadstore_size1[0]
  PIN loadstore_size1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 292.440 2200.000 293.040 ;
    END
  END loadstore_size1[1]
  PIN loadstore_size2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.640 4.000 252.240 ;
    END
  END loadstore_size2[0]
  PIN loadstore_size2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 15.214499 ;
    PORT
      LAYER met3 ;
        RECT 0.000 254.360 4.000 254.960 ;
    END
  END loadstore_size2[1]
  PIN new_PC0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1473.930 646.000 1474.210 650.000 ;
    END
  END new_PC0[0]
  PIN new_PC0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1524.530 646.000 1524.810 650.000 ;
    END
  END new_PC0[10]
  PIN new_PC0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1529.590 646.000 1529.870 650.000 ;
    END
  END new_PC0[11]
  PIN new_PC0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 3.042900 ;
    PORT
      LAYER met2 ;
        RECT 1534.650 646.000 1534.930 650.000 ;
    END
  END new_PC0[12]
  PIN new_PC0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 2.608200 ;
    PORT
      LAYER met2 ;
        RECT 1539.710 646.000 1539.990 650.000 ;
    END
  END new_PC0[13]
  PIN new_PC0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 3.042900 ;
    PORT
      LAYER met2 ;
        RECT 1544.770 646.000 1545.050 650.000 ;
    END
  END new_PC0[14]
  PIN new_PC0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 2.173500 ;
    PORT
      LAYER met2 ;
        RECT 1549.830 646.000 1550.110 650.000 ;
    END
  END new_PC0[15]
  PIN new_PC0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 5.216400 ;
    PORT
      LAYER met2 ;
        RECT 1554.890 646.000 1555.170 650.000 ;
    END
  END new_PC0[16]
  PIN new_PC0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1559.950 646.000 1560.230 650.000 ;
    END
  END new_PC0[17]
  PIN new_PC0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 5.216400 ;
    PORT
      LAYER met2 ;
        RECT 1565.010 646.000 1565.290 650.000 ;
    END
  END new_PC0[18]
  PIN new_PC0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 3.042900 ;
    PORT
      LAYER met2 ;
        RECT 1570.070 646.000 1570.350 650.000 ;
    END
  END new_PC0[19]
  PIN new_PC0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1478.990 646.000 1479.270 650.000 ;
    END
  END new_PC0[1]
  PIN new_PC0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 2.608200 ;
    PORT
      LAYER met2 ;
        RECT 1575.130 646.000 1575.410 650.000 ;
    END
  END new_PC0[20]
  PIN new_PC0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1580.190 646.000 1580.470 650.000 ;
    END
  END new_PC0[21]
  PIN new_PC0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1585.250 646.000 1585.530 650.000 ;
    END
  END new_PC0[22]
  PIN new_PC0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 4.347000 ;
    PORT
      LAYER met2 ;
        RECT 1590.310 646.000 1590.590 650.000 ;
    END
  END new_PC0[23]
  PIN new_PC0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1595.370 646.000 1595.650 650.000 ;
    END
  END new_PC0[24]
  PIN new_PC0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1600.430 646.000 1600.710 650.000 ;
    END
  END new_PC0[25]
  PIN new_PC0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met2 ;
        RECT 1605.490 646.000 1605.770 650.000 ;
    END
  END new_PC0[26]
  PIN new_PC0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 1610.550 646.000 1610.830 650.000 ;
    END
  END new_PC0[27]
  PIN new_PC0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1484.050 646.000 1484.330 650.000 ;
    END
  END new_PC0[2]
  PIN new_PC0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met2 ;
        RECT 1489.110 646.000 1489.390 650.000 ;
    END
  END new_PC0[3]
  PIN new_PC0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 5.651100 ;
    PORT
      LAYER met2 ;
        RECT 1494.170 646.000 1494.450 650.000 ;
    END
  END new_PC0[4]
  PIN new_PC0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 2.608200 ;
    PORT
      LAYER met2 ;
        RECT 1499.230 646.000 1499.510 650.000 ;
    END
  END new_PC0[5]
  PIN new_PC0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 5.216400 ;
    PORT
      LAYER met2 ;
        RECT 1504.290 646.000 1504.570 650.000 ;
    END
  END new_PC0[6]
  PIN new_PC0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1509.350 646.000 1509.630 650.000 ;
    END
  END new_PC0[7]
  PIN new_PC0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 4.347000 ;
    PORT
      LAYER met2 ;
        RECT 1514.410 646.000 1514.690 650.000 ;
    END
  END new_PC0[8]
  PIN new_PC0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 5.216400 ;
    PORT
      LAYER met2 ;
        RECT 1519.470 646.000 1519.750 650.000 ;
    END
  END new_PC0[9]
  PIN new_PC1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 3.042900 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 301.960 2200.000 302.560 ;
    END
  END new_PC1[0]
  PIN new_PC1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 5.216400 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 315.560 2200.000 316.160 ;
    END
  END new_PC1[10]
  PIN new_PC1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.347000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 316.920 2200.000 317.520 ;
    END
  END new_PC1[11]
  PIN new_PC1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 318.280 2200.000 318.880 ;
    END
  END new_PC1[12]
  PIN new_PC1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 5.651100 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 319.640 2200.000 320.240 ;
    END
  END new_PC1[13]
  PIN new_PC1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 321.000 2200.000 321.600 ;
    END
  END new_PC1[14]
  PIN new_PC1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 7.389900 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 322.360 2200.000 322.960 ;
    END
  END new_PC1[15]
  PIN new_PC1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 323.720 2200.000 324.320 ;
    END
  END new_PC1[16]
  PIN new_PC1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 325.080 2200.000 325.680 ;
    END
  END new_PC1[17]
  PIN new_PC1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 326.440 2200.000 327.040 ;
    END
  END new_PC1[18]
  PIN new_PC1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 327.800 2200.000 328.400 ;
    END
  END new_PC1[19]
  PIN new_PC1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 303.320 2200.000 303.920 ;
    END
  END new_PC1[1]
  PIN new_PC1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 3.042900 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 329.160 2200.000 329.760 ;
    END
  END new_PC1[20]
  PIN new_PC1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 330.520 2200.000 331.120 ;
    END
  END new_PC1[21]
  PIN new_PC1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 331.880 2200.000 332.480 ;
    END
  END new_PC1[22]
  PIN new_PC1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 7.389900 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 333.240 2200.000 333.840 ;
    END
  END new_PC1[23]
  PIN new_PC1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 2.173500 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 334.600 2200.000 335.200 ;
    END
  END new_PC1[24]
  PIN new_PC1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 335.960 2200.000 336.560 ;
    END
  END new_PC1[25]
  PIN new_PC1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 337.320 2200.000 337.920 ;
    END
  END new_PC1[26]
  PIN new_PC1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.980000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 338.680 2200.000 339.280 ;
    END
  END new_PC1[27]
  PIN new_PC1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 9.998099 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 304.680 2200.000 305.280 ;
    END
  END new_PC1[2]
  PIN new_PC1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 306.040 2200.000 306.640 ;
    END
  END new_PC1[3]
  PIN new_PC1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 3.042900 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 307.400 2200.000 308.000 ;
    END
  END new_PC1[4]
  PIN new_PC1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 308.760 2200.000 309.360 ;
    END
  END new_PC1[5]
  PIN new_PC1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 15.214499 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 310.120 2200.000 310.720 ;
    END
  END new_PC1[6]
  PIN new_PC1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 311.480 2200.000 312.080 ;
    END
  END new_PC1[7]
  PIN new_PC1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 3.042900 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 312.840 2200.000 313.440 ;
    END
  END new_PC1[8]
  PIN new_PC1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 5.216400 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 314.200 2200.000 314.800 ;
    END
  END new_PC1[9]
  PIN new_PC2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 273.400 4.000 274.000 ;
    END
  END new_PC2[0]
  PIN new_PC2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 300.600 4.000 301.200 ;
    END
  END new_PC2[10]
  PIN new_PC2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 303.320 4.000 303.920 ;
    END
  END new_PC2[11]
  PIN new_PC2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.040 4.000 306.640 ;
    END
  END new_PC2[12]
  PIN new_PC2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 308.760 4.000 309.360 ;
    END
  END new_PC2[13]
  PIN new_PC2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 311.480 4.000 312.080 ;
    END
  END new_PC2[14]
  PIN new_PC2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 314.200 4.000 314.800 ;
    END
  END new_PC2[15]
  PIN new_PC2[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.920 4.000 317.520 ;
    END
  END new_PC2[16]
  PIN new_PC2[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 319.640 4.000 320.240 ;
    END
  END new_PC2[17]
  PIN new_PC2[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 322.360 4.000 322.960 ;
    END
  END new_PC2[18]
  PIN new_PC2[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 9.998099 ;
    PORT
      LAYER met3 ;
        RECT 0.000 325.080 4.000 325.680 ;
    END
  END new_PC2[19]
  PIN new_PC2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 276.120 4.000 276.720 ;
    END
  END new_PC2[1]
  PIN new_PC2[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 327.800 4.000 328.400 ;
    END
  END new_PC2[20]
  PIN new_PC2[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 330.520 4.000 331.120 ;
    END
  END new_PC2[21]
  PIN new_PC2[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.240 4.000 333.840 ;
    END
  END new_PC2[22]
  PIN new_PC2[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 335.960 4.000 336.560 ;
    END
  END new_PC2[23]
  PIN new_PC2[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 338.680 4.000 339.280 ;
    END
  END new_PC2[24]
  PIN new_PC2[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 5.651100 ;
    PORT
      LAYER met3 ;
        RECT 0.000 341.400 4.000 342.000 ;
    END
  END new_PC2[25]
  PIN new_PC2[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.347000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 344.120 4.000 344.720 ;
    END
  END new_PC2[26]
  PIN new_PC2[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.840 4.000 347.440 ;
    END
  END new_PC2[27]
  PIN new_PC2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.840 4.000 279.440 ;
    END
  END new_PC2[2]
  PIN new_PC2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 281.560 4.000 282.160 ;
    END
  END new_PC2[3]
  PIN new_PC2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 284.280 4.000 284.880 ;
    END
  END new_PC2[4]
  PIN new_PC2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 287.000 4.000 287.600 ;
    END
  END new_PC2[5]
  PIN new_PC2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.720 4.000 290.320 ;
    END
  END new_PC2[6]
  PIN new_PC2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.440 4.000 293.040 ;
    END
  END new_PC2[7]
  PIN new_PC2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.160 4.000 295.760 ;
    END
  END new_PC2[8]
  PIN new_PC2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 297.880 4.000 298.480 ;
    END
  END new_PC2[9]
  PIN pred_idx0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.696000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1220.930 646.000 1221.210 650.000 ;
    END
  END pred_idx0[0]
  PIN pred_idx0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.696000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1225.990 646.000 1226.270 650.000 ;
    END
  END pred_idx0[1]
  PIN pred_idx0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1231.050 646.000 1231.330 650.000 ;
    END
  END pred_idx0[2]
  PIN pred_idx1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.630000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 233.960 2200.000 234.560 ;
    END
  END pred_idx1[0]
  PIN pred_idx1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.630000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 235.320 2200.000 235.920 ;
    END
  END pred_idx1[1]
  PIN pred_idx1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 236.680 2200.000 237.280 ;
    END
  END pred_idx1[2]
  PIN pred_idx2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.630000 ;
    ANTENNADIFFAREA 2.608200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.400 4.000 138.000 ;
    END
  END pred_idx2[0]
  PIN pred_idx2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.630000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.120 4.000 140.720 ;
    END
  END pred_idx2[1]
  PIN pred_idx2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END pred_idx2[2]
  PIN pred_val0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.962500 ;
    PORT
      LAYER met2 ;
        RECT 2157.030 646.000 2157.310 650.000 ;
    END
  END pred_val0
  PIN pred_val1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.962500 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 485.560 2200.000 486.160 ;
    END
  END pred_val1
  PIN pred_val2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.962500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 640.600 4.000 641.200 ;
    END
  END pred_val2
  PIN reg1_idx0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.574500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 972.990 646.000 973.270 650.000 ;
    END
  END reg1_idx0[0]
  PIN reg1_idx0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 978.050 646.000 978.330 650.000 ;
    END
  END reg1_idx0[1]
  PIN reg1_idx0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.970000 ;
    PORT
      LAYER met2 ;
        RECT 983.110 646.000 983.390 650.000 ;
    END
  END reg1_idx0[2]
  PIN reg1_idx0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.383000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 988.170 646.000 988.450 650.000 ;
    END
  END reg1_idx0[3]
  PIN reg1_idx0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.293000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 993.230 646.000 993.510 650.000 ;
    END
  END reg1_idx0[4]
  PIN reg1_idx1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.406000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 167.320 2200.000 167.920 ;
    END
  END reg1_idx1[0]
  PIN reg1_idx1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.574500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 168.680 2200.000 169.280 ;
    END
  END reg1_idx1[1]
  PIN reg1_idx1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.722500 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 170.040 2200.000 170.640 ;
    END
  END reg1_idx1[2]
  PIN reg1_idx1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.383000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 171.400 2200.000 172.000 ;
    END
  END reg1_idx1[3]
  PIN reg1_idx1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.293000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 172.760 2200.000 173.360 ;
    END
  END reg1_idx1[4]
  PIN reg1_idx2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.842000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.120 4.000 4.720 ;
    END
  END reg1_idx2[0]
  PIN reg1_idx2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.475000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END reg1_idx2[1]
  PIN reg1_idx2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 9.560 4.000 10.160 ;
    END
  END reg1_idx2[2]
  PIN reg1_idx2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.383000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 4.000 12.880 ;
    END
  END reg1_idx2[3]
  PIN reg1_idx2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.293000 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.000 4.000 15.600 ;
    END
  END reg1_idx2[4]
  PIN reg1_val0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1833.190 646.000 1833.470 650.000 ;
    END
  END reg1_val0[0]
  PIN reg1_val0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1883.790 646.000 1884.070 650.000 ;
    END
  END reg1_val0[10]
  PIN reg1_val0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1888.850 646.000 1889.130 650.000 ;
    END
  END reg1_val0[11]
  PIN reg1_val0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1893.910 646.000 1894.190 650.000 ;
    END
  END reg1_val0[12]
  PIN reg1_val0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1898.970 646.000 1899.250 650.000 ;
    END
  END reg1_val0[13]
  PIN reg1_val0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1904.030 646.000 1904.310 650.000 ;
    END
  END reg1_val0[14]
  PIN reg1_val0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1909.090 646.000 1909.370 650.000 ;
    END
  END reg1_val0[15]
  PIN reg1_val0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1914.150 646.000 1914.430 650.000 ;
    END
  END reg1_val0[16]
  PIN reg1_val0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1919.210 646.000 1919.490 650.000 ;
    END
  END reg1_val0[17]
  PIN reg1_val0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1924.270 646.000 1924.550 650.000 ;
    END
  END reg1_val0[18]
  PIN reg1_val0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1929.330 646.000 1929.610 650.000 ;
    END
  END reg1_val0[19]
  PIN reg1_val0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1838.250 646.000 1838.530 650.000 ;
    END
  END reg1_val0[1]
  PIN reg1_val0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1934.390 646.000 1934.670 650.000 ;
    END
  END reg1_val0[20]
  PIN reg1_val0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1939.450 646.000 1939.730 650.000 ;
    END
  END reg1_val0[21]
  PIN reg1_val0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1944.510 646.000 1944.790 650.000 ;
    END
  END reg1_val0[22]
  PIN reg1_val0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1949.570 646.000 1949.850 650.000 ;
    END
  END reg1_val0[23]
  PIN reg1_val0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1954.630 646.000 1954.910 650.000 ;
    END
  END reg1_val0[24]
  PIN reg1_val0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1959.690 646.000 1959.970 650.000 ;
    END
  END reg1_val0[25]
  PIN reg1_val0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1964.750 646.000 1965.030 650.000 ;
    END
  END reg1_val0[26]
  PIN reg1_val0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1969.810 646.000 1970.090 650.000 ;
    END
  END reg1_val0[27]
  PIN reg1_val0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1974.870 646.000 1975.150 650.000 ;
    END
  END reg1_val0[28]
  PIN reg1_val0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1979.930 646.000 1980.210 650.000 ;
    END
  END reg1_val0[29]
  PIN reg1_val0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1843.310 646.000 1843.590 650.000 ;
    END
  END reg1_val0[2]
  PIN reg1_val0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1984.990 646.000 1985.270 650.000 ;
    END
  END reg1_val0[30]
  PIN reg1_val0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1990.050 646.000 1990.330 650.000 ;
    END
  END reg1_val0[31]
  PIN reg1_val0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1848.370 646.000 1848.650 650.000 ;
    END
  END reg1_val0[3]
  PIN reg1_val0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1853.430 646.000 1853.710 650.000 ;
    END
  END reg1_val0[4]
  PIN reg1_val0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1858.490 646.000 1858.770 650.000 ;
    END
  END reg1_val0[5]
  PIN reg1_val0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1863.550 646.000 1863.830 650.000 ;
    END
  END reg1_val0[6]
  PIN reg1_val0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1868.610 646.000 1868.890 650.000 ;
    END
  END reg1_val0[7]
  PIN reg1_val0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1873.670 646.000 1873.950 650.000 ;
    END
  END reg1_val0[8]
  PIN reg1_val0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1878.730 646.000 1879.010 650.000 ;
    END
  END reg1_val0[9]
  PIN reg1_val1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 398.520 2200.000 399.120 ;
    END
  END reg1_val1[0]
  PIN reg1_val1[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 412.120 2200.000 412.720 ;
    END
  END reg1_val1[10]
  PIN reg1_val1[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 413.480 2200.000 414.080 ;
    END
  END reg1_val1[11]
  PIN reg1_val1[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 414.840 2200.000 415.440 ;
    END
  END reg1_val1[12]
  PIN reg1_val1[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 416.200 2200.000 416.800 ;
    END
  END reg1_val1[13]
  PIN reg1_val1[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 417.560 2200.000 418.160 ;
    END
  END reg1_val1[14]
  PIN reg1_val1[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 418.920 2200.000 419.520 ;
    END
  END reg1_val1[15]
  PIN reg1_val1[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 420.280 2200.000 420.880 ;
    END
  END reg1_val1[16]
  PIN reg1_val1[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 421.640 2200.000 422.240 ;
    END
  END reg1_val1[17]
  PIN reg1_val1[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 423.000 2200.000 423.600 ;
    END
  END reg1_val1[18]
  PIN reg1_val1[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 424.360 2200.000 424.960 ;
    END
  END reg1_val1[19]
  PIN reg1_val1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 399.880 2200.000 400.480 ;
    END
  END reg1_val1[1]
  PIN reg1_val1[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 425.720 2200.000 426.320 ;
    END
  END reg1_val1[20]
  PIN reg1_val1[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 427.080 2200.000 427.680 ;
    END
  END reg1_val1[21]
  PIN reg1_val1[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 428.440 2200.000 429.040 ;
    END
  END reg1_val1[22]
  PIN reg1_val1[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 429.800 2200.000 430.400 ;
    END
  END reg1_val1[23]
  PIN reg1_val1[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 431.160 2200.000 431.760 ;
    END
  END reg1_val1[24]
  PIN reg1_val1[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 432.520 2200.000 433.120 ;
    END
  END reg1_val1[25]
  PIN reg1_val1[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 433.880 2200.000 434.480 ;
    END
  END reg1_val1[26]
  PIN reg1_val1[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 435.240 2200.000 435.840 ;
    END
  END reg1_val1[27]
  PIN reg1_val1[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 436.600 2200.000 437.200 ;
    END
  END reg1_val1[28]
  PIN reg1_val1[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 437.960 2200.000 438.560 ;
    END
  END reg1_val1[29]
  PIN reg1_val1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 401.240 2200.000 401.840 ;
    END
  END reg1_val1[2]
  PIN reg1_val1[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 439.320 2200.000 439.920 ;
    END
  END reg1_val1[30]
  PIN reg1_val1[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 440.680 2200.000 441.280 ;
    END
  END reg1_val1[31]
  PIN reg1_val1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 402.600 2200.000 403.200 ;
    END
  END reg1_val1[3]
  PIN reg1_val1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 403.960 2200.000 404.560 ;
    END
  END reg1_val1[4]
  PIN reg1_val1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 405.320 2200.000 405.920 ;
    END
  END reg1_val1[5]
  PIN reg1_val1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 406.680 2200.000 407.280 ;
    END
  END reg1_val1[6]
  PIN reg1_val1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 408.040 2200.000 408.640 ;
    END
  END reg1_val1[7]
  PIN reg1_val1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 409.400 2200.000 410.000 ;
    END
  END reg1_val1[8]
  PIN reg1_val1[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 410.760 2200.000 411.360 ;
    END
  END reg1_val1[9]
  PIN reg1_val2[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 466.520 4.000 467.120 ;
    END
  END reg1_val2[0]
  PIN reg1_val2[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 493.720 4.000 494.320 ;
    END
  END reg1_val2[10]
  PIN reg1_val2[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 496.440 4.000 497.040 ;
    END
  END reg1_val2[11]
  PIN reg1_val2[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 499.160 4.000 499.760 ;
    END
  END reg1_val2[12]
  PIN reg1_val2[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 501.880 4.000 502.480 ;
    END
  END reg1_val2[13]
  PIN reg1_val2[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 504.600 4.000 505.200 ;
    END
  END reg1_val2[14]
  PIN reg1_val2[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 507.320 4.000 507.920 ;
    END
  END reg1_val2[15]
  PIN reg1_val2[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 510.040 4.000 510.640 ;
    END
  END reg1_val2[16]
  PIN reg1_val2[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 512.760 4.000 513.360 ;
    END
  END reg1_val2[17]
  PIN reg1_val2[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 515.480 4.000 516.080 ;
    END
  END reg1_val2[18]
  PIN reg1_val2[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 518.200 4.000 518.800 ;
    END
  END reg1_val2[19]
  PIN reg1_val2[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 469.240 4.000 469.840 ;
    END
  END reg1_val2[1]
  PIN reg1_val2[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 520.920 4.000 521.520 ;
    END
  END reg1_val2[20]
  PIN reg1_val2[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 523.640 4.000 524.240 ;
    END
  END reg1_val2[21]
  PIN reg1_val2[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 526.360 4.000 526.960 ;
    END
  END reg1_val2[22]
  PIN reg1_val2[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 529.080 4.000 529.680 ;
    END
  END reg1_val2[23]
  PIN reg1_val2[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 531.800 4.000 532.400 ;
    END
  END reg1_val2[24]
  PIN reg1_val2[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 534.520 4.000 535.120 ;
    END
  END reg1_val2[25]
  PIN reg1_val2[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 537.240 4.000 537.840 ;
    END
  END reg1_val2[26]
  PIN reg1_val2[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 539.960 4.000 540.560 ;
    END
  END reg1_val2[27]
  PIN reg1_val2[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 542.680 4.000 543.280 ;
    END
  END reg1_val2[28]
  PIN reg1_val2[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 545.400 4.000 546.000 ;
    END
  END reg1_val2[29]
  PIN reg1_val2[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 471.960 4.000 472.560 ;
    END
  END reg1_val2[2]
  PIN reg1_val2[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 548.120 4.000 548.720 ;
    END
  END reg1_val2[30]
  PIN reg1_val2[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 550.840 4.000 551.440 ;
    END
  END reg1_val2[31]
  PIN reg1_val2[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 474.680 4.000 475.280 ;
    END
  END reg1_val2[3]
  PIN reg1_val2[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 477.400 4.000 478.000 ;
    END
  END reg1_val2[4]
  PIN reg1_val2[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 480.120 4.000 480.720 ;
    END
  END reg1_val2[5]
  PIN reg1_val2[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 482.840 4.000 483.440 ;
    END
  END reg1_val2[6]
  PIN reg1_val2[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 485.560 4.000 486.160 ;
    END
  END reg1_val2[7]
  PIN reg1_val2[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 488.280 4.000 488.880 ;
    END
  END reg1_val2[8]
  PIN reg1_val2[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 491.000 4.000 491.600 ;
    END
  END reg1_val2[9]
  PIN reg2_idx0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 998.290 646.000 998.570 650.000 ;
    END
  END reg2_idx0[0]
  PIN reg2_idx0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.337000 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met2 ;
        RECT 1003.350 646.000 1003.630 650.000 ;
    END
  END reg2_idx0[1]
  PIN reg2_idx0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.684000 ;
    PORT
      LAYER met2 ;
        RECT 1008.410 646.000 1008.690 650.000 ;
    END
  END reg2_idx0[2]
  PIN reg2_idx0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.383000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1013.470 646.000 1013.750 650.000 ;
    END
  END reg2_idx0[3]
  PIN reg2_idx0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.293000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1018.530 646.000 1018.810 650.000 ;
    END
  END reg2_idx0[4]
  PIN reg2_idx1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.524500 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 174.120 2200.000 174.720 ;
    END
  END reg2_idx1[0]
  PIN reg2_idx1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.347000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 175.480 2200.000 176.080 ;
    END
  END reg2_idx1[1]
  PIN reg2_idx1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.189000 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 176.840 2200.000 177.440 ;
    END
  END reg2_idx1[2]
  PIN reg2_idx1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.383000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 178.200 2200.000 178.800 ;
    END
  END reg2_idx1[3]
  PIN reg2_idx1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.293000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 179.560 2200.000 180.160 ;
    END
  END reg2_idx1[4]
  PIN reg2_idx2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.732500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.720 4.000 18.320 ;
    END
  END reg2_idx2[0]
  PIN reg2_idx2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.481000 ;
    ANTENNADIFFAREA 3.477600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END reg2_idx2[1]
  PIN reg2_idx2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.722500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.160 4.000 23.760 ;
    END
  END reg2_idx2[2]
  PIN reg2_idx2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.383000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 4.000 26.480 ;
    END
  END reg2_idx2[3]
  PIN reg2_idx2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.293000 ;
    ANTENNADIFFAREA 5.216400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.600 4.000 29.200 ;
    END
  END reg2_idx2[4]
  PIN reg2_val0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1995.110 646.000 1995.390 650.000 ;
    END
  END reg2_val0[0]
  PIN reg2_val0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 2045.710 646.000 2045.990 650.000 ;
    END
  END reg2_val0[10]
  PIN reg2_val0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 2050.770 646.000 2051.050 650.000 ;
    END
  END reg2_val0[11]
  PIN reg2_val0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 2055.830 646.000 2056.110 650.000 ;
    END
  END reg2_val0[12]
  PIN reg2_val0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 2060.890 646.000 2061.170 650.000 ;
    END
  END reg2_val0[13]
  PIN reg2_val0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 2065.950 646.000 2066.230 650.000 ;
    END
  END reg2_val0[14]
  PIN reg2_val0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 2071.010 646.000 2071.290 650.000 ;
    END
  END reg2_val0[15]
  PIN reg2_val0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 2076.070 646.000 2076.350 650.000 ;
    END
  END reg2_val0[16]
  PIN reg2_val0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 2081.130 646.000 2081.410 650.000 ;
    END
  END reg2_val0[17]
  PIN reg2_val0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 2086.190 646.000 2086.470 650.000 ;
    END
  END reg2_val0[18]
  PIN reg2_val0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 2091.250 646.000 2091.530 650.000 ;
    END
  END reg2_val0[19]
  PIN reg2_val0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 2000.170 646.000 2000.450 650.000 ;
    END
  END reg2_val0[1]
  PIN reg2_val0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 2096.310 646.000 2096.590 650.000 ;
    END
  END reg2_val0[20]
  PIN reg2_val0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 2101.370 646.000 2101.650 650.000 ;
    END
  END reg2_val0[21]
  PIN reg2_val0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 2106.430 646.000 2106.710 650.000 ;
    END
  END reg2_val0[22]
  PIN reg2_val0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 2111.490 646.000 2111.770 650.000 ;
    END
  END reg2_val0[23]
  PIN reg2_val0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 2116.550 646.000 2116.830 650.000 ;
    END
  END reg2_val0[24]
  PIN reg2_val0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 2121.610 646.000 2121.890 650.000 ;
    END
  END reg2_val0[25]
  PIN reg2_val0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 2126.670 646.000 2126.950 650.000 ;
    END
  END reg2_val0[26]
  PIN reg2_val0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 2131.730 646.000 2132.010 650.000 ;
    END
  END reg2_val0[27]
  PIN reg2_val0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 2136.790 646.000 2137.070 650.000 ;
    END
  END reg2_val0[28]
  PIN reg2_val0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 2141.850 646.000 2142.130 650.000 ;
    END
  END reg2_val0[29]
  PIN reg2_val0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 2005.230 646.000 2005.510 650.000 ;
    END
  END reg2_val0[2]
  PIN reg2_val0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 2146.910 646.000 2147.190 650.000 ;
    END
  END reg2_val0[30]
  PIN reg2_val0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 2151.970 646.000 2152.250 650.000 ;
    END
  END reg2_val0[31]
  PIN reg2_val0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 2010.290 646.000 2010.570 650.000 ;
    END
  END reg2_val0[3]
  PIN reg2_val0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 2015.350 646.000 2015.630 650.000 ;
    END
  END reg2_val0[4]
  PIN reg2_val0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 2020.410 646.000 2020.690 650.000 ;
    END
  END reg2_val0[5]
  PIN reg2_val0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 2025.470 646.000 2025.750 650.000 ;
    END
  END reg2_val0[6]
  PIN reg2_val0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 2030.530 646.000 2030.810 650.000 ;
    END
  END reg2_val0[7]
  PIN reg2_val0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 2035.590 646.000 2035.870 650.000 ;
    END
  END reg2_val0[8]
  PIN reg2_val0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 2040.650 646.000 2040.930 650.000 ;
    END
  END reg2_val0[9]
  PIN reg2_val1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 442.040 2200.000 442.640 ;
    END
  END reg2_val1[0]
  PIN reg2_val1[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 455.640 2200.000 456.240 ;
    END
  END reg2_val1[10]
  PIN reg2_val1[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 457.000 2200.000 457.600 ;
    END
  END reg2_val1[11]
  PIN reg2_val1[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 458.360 2200.000 458.960 ;
    END
  END reg2_val1[12]
  PIN reg2_val1[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 459.720 2200.000 460.320 ;
    END
  END reg2_val1[13]
  PIN reg2_val1[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 461.080 2200.000 461.680 ;
    END
  END reg2_val1[14]
  PIN reg2_val1[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 462.440 2200.000 463.040 ;
    END
  END reg2_val1[15]
  PIN reg2_val1[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 463.800 2200.000 464.400 ;
    END
  END reg2_val1[16]
  PIN reg2_val1[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 465.160 2200.000 465.760 ;
    END
  END reg2_val1[17]
  PIN reg2_val1[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 466.520 2200.000 467.120 ;
    END
  END reg2_val1[18]
  PIN reg2_val1[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 467.880 2200.000 468.480 ;
    END
  END reg2_val1[19]
  PIN reg2_val1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 443.400 2200.000 444.000 ;
    END
  END reg2_val1[1]
  PIN reg2_val1[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 469.240 2200.000 469.840 ;
    END
  END reg2_val1[20]
  PIN reg2_val1[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 470.600 2200.000 471.200 ;
    END
  END reg2_val1[21]
  PIN reg2_val1[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 471.960 2200.000 472.560 ;
    END
  END reg2_val1[22]
  PIN reg2_val1[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 473.320 2200.000 473.920 ;
    END
  END reg2_val1[23]
  PIN reg2_val1[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 474.680 2200.000 475.280 ;
    END
  END reg2_val1[24]
  PIN reg2_val1[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 476.040 2200.000 476.640 ;
    END
  END reg2_val1[25]
  PIN reg2_val1[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 477.400 2200.000 478.000 ;
    END
  END reg2_val1[26]
  PIN reg2_val1[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 478.760 2200.000 479.360 ;
    END
  END reg2_val1[27]
  PIN reg2_val1[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 480.120 2200.000 480.720 ;
    END
  END reg2_val1[28]
  PIN reg2_val1[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 481.480 2200.000 482.080 ;
    END
  END reg2_val1[29]
  PIN reg2_val1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 444.760 2200.000 445.360 ;
    END
  END reg2_val1[2]
  PIN reg2_val1[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 482.840 2200.000 483.440 ;
    END
  END reg2_val1[30]
  PIN reg2_val1[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 484.200 2200.000 484.800 ;
    END
  END reg2_val1[31]
  PIN reg2_val1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 446.120 2200.000 446.720 ;
    END
  END reg2_val1[3]
  PIN reg2_val1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 447.480 2200.000 448.080 ;
    END
  END reg2_val1[4]
  PIN reg2_val1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 448.840 2200.000 449.440 ;
    END
  END reg2_val1[5]
  PIN reg2_val1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 450.200 2200.000 450.800 ;
    END
  END reg2_val1[6]
  PIN reg2_val1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 451.560 2200.000 452.160 ;
    END
  END reg2_val1[7]
  PIN reg2_val1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 452.920 2200.000 453.520 ;
    END
  END reg2_val1[8]
  PIN reg2_val1[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 454.280 2200.000 454.880 ;
    END
  END reg2_val1[9]
  PIN reg2_val2[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 553.560 4.000 554.160 ;
    END
  END reg2_val2[0]
  PIN reg2_val2[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 580.760 4.000 581.360 ;
    END
  END reg2_val2[10]
  PIN reg2_val2[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 583.480 4.000 584.080 ;
    END
  END reg2_val2[11]
  PIN reg2_val2[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 586.200 4.000 586.800 ;
    END
  END reg2_val2[12]
  PIN reg2_val2[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 588.920 4.000 589.520 ;
    END
  END reg2_val2[13]
  PIN reg2_val2[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 591.640 4.000 592.240 ;
    END
  END reg2_val2[14]
  PIN reg2_val2[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 594.360 4.000 594.960 ;
    END
  END reg2_val2[15]
  PIN reg2_val2[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 597.080 4.000 597.680 ;
    END
  END reg2_val2[16]
  PIN reg2_val2[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 599.800 4.000 600.400 ;
    END
  END reg2_val2[17]
  PIN reg2_val2[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 602.520 4.000 603.120 ;
    END
  END reg2_val2[18]
  PIN reg2_val2[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 605.240 4.000 605.840 ;
    END
  END reg2_val2[19]
  PIN reg2_val2[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 556.280 4.000 556.880 ;
    END
  END reg2_val2[1]
  PIN reg2_val2[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 607.960 4.000 608.560 ;
    END
  END reg2_val2[20]
  PIN reg2_val2[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 610.680 4.000 611.280 ;
    END
  END reg2_val2[21]
  PIN reg2_val2[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 613.400 4.000 614.000 ;
    END
  END reg2_val2[22]
  PIN reg2_val2[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 616.120 4.000 616.720 ;
    END
  END reg2_val2[23]
  PIN reg2_val2[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 618.840 4.000 619.440 ;
    END
  END reg2_val2[24]
  PIN reg2_val2[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 621.560 4.000 622.160 ;
    END
  END reg2_val2[25]
  PIN reg2_val2[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 624.280 4.000 624.880 ;
    END
  END reg2_val2[26]
  PIN reg2_val2[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 627.000 4.000 627.600 ;
    END
  END reg2_val2[27]
  PIN reg2_val2[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 629.720 4.000 630.320 ;
    END
  END reg2_val2[28]
  PIN reg2_val2[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 632.440 4.000 633.040 ;
    END
  END reg2_val2[29]
  PIN reg2_val2[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 559.000 4.000 559.600 ;
    END
  END reg2_val2[2]
  PIN reg2_val2[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 635.160 4.000 635.760 ;
    END
  END reg2_val2[30]
  PIN reg2_val2[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 637.880 4.000 638.480 ;
    END
  END reg2_val2[31]
  PIN reg2_val2[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 561.720 4.000 562.320 ;
    END
  END reg2_val2[3]
  PIN reg2_val2[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 564.440 4.000 565.040 ;
    END
  END reg2_val2[4]
  PIN reg2_val2[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 567.160 4.000 567.760 ;
    END
  END reg2_val2[5]
  PIN reg2_val2[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 569.880 4.000 570.480 ;
    END
  END reg2_val2[6]
  PIN reg2_val2[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 572.600 4.000 573.200 ;
    END
  END reg2_val2[7]
  PIN reg2_val2[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 575.320 4.000 575.920 ;
    END
  END reg2_val2[8]
  PIN reg2_val2[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 578.040 4.000 578.640 ;
    END
  END reg2_val2[9]
  PIN rst_eu
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.862000 ;
    PORT
      LAYER met2 ;
        RECT 826.250 646.000 826.530 650.000 ;
    END
  END rst_eu
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.086000 ;
    PORT
      LAYER met2 ;
        RECT 2113.330 0.000 2113.610 4.000 ;
    END
  END rst_n
  PIN sign_extend0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1428.390 646.000 1428.670 650.000 ;
    END
  END sign_extend0
  PIN sign_extend1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 7.824600 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 289.720 2200.000 290.320 ;
    END
  END sign_extend1
  PIN sign_extend2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 24.777899 ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.920 4.000 249.520 ;
    END
  END sign_extend2
  PIN take_branch0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.485000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1468.870 646.000 1469.150 650.000 ;
    END
  END take_branch0
  PIN take_branch1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.406000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 300.600 2200.000 301.200 ;
    END
  END take_branch1
  PIN take_branch2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 270.680 4.000 271.280 ;
    END
  END take_branch2
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 636.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 636.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 636.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 636.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 636.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 636.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 636.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 636.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 636.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 636.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.040 10.640 1558.640 636.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1710.640 10.640 1712.240 636.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1864.240 10.640 1865.840 636.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 2017.840 10.640 2019.440 636.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 2171.440 10.640 2173.040 636.720 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 636.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 636.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 636.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 636.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 636.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 636.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 636.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 636.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 636.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 636.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1633.840 10.640 1635.440 636.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1787.440 10.640 1789.040 636.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1941.040 10.640 1942.640 636.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 2094.640 10.640 2096.240 636.720 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 2104.590 0.000 2104.870 4.000 ;
    END
  END wb_clk_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2194.200 636.565 ;
      LAYER met1 ;
        RECT 5.520 10.240 2197.350 649.980 ;
      LAYER met2 ;
        RECT 15.730 645.720 36.610 649.925 ;
        RECT 37.450 645.720 41.670 649.925 ;
        RECT 42.510 645.720 46.730 649.925 ;
        RECT 47.570 645.720 51.790 649.925 ;
        RECT 52.630 645.720 56.850 649.925 ;
        RECT 57.690 645.720 61.910 649.925 ;
        RECT 62.750 645.720 66.970 649.925 ;
        RECT 67.810 645.720 72.030 649.925 ;
        RECT 72.870 645.720 77.090 649.925 ;
        RECT 77.930 645.720 82.150 649.925 ;
        RECT 82.990 645.720 87.210 649.925 ;
        RECT 88.050 645.720 92.270 649.925 ;
        RECT 93.110 645.720 97.330 649.925 ;
        RECT 98.170 645.720 102.390 649.925 ;
        RECT 103.230 645.720 107.450 649.925 ;
        RECT 108.290 645.720 112.510 649.925 ;
        RECT 113.350 645.720 117.570 649.925 ;
        RECT 118.410 645.720 122.630 649.925 ;
        RECT 123.470 645.720 127.690 649.925 ;
        RECT 128.530 645.720 132.750 649.925 ;
        RECT 133.590 645.720 137.810 649.925 ;
        RECT 138.650 645.720 142.870 649.925 ;
        RECT 143.710 645.720 147.930 649.925 ;
        RECT 148.770 645.720 152.990 649.925 ;
        RECT 153.830 645.720 158.050 649.925 ;
        RECT 158.890 645.720 163.110 649.925 ;
        RECT 163.950 645.720 168.170 649.925 ;
        RECT 169.010 645.720 173.230 649.925 ;
        RECT 174.070 645.720 178.290 649.925 ;
        RECT 179.130 645.720 183.350 649.925 ;
        RECT 184.190 645.720 188.410 649.925 ;
        RECT 189.250 645.720 193.470 649.925 ;
        RECT 194.310 645.720 198.530 649.925 ;
        RECT 199.370 645.720 203.590 649.925 ;
        RECT 204.430 645.720 208.650 649.925 ;
        RECT 209.490 645.720 213.710 649.925 ;
        RECT 214.550 645.720 218.770 649.925 ;
        RECT 219.610 645.720 223.830 649.925 ;
        RECT 224.670 645.720 228.890 649.925 ;
        RECT 229.730 645.720 233.950 649.925 ;
        RECT 234.790 645.720 239.010 649.925 ;
        RECT 239.850 645.720 244.070 649.925 ;
        RECT 244.910 645.720 249.130 649.925 ;
        RECT 249.970 645.720 254.190 649.925 ;
        RECT 255.030 645.720 259.250 649.925 ;
        RECT 260.090 645.720 264.310 649.925 ;
        RECT 265.150 645.720 269.370 649.925 ;
        RECT 270.210 645.720 274.430 649.925 ;
        RECT 275.270 645.720 279.490 649.925 ;
        RECT 280.330 645.720 284.550 649.925 ;
        RECT 285.390 645.720 289.610 649.925 ;
        RECT 290.450 645.720 294.670 649.925 ;
        RECT 295.510 645.720 299.730 649.925 ;
        RECT 300.570 645.720 304.790 649.925 ;
        RECT 305.630 645.720 309.850 649.925 ;
        RECT 310.690 645.720 314.910 649.925 ;
        RECT 315.750 645.720 319.970 649.925 ;
        RECT 320.810 645.720 325.030 649.925 ;
        RECT 325.870 645.720 330.090 649.925 ;
        RECT 330.930 645.720 335.150 649.925 ;
        RECT 335.990 645.720 340.210 649.925 ;
        RECT 341.050 645.720 345.270 649.925 ;
        RECT 346.110 645.720 350.330 649.925 ;
        RECT 351.170 645.720 355.390 649.925 ;
        RECT 356.230 645.720 360.450 649.925 ;
        RECT 361.290 645.720 365.510 649.925 ;
        RECT 366.350 645.720 370.570 649.925 ;
        RECT 371.410 645.720 375.630 649.925 ;
        RECT 376.470 645.720 380.690 649.925 ;
        RECT 381.530 645.720 385.750 649.925 ;
        RECT 386.590 645.720 390.810 649.925 ;
        RECT 391.650 645.720 395.870 649.925 ;
        RECT 396.710 645.720 400.930 649.925 ;
        RECT 401.770 645.720 405.990 649.925 ;
        RECT 406.830 645.720 411.050 649.925 ;
        RECT 411.890 645.720 416.110 649.925 ;
        RECT 416.950 645.720 421.170 649.925 ;
        RECT 422.010 645.720 426.230 649.925 ;
        RECT 427.070 645.720 431.290 649.925 ;
        RECT 432.130 645.720 436.350 649.925 ;
        RECT 437.190 645.720 441.410 649.925 ;
        RECT 442.250 645.720 446.470 649.925 ;
        RECT 447.310 645.720 451.530 649.925 ;
        RECT 452.370 645.720 456.590 649.925 ;
        RECT 457.430 645.720 461.650 649.925 ;
        RECT 462.490 645.720 466.710 649.925 ;
        RECT 467.550 645.720 471.770 649.925 ;
        RECT 472.610 645.720 476.830 649.925 ;
        RECT 477.670 645.720 481.890 649.925 ;
        RECT 482.730 645.720 486.950 649.925 ;
        RECT 487.790 645.720 492.010 649.925 ;
        RECT 492.850 645.720 497.070 649.925 ;
        RECT 497.910 645.720 502.130 649.925 ;
        RECT 502.970 645.720 507.190 649.925 ;
        RECT 508.030 645.720 512.250 649.925 ;
        RECT 513.090 645.720 517.310 649.925 ;
        RECT 518.150 645.720 522.370 649.925 ;
        RECT 523.210 645.720 527.430 649.925 ;
        RECT 528.270 645.720 532.490 649.925 ;
        RECT 533.330 645.720 537.550 649.925 ;
        RECT 538.390 645.720 542.610 649.925 ;
        RECT 543.450 645.720 547.670 649.925 ;
        RECT 548.510 645.720 552.730 649.925 ;
        RECT 553.570 645.720 557.790 649.925 ;
        RECT 558.630 645.720 562.850 649.925 ;
        RECT 563.690 645.720 567.910 649.925 ;
        RECT 568.750 645.720 572.970 649.925 ;
        RECT 573.810 645.720 578.030 649.925 ;
        RECT 578.870 645.720 583.090 649.925 ;
        RECT 583.930 645.720 588.150 649.925 ;
        RECT 588.990 645.720 593.210 649.925 ;
        RECT 594.050 645.720 598.270 649.925 ;
        RECT 599.110 645.720 603.330 649.925 ;
        RECT 604.170 645.720 608.390 649.925 ;
        RECT 609.230 645.720 613.450 649.925 ;
        RECT 614.290 645.720 618.510 649.925 ;
        RECT 619.350 645.720 623.570 649.925 ;
        RECT 624.410 645.720 628.630 649.925 ;
        RECT 629.470 645.720 633.690 649.925 ;
        RECT 634.530 645.720 638.750 649.925 ;
        RECT 639.590 645.720 643.810 649.925 ;
        RECT 644.650 645.720 648.870 649.925 ;
        RECT 649.710 645.720 653.930 649.925 ;
        RECT 654.770 645.720 658.990 649.925 ;
        RECT 659.830 645.720 664.050 649.925 ;
        RECT 664.890 645.720 669.110 649.925 ;
        RECT 669.950 645.720 674.170 649.925 ;
        RECT 675.010 645.720 679.230 649.925 ;
        RECT 680.070 645.720 684.290 649.925 ;
        RECT 685.130 645.720 689.350 649.925 ;
        RECT 690.190 645.720 694.410 649.925 ;
        RECT 695.250 645.720 699.470 649.925 ;
        RECT 700.310 645.720 704.530 649.925 ;
        RECT 705.370 645.720 709.590 649.925 ;
        RECT 710.430 645.720 714.650 649.925 ;
        RECT 715.490 645.720 719.710 649.925 ;
        RECT 720.550 645.720 724.770 649.925 ;
        RECT 725.610 645.720 729.830 649.925 ;
        RECT 730.670 645.720 734.890 649.925 ;
        RECT 735.730 645.720 739.950 649.925 ;
        RECT 740.790 645.720 745.010 649.925 ;
        RECT 745.850 645.720 750.070 649.925 ;
        RECT 750.910 645.720 755.130 649.925 ;
        RECT 755.970 645.720 760.190 649.925 ;
        RECT 761.030 645.720 765.250 649.925 ;
        RECT 766.090 645.720 770.310 649.925 ;
        RECT 771.150 645.720 775.370 649.925 ;
        RECT 776.210 645.720 780.430 649.925 ;
        RECT 781.270 645.720 785.490 649.925 ;
        RECT 786.330 645.720 790.550 649.925 ;
        RECT 791.390 645.720 795.610 649.925 ;
        RECT 796.450 645.720 800.670 649.925 ;
        RECT 801.510 645.720 805.730 649.925 ;
        RECT 806.570 645.720 810.790 649.925 ;
        RECT 811.630 645.720 815.850 649.925 ;
        RECT 816.690 645.720 820.910 649.925 ;
        RECT 821.750 645.720 825.970 649.925 ;
        RECT 826.810 645.720 831.030 649.925 ;
        RECT 831.870 645.720 836.090 649.925 ;
        RECT 836.930 645.720 841.150 649.925 ;
        RECT 841.990 645.720 846.210 649.925 ;
        RECT 847.050 645.720 851.270 649.925 ;
        RECT 852.110 645.720 856.330 649.925 ;
        RECT 857.170 645.720 861.390 649.925 ;
        RECT 862.230 645.720 866.450 649.925 ;
        RECT 867.290 645.720 871.510 649.925 ;
        RECT 872.350 645.720 876.570 649.925 ;
        RECT 877.410 645.720 881.630 649.925 ;
        RECT 882.470 645.720 886.690 649.925 ;
        RECT 887.530 645.720 891.750 649.925 ;
        RECT 892.590 645.720 896.810 649.925 ;
        RECT 897.650 645.720 901.870 649.925 ;
        RECT 902.710 645.720 906.930 649.925 ;
        RECT 907.770 645.720 911.990 649.925 ;
        RECT 912.830 645.720 917.050 649.925 ;
        RECT 917.890 645.720 922.110 649.925 ;
        RECT 922.950 645.720 927.170 649.925 ;
        RECT 928.010 645.720 932.230 649.925 ;
        RECT 933.070 645.720 937.290 649.925 ;
        RECT 938.130 645.720 942.350 649.925 ;
        RECT 943.190 645.720 947.410 649.925 ;
        RECT 948.250 645.720 952.470 649.925 ;
        RECT 953.310 645.720 957.530 649.925 ;
        RECT 958.370 645.720 962.590 649.925 ;
        RECT 963.430 645.720 967.650 649.925 ;
        RECT 968.490 645.720 972.710 649.925 ;
        RECT 973.550 645.720 977.770 649.925 ;
        RECT 978.610 645.720 982.830 649.925 ;
        RECT 983.670 645.720 987.890 649.925 ;
        RECT 988.730 645.720 992.950 649.925 ;
        RECT 993.790 645.720 998.010 649.925 ;
        RECT 998.850 645.720 1003.070 649.925 ;
        RECT 1003.910 645.720 1008.130 649.925 ;
        RECT 1008.970 645.720 1013.190 649.925 ;
        RECT 1014.030 645.720 1018.250 649.925 ;
        RECT 1019.090 645.720 1023.310 649.925 ;
        RECT 1024.150 645.720 1028.370 649.925 ;
        RECT 1029.210 645.720 1033.430 649.925 ;
        RECT 1034.270 645.720 1038.490 649.925 ;
        RECT 1039.330 645.720 1043.550 649.925 ;
        RECT 1044.390 645.720 1048.610 649.925 ;
        RECT 1049.450 645.720 1053.670 649.925 ;
        RECT 1054.510 645.720 1058.730 649.925 ;
        RECT 1059.570 645.720 1063.790 649.925 ;
        RECT 1064.630 645.720 1068.850 649.925 ;
        RECT 1069.690 645.720 1073.910 649.925 ;
        RECT 1074.750 645.720 1078.970 649.925 ;
        RECT 1079.810 645.720 1084.030 649.925 ;
        RECT 1084.870 645.720 1089.090 649.925 ;
        RECT 1089.930 645.720 1094.150 649.925 ;
        RECT 1094.990 645.720 1099.210 649.925 ;
        RECT 1100.050 645.720 1104.270 649.925 ;
        RECT 1105.110 645.720 1109.330 649.925 ;
        RECT 1110.170 645.720 1114.390 649.925 ;
        RECT 1115.230 645.720 1119.450 649.925 ;
        RECT 1120.290 645.720 1124.510 649.925 ;
        RECT 1125.350 645.720 1129.570 649.925 ;
        RECT 1130.410 645.720 1134.630 649.925 ;
        RECT 1135.470 645.720 1139.690 649.925 ;
        RECT 1140.530 645.720 1144.750 649.925 ;
        RECT 1145.590 645.720 1149.810 649.925 ;
        RECT 1150.650 645.720 1154.870 649.925 ;
        RECT 1155.710 645.720 1159.930 649.925 ;
        RECT 1160.770 645.720 1164.990 649.925 ;
        RECT 1165.830 645.720 1170.050 649.925 ;
        RECT 1170.890 645.720 1175.110 649.925 ;
        RECT 1175.950 645.720 1180.170 649.925 ;
        RECT 1181.010 645.720 1185.230 649.925 ;
        RECT 1186.070 645.720 1190.290 649.925 ;
        RECT 1191.130 645.720 1195.350 649.925 ;
        RECT 1196.190 645.720 1200.410 649.925 ;
        RECT 1201.250 645.720 1205.470 649.925 ;
        RECT 1206.310 645.720 1210.530 649.925 ;
        RECT 1211.370 645.720 1215.590 649.925 ;
        RECT 1216.430 645.720 1220.650 649.925 ;
        RECT 1221.490 645.720 1225.710 649.925 ;
        RECT 1226.550 645.720 1230.770 649.925 ;
        RECT 1231.610 645.720 1235.830 649.925 ;
        RECT 1236.670 645.720 1240.890 649.925 ;
        RECT 1241.730 645.720 1245.950 649.925 ;
        RECT 1246.790 645.720 1251.010 649.925 ;
        RECT 1251.850 645.720 1256.070 649.925 ;
        RECT 1256.910 645.720 1261.130 649.925 ;
        RECT 1261.970 645.720 1266.190 649.925 ;
        RECT 1267.030 645.720 1271.250 649.925 ;
        RECT 1272.090 645.720 1276.310 649.925 ;
        RECT 1277.150 645.720 1281.370 649.925 ;
        RECT 1282.210 645.720 1286.430 649.925 ;
        RECT 1287.270 645.720 1291.490 649.925 ;
        RECT 1292.330 645.720 1296.550 649.925 ;
        RECT 1297.390 645.720 1301.610 649.925 ;
        RECT 1302.450 645.720 1306.670 649.925 ;
        RECT 1307.510 645.720 1311.730 649.925 ;
        RECT 1312.570 645.720 1316.790 649.925 ;
        RECT 1317.630 645.720 1321.850 649.925 ;
        RECT 1322.690 645.720 1326.910 649.925 ;
        RECT 1327.750 645.720 1331.970 649.925 ;
        RECT 1332.810 645.720 1337.030 649.925 ;
        RECT 1337.870 645.720 1342.090 649.925 ;
        RECT 1342.930 645.720 1347.150 649.925 ;
        RECT 1347.990 645.720 1352.210 649.925 ;
        RECT 1353.050 645.720 1357.270 649.925 ;
        RECT 1358.110 645.720 1362.330 649.925 ;
        RECT 1363.170 645.720 1367.390 649.925 ;
        RECT 1368.230 645.720 1372.450 649.925 ;
        RECT 1373.290 645.720 1377.510 649.925 ;
        RECT 1378.350 645.720 1382.570 649.925 ;
        RECT 1383.410 645.720 1387.630 649.925 ;
        RECT 1388.470 645.720 1392.690 649.925 ;
        RECT 1393.530 645.720 1397.750 649.925 ;
        RECT 1398.590 645.720 1402.810 649.925 ;
        RECT 1403.650 645.720 1407.870 649.925 ;
        RECT 1408.710 645.720 1412.930 649.925 ;
        RECT 1413.770 645.720 1417.990 649.925 ;
        RECT 1418.830 645.720 1423.050 649.925 ;
        RECT 1423.890 645.720 1428.110 649.925 ;
        RECT 1428.950 645.720 1433.170 649.925 ;
        RECT 1434.010 645.720 1438.230 649.925 ;
        RECT 1439.070 645.720 1443.290 649.925 ;
        RECT 1444.130 645.720 1448.350 649.925 ;
        RECT 1449.190 645.720 1453.410 649.925 ;
        RECT 1454.250 645.720 1458.470 649.925 ;
        RECT 1459.310 645.720 1463.530 649.925 ;
        RECT 1464.370 645.720 1468.590 649.925 ;
        RECT 1469.430 645.720 1473.650 649.925 ;
        RECT 1474.490 645.720 1478.710 649.925 ;
        RECT 1479.550 645.720 1483.770 649.925 ;
        RECT 1484.610 645.720 1488.830 649.925 ;
        RECT 1489.670 645.720 1493.890 649.925 ;
        RECT 1494.730 645.720 1498.950 649.925 ;
        RECT 1499.790 645.720 1504.010 649.925 ;
        RECT 1504.850 645.720 1509.070 649.925 ;
        RECT 1509.910 645.720 1514.130 649.925 ;
        RECT 1514.970 645.720 1519.190 649.925 ;
        RECT 1520.030 645.720 1524.250 649.925 ;
        RECT 1525.090 645.720 1529.310 649.925 ;
        RECT 1530.150 645.720 1534.370 649.925 ;
        RECT 1535.210 645.720 1539.430 649.925 ;
        RECT 1540.270 645.720 1544.490 649.925 ;
        RECT 1545.330 645.720 1549.550 649.925 ;
        RECT 1550.390 645.720 1554.610 649.925 ;
        RECT 1555.450 645.720 1559.670 649.925 ;
        RECT 1560.510 645.720 1564.730 649.925 ;
        RECT 1565.570 645.720 1569.790 649.925 ;
        RECT 1570.630 645.720 1574.850 649.925 ;
        RECT 1575.690 645.720 1579.910 649.925 ;
        RECT 1580.750 645.720 1584.970 649.925 ;
        RECT 1585.810 645.720 1590.030 649.925 ;
        RECT 1590.870 645.720 1595.090 649.925 ;
        RECT 1595.930 645.720 1600.150 649.925 ;
        RECT 1600.990 645.720 1605.210 649.925 ;
        RECT 1606.050 645.720 1610.270 649.925 ;
        RECT 1611.110 645.720 1615.330 649.925 ;
        RECT 1616.170 645.720 1620.390 649.925 ;
        RECT 1621.230 645.720 1625.450 649.925 ;
        RECT 1626.290 645.720 1630.510 649.925 ;
        RECT 1631.350 645.720 1635.570 649.925 ;
        RECT 1636.410 645.720 1640.630 649.925 ;
        RECT 1641.470 645.720 1645.690 649.925 ;
        RECT 1646.530 645.720 1650.750 649.925 ;
        RECT 1651.590 645.720 1655.810 649.925 ;
        RECT 1656.650 645.720 1660.870 649.925 ;
        RECT 1661.710 645.720 1665.930 649.925 ;
        RECT 1666.770 645.720 1670.990 649.925 ;
        RECT 1671.830 645.720 1676.050 649.925 ;
        RECT 1676.890 645.720 1681.110 649.925 ;
        RECT 1681.950 645.720 1686.170 649.925 ;
        RECT 1687.010 645.720 1691.230 649.925 ;
        RECT 1692.070 645.720 1696.290 649.925 ;
        RECT 1697.130 645.720 1701.350 649.925 ;
        RECT 1702.190 645.720 1706.410 649.925 ;
        RECT 1707.250 645.720 1711.470 649.925 ;
        RECT 1712.310 645.720 1716.530 649.925 ;
        RECT 1717.370 645.720 1721.590 649.925 ;
        RECT 1722.430 645.720 1726.650 649.925 ;
        RECT 1727.490 645.720 1731.710 649.925 ;
        RECT 1732.550 645.720 1736.770 649.925 ;
        RECT 1737.610 645.720 1741.830 649.925 ;
        RECT 1742.670 645.720 1746.890 649.925 ;
        RECT 1747.730 645.720 1751.950 649.925 ;
        RECT 1752.790 645.720 1757.010 649.925 ;
        RECT 1757.850 645.720 1762.070 649.925 ;
        RECT 1762.910 645.720 1767.130 649.925 ;
        RECT 1767.970 645.720 1772.190 649.925 ;
        RECT 1773.030 645.720 1777.250 649.925 ;
        RECT 1778.090 645.720 1782.310 649.925 ;
        RECT 1783.150 645.720 1787.370 649.925 ;
        RECT 1788.210 645.720 1792.430 649.925 ;
        RECT 1793.270 645.720 1797.490 649.925 ;
        RECT 1798.330 645.720 1802.550 649.925 ;
        RECT 1803.390 645.720 1807.610 649.925 ;
        RECT 1808.450 645.720 1812.670 649.925 ;
        RECT 1813.510 645.720 1817.730 649.925 ;
        RECT 1818.570 645.720 1822.790 649.925 ;
        RECT 1823.630 645.720 1827.850 649.925 ;
        RECT 1828.690 645.720 1832.910 649.925 ;
        RECT 1833.750 645.720 1837.970 649.925 ;
        RECT 1838.810 645.720 1843.030 649.925 ;
        RECT 1843.870 645.720 1848.090 649.925 ;
        RECT 1848.930 645.720 1853.150 649.925 ;
        RECT 1853.990 645.720 1858.210 649.925 ;
        RECT 1859.050 645.720 1863.270 649.925 ;
        RECT 1864.110 645.720 1868.330 649.925 ;
        RECT 1869.170 645.720 1873.390 649.925 ;
        RECT 1874.230 645.720 1878.450 649.925 ;
        RECT 1879.290 645.720 1883.510 649.925 ;
        RECT 1884.350 645.720 1888.570 649.925 ;
        RECT 1889.410 645.720 1893.630 649.925 ;
        RECT 1894.470 645.720 1898.690 649.925 ;
        RECT 1899.530 645.720 1903.750 649.925 ;
        RECT 1904.590 645.720 1908.810 649.925 ;
        RECT 1909.650 645.720 1913.870 649.925 ;
        RECT 1914.710 645.720 1918.930 649.925 ;
        RECT 1919.770 645.720 1923.990 649.925 ;
        RECT 1924.830 645.720 1929.050 649.925 ;
        RECT 1929.890 645.720 1934.110 649.925 ;
        RECT 1934.950 645.720 1939.170 649.925 ;
        RECT 1940.010 645.720 1944.230 649.925 ;
        RECT 1945.070 645.720 1949.290 649.925 ;
        RECT 1950.130 645.720 1954.350 649.925 ;
        RECT 1955.190 645.720 1959.410 649.925 ;
        RECT 1960.250 645.720 1964.470 649.925 ;
        RECT 1965.310 645.720 1969.530 649.925 ;
        RECT 1970.370 645.720 1974.590 649.925 ;
        RECT 1975.430 645.720 1979.650 649.925 ;
        RECT 1980.490 645.720 1984.710 649.925 ;
        RECT 1985.550 645.720 1989.770 649.925 ;
        RECT 1990.610 645.720 1994.830 649.925 ;
        RECT 1995.670 645.720 1999.890 649.925 ;
        RECT 2000.730 645.720 2004.950 649.925 ;
        RECT 2005.790 645.720 2010.010 649.925 ;
        RECT 2010.850 645.720 2015.070 649.925 ;
        RECT 2015.910 645.720 2020.130 649.925 ;
        RECT 2020.970 645.720 2025.190 649.925 ;
        RECT 2026.030 645.720 2030.250 649.925 ;
        RECT 2031.090 645.720 2035.310 649.925 ;
        RECT 2036.150 645.720 2040.370 649.925 ;
        RECT 2041.210 645.720 2045.430 649.925 ;
        RECT 2046.270 645.720 2050.490 649.925 ;
        RECT 2051.330 645.720 2055.550 649.925 ;
        RECT 2056.390 645.720 2060.610 649.925 ;
        RECT 2061.450 645.720 2065.670 649.925 ;
        RECT 2066.510 645.720 2070.730 649.925 ;
        RECT 2071.570 645.720 2075.790 649.925 ;
        RECT 2076.630 645.720 2080.850 649.925 ;
        RECT 2081.690 645.720 2085.910 649.925 ;
        RECT 2086.750 645.720 2090.970 649.925 ;
        RECT 2091.810 645.720 2096.030 649.925 ;
        RECT 2096.870 645.720 2101.090 649.925 ;
        RECT 2101.930 645.720 2106.150 649.925 ;
        RECT 2106.990 645.720 2111.210 649.925 ;
        RECT 2112.050 645.720 2116.270 649.925 ;
        RECT 2117.110 645.720 2121.330 649.925 ;
        RECT 2122.170 645.720 2126.390 649.925 ;
        RECT 2127.230 645.720 2131.450 649.925 ;
        RECT 2132.290 645.720 2136.510 649.925 ;
        RECT 2137.350 645.720 2141.570 649.925 ;
        RECT 2142.410 645.720 2146.630 649.925 ;
        RECT 2147.470 645.720 2151.690 649.925 ;
        RECT 2152.530 645.720 2156.750 649.925 ;
        RECT 2157.590 645.720 2161.810 649.925 ;
        RECT 2162.650 645.720 2197.320 649.925 ;
        RECT 15.730 4.280 2197.320 645.720 ;
        RECT 15.730 3.670 41.670 4.280 ;
        RECT 42.510 3.670 50.410 4.280 ;
        RECT 51.250 3.670 59.150 4.280 ;
        RECT 59.990 3.670 67.890 4.280 ;
        RECT 68.730 3.670 76.630 4.280 ;
        RECT 77.470 3.670 85.370 4.280 ;
        RECT 86.210 3.670 94.110 4.280 ;
        RECT 94.950 3.670 102.850 4.280 ;
        RECT 103.690 3.670 111.590 4.280 ;
        RECT 112.430 3.670 120.330 4.280 ;
        RECT 121.170 3.670 129.070 4.280 ;
        RECT 129.910 3.670 137.810 4.280 ;
        RECT 138.650 3.670 146.550 4.280 ;
        RECT 147.390 3.670 155.290 4.280 ;
        RECT 156.130 3.670 164.030 4.280 ;
        RECT 164.870 3.670 172.770 4.280 ;
        RECT 173.610 3.670 181.510 4.280 ;
        RECT 182.350 3.670 190.250 4.280 ;
        RECT 191.090 3.670 198.990 4.280 ;
        RECT 199.830 3.670 207.730 4.280 ;
        RECT 208.570 3.670 216.470 4.280 ;
        RECT 217.310 3.670 225.210 4.280 ;
        RECT 226.050 3.670 233.950 4.280 ;
        RECT 234.790 3.670 242.690 4.280 ;
        RECT 243.530 3.670 251.430 4.280 ;
        RECT 252.270 3.670 260.170 4.280 ;
        RECT 261.010 3.670 268.910 4.280 ;
        RECT 269.750 3.670 277.650 4.280 ;
        RECT 278.490 3.670 286.390 4.280 ;
        RECT 287.230 3.670 295.130 4.280 ;
        RECT 295.970 3.670 303.870 4.280 ;
        RECT 304.710 3.670 312.610 4.280 ;
        RECT 313.450 3.670 321.350 4.280 ;
        RECT 322.190 3.670 330.090 4.280 ;
        RECT 330.930 3.670 338.830 4.280 ;
        RECT 339.670 3.670 347.570 4.280 ;
        RECT 348.410 3.670 356.310 4.280 ;
        RECT 357.150 3.670 365.050 4.280 ;
        RECT 365.890 3.670 373.790 4.280 ;
        RECT 374.630 3.670 382.530 4.280 ;
        RECT 383.370 3.670 391.270 4.280 ;
        RECT 392.110 3.670 400.010 4.280 ;
        RECT 400.850 3.670 408.750 4.280 ;
        RECT 409.590 3.670 417.490 4.280 ;
        RECT 418.330 3.670 426.230 4.280 ;
        RECT 427.070 3.670 434.970 4.280 ;
        RECT 435.810 3.670 443.710 4.280 ;
        RECT 444.550 3.670 452.450 4.280 ;
        RECT 453.290 3.670 461.190 4.280 ;
        RECT 462.030 3.670 469.930 4.280 ;
        RECT 470.770 3.670 478.670 4.280 ;
        RECT 479.510 3.670 487.410 4.280 ;
        RECT 488.250 3.670 496.150 4.280 ;
        RECT 496.990 3.670 504.890 4.280 ;
        RECT 505.730 3.670 513.630 4.280 ;
        RECT 514.470 3.670 522.370 4.280 ;
        RECT 523.210 3.670 531.110 4.280 ;
        RECT 531.950 3.670 539.850 4.280 ;
        RECT 540.690 3.670 548.590 4.280 ;
        RECT 549.430 3.670 557.330 4.280 ;
        RECT 558.170 3.670 566.070 4.280 ;
        RECT 566.910 3.670 574.810 4.280 ;
        RECT 575.650 3.670 583.550 4.280 ;
        RECT 584.390 3.670 592.290 4.280 ;
        RECT 593.130 3.670 601.030 4.280 ;
        RECT 601.870 3.670 609.770 4.280 ;
        RECT 610.610 3.670 618.510 4.280 ;
        RECT 619.350 3.670 627.250 4.280 ;
        RECT 628.090 3.670 635.990 4.280 ;
        RECT 636.830 3.670 644.730 4.280 ;
        RECT 645.570 3.670 653.470 4.280 ;
        RECT 654.310 3.670 662.210 4.280 ;
        RECT 663.050 3.670 670.950 4.280 ;
        RECT 671.790 3.670 679.690 4.280 ;
        RECT 680.530 3.670 688.430 4.280 ;
        RECT 689.270 3.670 697.170 4.280 ;
        RECT 698.010 3.670 705.910 4.280 ;
        RECT 706.750 3.670 714.650 4.280 ;
        RECT 715.490 3.670 723.390 4.280 ;
        RECT 724.230 3.670 732.130 4.280 ;
        RECT 732.970 3.670 740.870 4.280 ;
        RECT 741.710 3.670 749.610 4.280 ;
        RECT 750.450 3.670 758.350 4.280 ;
        RECT 759.190 3.670 767.090 4.280 ;
        RECT 767.930 3.670 775.830 4.280 ;
        RECT 776.670 3.670 784.570 4.280 ;
        RECT 785.410 3.670 793.310 4.280 ;
        RECT 794.150 3.670 802.050 4.280 ;
        RECT 802.890 3.670 810.790 4.280 ;
        RECT 811.630 3.670 819.530 4.280 ;
        RECT 820.370 3.670 828.270 4.280 ;
        RECT 829.110 3.670 837.010 4.280 ;
        RECT 837.850 3.670 845.750 4.280 ;
        RECT 846.590 3.670 854.490 4.280 ;
        RECT 855.330 3.670 863.230 4.280 ;
        RECT 864.070 3.670 871.970 4.280 ;
        RECT 872.810 3.670 880.710 4.280 ;
        RECT 881.550 3.670 889.450 4.280 ;
        RECT 890.290 3.670 898.190 4.280 ;
        RECT 899.030 3.670 906.930 4.280 ;
        RECT 907.770 3.670 915.670 4.280 ;
        RECT 916.510 3.670 924.410 4.280 ;
        RECT 925.250 3.670 933.150 4.280 ;
        RECT 933.990 3.670 941.890 4.280 ;
        RECT 942.730 3.670 950.630 4.280 ;
        RECT 951.470 3.670 959.370 4.280 ;
        RECT 960.210 3.670 968.110 4.280 ;
        RECT 968.950 3.670 976.850 4.280 ;
        RECT 977.690 3.670 985.590 4.280 ;
        RECT 986.430 3.670 994.330 4.280 ;
        RECT 995.170 3.670 1003.070 4.280 ;
        RECT 1003.910 3.670 1011.810 4.280 ;
        RECT 1012.650 3.670 1020.550 4.280 ;
        RECT 1021.390 3.670 1029.290 4.280 ;
        RECT 1030.130 3.670 1038.030 4.280 ;
        RECT 1038.870 3.670 1046.770 4.280 ;
        RECT 1047.610 3.670 1055.510 4.280 ;
        RECT 1056.350 3.670 1064.250 4.280 ;
        RECT 1065.090 3.670 1072.990 4.280 ;
        RECT 1073.830 3.670 1081.730 4.280 ;
        RECT 1082.570 3.670 1090.470 4.280 ;
        RECT 1091.310 3.670 1099.210 4.280 ;
        RECT 1100.050 3.670 1107.950 4.280 ;
        RECT 1108.790 3.670 1116.690 4.280 ;
        RECT 1117.530 3.670 1125.430 4.280 ;
        RECT 1126.270 3.670 1134.170 4.280 ;
        RECT 1135.010 3.670 1142.910 4.280 ;
        RECT 1143.750 3.670 1151.650 4.280 ;
        RECT 1152.490 3.670 1160.390 4.280 ;
        RECT 1161.230 3.670 1169.130 4.280 ;
        RECT 1169.970 3.670 1177.870 4.280 ;
        RECT 1178.710 3.670 1186.610 4.280 ;
        RECT 1187.450 3.670 1195.350 4.280 ;
        RECT 1196.190 3.670 1204.090 4.280 ;
        RECT 1204.930 3.670 1212.830 4.280 ;
        RECT 1213.670 3.670 1221.570 4.280 ;
        RECT 1222.410 3.670 1230.310 4.280 ;
        RECT 1231.150 3.670 1239.050 4.280 ;
        RECT 1239.890 3.670 1247.790 4.280 ;
        RECT 1248.630 3.670 1256.530 4.280 ;
        RECT 1257.370 3.670 1265.270 4.280 ;
        RECT 1266.110 3.670 1274.010 4.280 ;
        RECT 1274.850 3.670 1282.750 4.280 ;
        RECT 1283.590 3.670 1291.490 4.280 ;
        RECT 1292.330 3.670 1300.230 4.280 ;
        RECT 1301.070 3.670 1308.970 4.280 ;
        RECT 1309.810 3.670 1317.710 4.280 ;
        RECT 1318.550 3.670 1326.450 4.280 ;
        RECT 1327.290 3.670 1335.190 4.280 ;
        RECT 1336.030 3.670 1343.930 4.280 ;
        RECT 1344.770 3.670 1352.670 4.280 ;
        RECT 1353.510 3.670 1361.410 4.280 ;
        RECT 1362.250 3.670 1370.150 4.280 ;
        RECT 1370.990 3.670 1378.890 4.280 ;
        RECT 1379.730 3.670 1387.630 4.280 ;
        RECT 1388.470 3.670 1396.370 4.280 ;
        RECT 1397.210 3.670 1405.110 4.280 ;
        RECT 1405.950 3.670 1413.850 4.280 ;
        RECT 1414.690 3.670 1422.590 4.280 ;
        RECT 1423.430 3.670 1431.330 4.280 ;
        RECT 1432.170 3.670 1440.070 4.280 ;
        RECT 1440.910 3.670 1448.810 4.280 ;
        RECT 1449.650 3.670 1457.550 4.280 ;
        RECT 1458.390 3.670 1466.290 4.280 ;
        RECT 1467.130 3.670 1475.030 4.280 ;
        RECT 1475.870 3.670 1483.770 4.280 ;
        RECT 1484.610 3.670 1492.510 4.280 ;
        RECT 1493.350 3.670 1501.250 4.280 ;
        RECT 1502.090 3.670 1509.990 4.280 ;
        RECT 1510.830 3.670 1518.730 4.280 ;
        RECT 1519.570 3.670 1527.470 4.280 ;
        RECT 1528.310 3.670 1536.210 4.280 ;
        RECT 1537.050 3.670 1544.950 4.280 ;
        RECT 1545.790 3.670 1553.690 4.280 ;
        RECT 1554.530 3.670 1562.430 4.280 ;
        RECT 1563.270 3.670 1571.170 4.280 ;
        RECT 1572.010 3.670 1579.910 4.280 ;
        RECT 1580.750 3.670 1588.650 4.280 ;
        RECT 1589.490 3.670 1597.390 4.280 ;
        RECT 1598.230 3.670 1606.130 4.280 ;
        RECT 1606.970 3.670 1614.870 4.280 ;
        RECT 1615.710 3.670 1623.610 4.280 ;
        RECT 1624.450 3.670 1632.350 4.280 ;
        RECT 1633.190 3.670 1641.090 4.280 ;
        RECT 1641.930 3.670 1649.830 4.280 ;
        RECT 1650.670 3.670 1658.570 4.280 ;
        RECT 1659.410 3.670 1667.310 4.280 ;
        RECT 1668.150 3.670 1676.050 4.280 ;
        RECT 1676.890 3.670 1684.790 4.280 ;
        RECT 1685.630 3.670 1693.530 4.280 ;
        RECT 1694.370 3.670 1702.270 4.280 ;
        RECT 1703.110 3.670 1711.010 4.280 ;
        RECT 1711.850 3.670 1719.750 4.280 ;
        RECT 1720.590 3.670 1728.490 4.280 ;
        RECT 1729.330 3.670 1737.230 4.280 ;
        RECT 1738.070 3.670 1745.970 4.280 ;
        RECT 1746.810 3.670 1754.710 4.280 ;
        RECT 1755.550 3.670 1763.450 4.280 ;
        RECT 1764.290 3.670 1772.190 4.280 ;
        RECT 1773.030 3.670 1780.930 4.280 ;
        RECT 1781.770 3.670 1789.670 4.280 ;
        RECT 1790.510 3.670 1798.410 4.280 ;
        RECT 1799.250 3.670 1807.150 4.280 ;
        RECT 1807.990 3.670 1815.890 4.280 ;
        RECT 1816.730 3.670 1824.630 4.280 ;
        RECT 1825.470 3.670 1833.370 4.280 ;
        RECT 1834.210 3.670 1842.110 4.280 ;
        RECT 1842.950 3.670 1850.850 4.280 ;
        RECT 1851.690 3.670 1859.590 4.280 ;
        RECT 1860.430 3.670 1868.330 4.280 ;
        RECT 1869.170 3.670 1877.070 4.280 ;
        RECT 1877.910 3.670 1885.810 4.280 ;
        RECT 1886.650 3.670 1894.550 4.280 ;
        RECT 1895.390 3.670 1903.290 4.280 ;
        RECT 1904.130 3.670 1912.030 4.280 ;
        RECT 1912.870 3.670 1920.770 4.280 ;
        RECT 1921.610 3.670 1929.510 4.280 ;
        RECT 1930.350 3.670 1938.250 4.280 ;
        RECT 1939.090 3.670 1946.990 4.280 ;
        RECT 1947.830 3.670 1955.730 4.280 ;
        RECT 1956.570 3.670 1964.470 4.280 ;
        RECT 1965.310 3.670 1973.210 4.280 ;
        RECT 1974.050 3.670 1981.950 4.280 ;
        RECT 1982.790 3.670 1990.690 4.280 ;
        RECT 1991.530 3.670 1999.430 4.280 ;
        RECT 2000.270 3.670 2008.170 4.280 ;
        RECT 2009.010 3.670 2016.910 4.280 ;
        RECT 2017.750 3.670 2025.650 4.280 ;
        RECT 2026.490 3.670 2034.390 4.280 ;
        RECT 2035.230 3.670 2043.130 4.280 ;
        RECT 2043.970 3.670 2051.870 4.280 ;
        RECT 2052.710 3.670 2060.610 4.280 ;
        RECT 2061.450 3.670 2069.350 4.280 ;
        RECT 2070.190 3.670 2078.090 4.280 ;
        RECT 2078.930 3.670 2086.830 4.280 ;
        RECT 2087.670 3.670 2095.570 4.280 ;
        RECT 2096.410 3.670 2104.310 4.280 ;
        RECT 2105.150 3.670 2113.050 4.280 ;
        RECT 2113.890 3.670 2121.790 4.280 ;
        RECT 2122.630 3.670 2130.530 4.280 ;
        RECT 2131.370 3.670 2139.270 4.280 ;
        RECT 2140.110 3.670 2148.010 4.280 ;
        RECT 2148.850 3.670 2156.750 4.280 ;
        RECT 2157.590 3.670 2197.320 4.280 ;
      LAYER met3 ;
        RECT 4.000 644.320 2196.000 649.905 ;
        RECT 4.400 642.920 2196.000 644.320 ;
        RECT 4.000 641.600 2196.000 642.920 ;
        RECT 4.400 640.200 2196.000 641.600 ;
        RECT 4.000 638.880 2196.000 640.200 ;
        RECT 4.400 637.480 2196.000 638.880 ;
        RECT 4.000 636.160 2196.000 637.480 ;
        RECT 4.400 634.760 2196.000 636.160 ;
        RECT 4.000 633.440 2196.000 634.760 ;
        RECT 4.400 632.040 2196.000 633.440 ;
        RECT 4.000 630.720 2196.000 632.040 ;
        RECT 4.400 629.320 2196.000 630.720 ;
        RECT 4.000 628.000 2196.000 629.320 ;
        RECT 4.400 626.600 2196.000 628.000 ;
        RECT 4.000 625.280 2196.000 626.600 ;
        RECT 4.400 623.880 2196.000 625.280 ;
        RECT 4.000 622.560 2196.000 623.880 ;
        RECT 4.400 621.160 2196.000 622.560 ;
        RECT 4.000 619.840 2196.000 621.160 ;
        RECT 4.400 618.440 2196.000 619.840 ;
        RECT 4.000 617.120 2196.000 618.440 ;
        RECT 4.400 615.720 2196.000 617.120 ;
        RECT 4.000 614.400 2196.000 615.720 ;
        RECT 4.400 613.000 2196.000 614.400 ;
        RECT 4.000 611.680 2196.000 613.000 ;
        RECT 4.400 610.280 2196.000 611.680 ;
        RECT 4.000 608.960 2196.000 610.280 ;
        RECT 4.400 607.560 2196.000 608.960 ;
        RECT 4.000 606.240 2196.000 607.560 ;
        RECT 4.400 604.840 2196.000 606.240 ;
        RECT 4.000 603.520 2196.000 604.840 ;
        RECT 4.400 602.120 2196.000 603.520 ;
        RECT 4.000 600.800 2196.000 602.120 ;
        RECT 4.400 599.400 2196.000 600.800 ;
        RECT 4.000 598.080 2196.000 599.400 ;
        RECT 4.400 596.680 2196.000 598.080 ;
        RECT 4.000 595.360 2196.000 596.680 ;
        RECT 4.400 593.960 2196.000 595.360 ;
        RECT 4.000 592.640 2196.000 593.960 ;
        RECT 4.400 591.240 2196.000 592.640 ;
        RECT 4.000 589.920 2196.000 591.240 ;
        RECT 4.400 588.520 2196.000 589.920 ;
        RECT 4.000 587.200 2196.000 588.520 ;
        RECT 4.400 585.800 2196.000 587.200 ;
        RECT 4.000 584.480 2196.000 585.800 ;
        RECT 4.400 583.080 2196.000 584.480 ;
        RECT 4.000 581.760 2196.000 583.080 ;
        RECT 4.400 580.360 2196.000 581.760 ;
        RECT 4.000 579.040 2196.000 580.360 ;
        RECT 4.400 577.640 2196.000 579.040 ;
        RECT 4.000 576.320 2196.000 577.640 ;
        RECT 4.400 574.920 2196.000 576.320 ;
        RECT 4.000 573.600 2196.000 574.920 ;
        RECT 4.400 572.200 2196.000 573.600 ;
        RECT 4.000 570.880 2196.000 572.200 ;
        RECT 4.400 569.480 2196.000 570.880 ;
        RECT 4.000 568.160 2196.000 569.480 ;
        RECT 4.400 566.760 2196.000 568.160 ;
        RECT 4.000 565.440 2196.000 566.760 ;
        RECT 4.400 564.040 2196.000 565.440 ;
        RECT 4.000 562.720 2196.000 564.040 ;
        RECT 4.400 561.320 2196.000 562.720 ;
        RECT 4.000 560.000 2196.000 561.320 ;
        RECT 4.400 558.600 2196.000 560.000 ;
        RECT 4.000 557.280 2196.000 558.600 ;
        RECT 4.400 555.880 2196.000 557.280 ;
        RECT 4.000 554.560 2196.000 555.880 ;
        RECT 4.400 553.160 2196.000 554.560 ;
        RECT 4.000 551.840 2196.000 553.160 ;
        RECT 4.400 550.440 2196.000 551.840 ;
        RECT 4.000 549.120 2196.000 550.440 ;
        RECT 4.400 547.720 2196.000 549.120 ;
        RECT 4.000 546.400 2196.000 547.720 ;
        RECT 4.400 545.000 2196.000 546.400 ;
        RECT 4.000 543.680 2196.000 545.000 ;
        RECT 4.400 542.280 2196.000 543.680 ;
        RECT 4.000 540.960 2196.000 542.280 ;
        RECT 4.400 539.560 2196.000 540.960 ;
        RECT 4.000 538.240 2196.000 539.560 ;
        RECT 4.400 536.840 2196.000 538.240 ;
        RECT 4.000 535.520 2196.000 536.840 ;
        RECT 4.400 534.120 2196.000 535.520 ;
        RECT 4.000 532.800 2196.000 534.120 ;
        RECT 4.400 531.400 2196.000 532.800 ;
        RECT 4.000 530.080 2196.000 531.400 ;
        RECT 4.400 528.680 2196.000 530.080 ;
        RECT 4.000 527.360 2196.000 528.680 ;
        RECT 4.400 525.960 2196.000 527.360 ;
        RECT 4.000 524.640 2196.000 525.960 ;
        RECT 4.400 523.240 2196.000 524.640 ;
        RECT 4.000 521.920 2196.000 523.240 ;
        RECT 4.400 520.520 2196.000 521.920 ;
        RECT 4.000 519.200 2196.000 520.520 ;
        RECT 4.400 517.800 2196.000 519.200 ;
        RECT 4.000 516.480 2196.000 517.800 ;
        RECT 4.400 515.080 2196.000 516.480 ;
        RECT 4.000 513.760 2196.000 515.080 ;
        RECT 4.400 512.360 2196.000 513.760 ;
        RECT 4.000 511.040 2196.000 512.360 ;
        RECT 4.400 509.640 2196.000 511.040 ;
        RECT 4.000 508.320 2196.000 509.640 ;
        RECT 4.400 506.920 2196.000 508.320 ;
        RECT 4.000 505.600 2196.000 506.920 ;
        RECT 4.400 504.200 2196.000 505.600 ;
        RECT 4.000 502.880 2196.000 504.200 ;
        RECT 4.400 501.480 2196.000 502.880 ;
        RECT 4.000 500.160 2196.000 501.480 ;
        RECT 4.400 498.760 2196.000 500.160 ;
        RECT 4.000 497.440 2196.000 498.760 ;
        RECT 4.400 496.040 2196.000 497.440 ;
        RECT 4.000 494.720 2196.000 496.040 ;
        RECT 4.400 493.320 2196.000 494.720 ;
        RECT 4.000 492.000 2196.000 493.320 ;
        RECT 4.400 490.600 2196.000 492.000 ;
        RECT 4.000 489.280 2196.000 490.600 ;
        RECT 4.400 487.920 2196.000 489.280 ;
        RECT 4.400 487.880 2195.600 487.920 ;
        RECT 4.000 486.560 2195.600 487.880 ;
        RECT 4.400 485.160 2195.600 486.560 ;
        RECT 4.000 483.840 2195.600 485.160 ;
        RECT 4.400 482.440 2195.600 483.840 ;
        RECT 4.000 481.120 2195.600 482.440 ;
        RECT 4.400 479.720 2195.600 481.120 ;
        RECT 4.000 478.400 2195.600 479.720 ;
        RECT 4.400 477.000 2195.600 478.400 ;
        RECT 4.000 475.680 2195.600 477.000 ;
        RECT 4.400 474.280 2195.600 475.680 ;
        RECT 4.000 472.960 2195.600 474.280 ;
        RECT 4.400 471.560 2195.600 472.960 ;
        RECT 4.000 470.240 2195.600 471.560 ;
        RECT 4.400 468.840 2195.600 470.240 ;
        RECT 4.000 467.520 2195.600 468.840 ;
        RECT 4.400 466.120 2195.600 467.520 ;
        RECT 4.000 464.800 2195.600 466.120 ;
        RECT 4.400 463.400 2195.600 464.800 ;
        RECT 4.000 462.080 2195.600 463.400 ;
        RECT 4.400 460.680 2195.600 462.080 ;
        RECT 4.000 459.360 2195.600 460.680 ;
        RECT 4.400 457.960 2195.600 459.360 ;
        RECT 4.000 456.640 2195.600 457.960 ;
        RECT 4.400 455.240 2195.600 456.640 ;
        RECT 4.000 453.920 2195.600 455.240 ;
        RECT 4.400 452.520 2195.600 453.920 ;
        RECT 4.000 451.200 2195.600 452.520 ;
        RECT 4.400 449.800 2195.600 451.200 ;
        RECT 4.000 448.480 2195.600 449.800 ;
        RECT 4.400 447.080 2195.600 448.480 ;
        RECT 4.000 445.760 2195.600 447.080 ;
        RECT 4.400 444.360 2195.600 445.760 ;
        RECT 4.000 443.040 2195.600 444.360 ;
        RECT 4.400 441.640 2195.600 443.040 ;
        RECT 4.000 440.320 2195.600 441.640 ;
        RECT 4.400 438.920 2195.600 440.320 ;
        RECT 4.000 437.600 2195.600 438.920 ;
        RECT 4.400 436.200 2195.600 437.600 ;
        RECT 4.000 434.880 2195.600 436.200 ;
        RECT 4.400 433.480 2195.600 434.880 ;
        RECT 4.000 432.160 2195.600 433.480 ;
        RECT 4.400 430.760 2195.600 432.160 ;
        RECT 4.000 429.440 2195.600 430.760 ;
        RECT 4.400 428.040 2195.600 429.440 ;
        RECT 4.000 426.720 2195.600 428.040 ;
        RECT 4.400 425.320 2195.600 426.720 ;
        RECT 4.000 424.000 2195.600 425.320 ;
        RECT 4.400 422.600 2195.600 424.000 ;
        RECT 4.000 421.280 2195.600 422.600 ;
        RECT 4.400 419.880 2195.600 421.280 ;
        RECT 4.000 418.560 2195.600 419.880 ;
        RECT 4.400 417.160 2195.600 418.560 ;
        RECT 4.000 415.840 2195.600 417.160 ;
        RECT 4.400 414.440 2195.600 415.840 ;
        RECT 4.000 413.120 2195.600 414.440 ;
        RECT 4.400 411.720 2195.600 413.120 ;
        RECT 4.000 410.400 2195.600 411.720 ;
        RECT 4.400 409.000 2195.600 410.400 ;
        RECT 4.000 407.680 2195.600 409.000 ;
        RECT 4.400 406.280 2195.600 407.680 ;
        RECT 4.000 404.960 2195.600 406.280 ;
        RECT 4.400 403.560 2195.600 404.960 ;
        RECT 4.000 402.240 2195.600 403.560 ;
        RECT 4.400 400.840 2195.600 402.240 ;
        RECT 4.000 399.520 2195.600 400.840 ;
        RECT 4.400 398.120 2195.600 399.520 ;
        RECT 4.000 396.800 2195.600 398.120 ;
        RECT 4.400 395.400 2195.600 396.800 ;
        RECT 4.000 394.080 2195.600 395.400 ;
        RECT 4.400 392.680 2195.600 394.080 ;
        RECT 4.000 391.360 2195.600 392.680 ;
        RECT 4.400 389.960 2195.600 391.360 ;
        RECT 4.000 388.640 2195.600 389.960 ;
        RECT 4.400 387.240 2195.600 388.640 ;
        RECT 4.000 385.920 2195.600 387.240 ;
        RECT 4.400 384.520 2195.600 385.920 ;
        RECT 4.000 383.200 2195.600 384.520 ;
        RECT 4.400 381.800 2195.600 383.200 ;
        RECT 4.000 380.480 2195.600 381.800 ;
        RECT 4.400 379.080 2195.600 380.480 ;
        RECT 4.000 377.760 2195.600 379.080 ;
        RECT 4.400 376.360 2195.600 377.760 ;
        RECT 4.000 375.040 2195.600 376.360 ;
        RECT 4.400 373.640 2195.600 375.040 ;
        RECT 4.000 372.320 2195.600 373.640 ;
        RECT 4.400 370.920 2195.600 372.320 ;
        RECT 4.000 369.600 2195.600 370.920 ;
        RECT 4.400 368.200 2195.600 369.600 ;
        RECT 4.000 366.880 2195.600 368.200 ;
        RECT 4.400 365.480 2195.600 366.880 ;
        RECT 4.000 364.160 2195.600 365.480 ;
        RECT 4.400 362.760 2195.600 364.160 ;
        RECT 4.000 361.440 2195.600 362.760 ;
        RECT 4.400 360.040 2195.600 361.440 ;
        RECT 4.000 358.720 2195.600 360.040 ;
        RECT 4.400 357.320 2195.600 358.720 ;
        RECT 4.000 356.000 2195.600 357.320 ;
        RECT 4.400 354.600 2195.600 356.000 ;
        RECT 4.000 353.280 2195.600 354.600 ;
        RECT 4.400 351.880 2195.600 353.280 ;
        RECT 4.000 350.560 2195.600 351.880 ;
        RECT 4.400 349.160 2195.600 350.560 ;
        RECT 4.000 347.840 2195.600 349.160 ;
        RECT 4.400 346.440 2195.600 347.840 ;
        RECT 4.000 345.120 2195.600 346.440 ;
        RECT 4.400 343.720 2195.600 345.120 ;
        RECT 4.000 342.400 2195.600 343.720 ;
        RECT 4.400 341.000 2195.600 342.400 ;
        RECT 4.000 339.680 2195.600 341.000 ;
        RECT 4.400 338.280 2195.600 339.680 ;
        RECT 4.000 336.960 2195.600 338.280 ;
        RECT 4.400 335.560 2195.600 336.960 ;
        RECT 4.000 334.240 2195.600 335.560 ;
        RECT 4.400 332.840 2195.600 334.240 ;
        RECT 4.000 331.520 2195.600 332.840 ;
        RECT 4.400 330.120 2195.600 331.520 ;
        RECT 4.000 328.800 2195.600 330.120 ;
        RECT 4.400 327.400 2195.600 328.800 ;
        RECT 4.000 326.080 2195.600 327.400 ;
        RECT 4.400 324.680 2195.600 326.080 ;
        RECT 4.000 323.360 2195.600 324.680 ;
        RECT 4.400 321.960 2195.600 323.360 ;
        RECT 4.000 320.640 2195.600 321.960 ;
        RECT 4.400 319.240 2195.600 320.640 ;
        RECT 4.000 317.920 2195.600 319.240 ;
        RECT 4.400 316.520 2195.600 317.920 ;
        RECT 4.000 315.200 2195.600 316.520 ;
        RECT 4.400 313.800 2195.600 315.200 ;
        RECT 4.000 312.480 2195.600 313.800 ;
        RECT 4.400 311.080 2195.600 312.480 ;
        RECT 4.000 309.760 2195.600 311.080 ;
        RECT 4.400 308.360 2195.600 309.760 ;
        RECT 4.000 307.040 2195.600 308.360 ;
        RECT 4.400 305.640 2195.600 307.040 ;
        RECT 4.000 304.320 2195.600 305.640 ;
        RECT 4.400 302.920 2195.600 304.320 ;
        RECT 4.000 301.600 2195.600 302.920 ;
        RECT 4.400 300.200 2195.600 301.600 ;
        RECT 4.000 298.880 2195.600 300.200 ;
        RECT 4.400 297.480 2195.600 298.880 ;
        RECT 4.000 296.160 2195.600 297.480 ;
        RECT 4.400 294.760 2195.600 296.160 ;
        RECT 4.000 293.440 2195.600 294.760 ;
        RECT 4.400 292.040 2195.600 293.440 ;
        RECT 4.000 290.720 2195.600 292.040 ;
        RECT 4.400 289.320 2195.600 290.720 ;
        RECT 4.000 288.000 2195.600 289.320 ;
        RECT 4.400 286.600 2195.600 288.000 ;
        RECT 4.000 285.280 2195.600 286.600 ;
        RECT 4.400 283.880 2195.600 285.280 ;
        RECT 4.000 282.560 2195.600 283.880 ;
        RECT 4.400 281.160 2195.600 282.560 ;
        RECT 4.000 279.840 2195.600 281.160 ;
        RECT 4.400 278.440 2195.600 279.840 ;
        RECT 4.000 277.120 2195.600 278.440 ;
        RECT 4.400 275.720 2195.600 277.120 ;
        RECT 4.000 274.400 2195.600 275.720 ;
        RECT 4.400 273.000 2195.600 274.400 ;
        RECT 4.000 271.680 2195.600 273.000 ;
        RECT 4.400 270.280 2195.600 271.680 ;
        RECT 4.000 268.960 2195.600 270.280 ;
        RECT 4.400 267.560 2195.600 268.960 ;
        RECT 4.000 266.240 2195.600 267.560 ;
        RECT 4.400 264.840 2195.600 266.240 ;
        RECT 4.000 263.520 2195.600 264.840 ;
        RECT 4.400 262.120 2195.600 263.520 ;
        RECT 4.000 260.800 2195.600 262.120 ;
        RECT 4.400 259.400 2195.600 260.800 ;
        RECT 4.000 258.080 2195.600 259.400 ;
        RECT 4.400 256.680 2195.600 258.080 ;
        RECT 4.000 255.360 2195.600 256.680 ;
        RECT 4.400 253.960 2195.600 255.360 ;
        RECT 4.000 252.640 2195.600 253.960 ;
        RECT 4.400 251.240 2195.600 252.640 ;
        RECT 4.000 249.920 2195.600 251.240 ;
        RECT 4.400 248.520 2195.600 249.920 ;
        RECT 4.000 247.200 2195.600 248.520 ;
        RECT 4.400 245.800 2195.600 247.200 ;
        RECT 4.000 244.480 2195.600 245.800 ;
        RECT 4.400 243.080 2195.600 244.480 ;
        RECT 4.000 241.760 2195.600 243.080 ;
        RECT 4.400 240.360 2195.600 241.760 ;
        RECT 4.000 239.040 2195.600 240.360 ;
        RECT 4.400 237.640 2195.600 239.040 ;
        RECT 4.000 236.320 2195.600 237.640 ;
        RECT 4.400 234.920 2195.600 236.320 ;
        RECT 4.000 233.600 2195.600 234.920 ;
        RECT 4.400 232.200 2195.600 233.600 ;
        RECT 4.000 230.880 2195.600 232.200 ;
        RECT 4.400 229.480 2195.600 230.880 ;
        RECT 4.000 228.160 2195.600 229.480 ;
        RECT 4.400 226.760 2195.600 228.160 ;
        RECT 4.000 225.440 2195.600 226.760 ;
        RECT 4.400 224.040 2195.600 225.440 ;
        RECT 4.000 222.720 2195.600 224.040 ;
        RECT 4.400 221.320 2195.600 222.720 ;
        RECT 4.000 220.000 2195.600 221.320 ;
        RECT 4.400 218.600 2195.600 220.000 ;
        RECT 4.000 217.280 2195.600 218.600 ;
        RECT 4.400 215.880 2195.600 217.280 ;
        RECT 4.000 214.560 2195.600 215.880 ;
        RECT 4.400 213.160 2195.600 214.560 ;
        RECT 4.000 211.840 2195.600 213.160 ;
        RECT 4.400 210.440 2195.600 211.840 ;
        RECT 4.000 209.120 2195.600 210.440 ;
        RECT 4.400 207.720 2195.600 209.120 ;
        RECT 4.000 206.400 2195.600 207.720 ;
        RECT 4.400 205.000 2195.600 206.400 ;
        RECT 4.000 203.680 2195.600 205.000 ;
        RECT 4.400 202.280 2195.600 203.680 ;
        RECT 4.000 200.960 2195.600 202.280 ;
        RECT 4.400 199.560 2195.600 200.960 ;
        RECT 4.000 198.240 2195.600 199.560 ;
        RECT 4.400 196.840 2195.600 198.240 ;
        RECT 4.000 195.520 2195.600 196.840 ;
        RECT 4.400 194.120 2195.600 195.520 ;
        RECT 4.000 192.800 2195.600 194.120 ;
        RECT 4.400 191.400 2195.600 192.800 ;
        RECT 4.000 190.080 2195.600 191.400 ;
        RECT 4.400 188.680 2195.600 190.080 ;
        RECT 4.000 187.360 2195.600 188.680 ;
        RECT 4.400 185.960 2195.600 187.360 ;
        RECT 4.000 184.640 2195.600 185.960 ;
        RECT 4.400 183.240 2195.600 184.640 ;
        RECT 4.000 181.920 2195.600 183.240 ;
        RECT 4.400 180.520 2195.600 181.920 ;
        RECT 4.000 179.200 2195.600 180.520 ;
        RECT 4.400 177.800 2195.600 179.200 ;
        RECT 4.000 176.480 2195.600 177.800 ;
        RECT 4.400 175.080 2195.600 176.480 ;
        RECT 4.000 173.760 2195.600 175.080 ;
        RECT 4.400 172.360 2195.600 173.760 ;
        RECT 4.000 171.040 2195.600 172.360 ;
        RECT 4.400 169.640 2195.600 171.040 ;
        RECT 4.000 168.320 2195.600 169.640 ;
        RECT 4.400 166.920 2195.600 168.320 ;
        RECT 4.000 165.600 2195.600 166.920 ;
        RECT 4.400 164.200 2195.600 165.600 ;
        RECT 4.000 162.880 2195.600 164.200 ;
        RECT 4.400 161.480 2195.600 162.880 ;
        RECT 4.000 160.160 2196.000 161.480 ;
        RECT 4.400 158.760 2196.000 160.160 ;
        RECT 4.000 157.440 2196.000 158.760 ;
        RECT 4.400 156.040 2196.000 157.440 ;
        RECT 4.000 154.720 2196.000 156.040 ;
        RECT 4.400 153.320 2196.000 154.720 ;
        RECT 4.000 152.000 2196.000 153.320 ;
        RECT 4.400 150.600 2196.000 152.000 ;
        RECT 4.000 149.280 2196.000 150.600 ;
        RECT 4.400 147.880 2196.000 149.280 ;
        RECT 4.000 146.560 2196.000 147.880 ;
        RECT 4.400 145.160 2196.000 146.560 ;
        RECT 4.000 143.840 2196.000 145.160 ;
        RECT 4.400 142.440 2196.000 143.840 ;
        RECT 4.000 141.120 2196.000 142.440 ;
        RECT 4.400 139.720 2196.000 141.120 ;
        RECT 4.000 138.400 2196.000 139.720 ;
        RECT 4.400 137.000 2196.000 138.400 ;
        RECT 4.000 135.680 2196.000 137.000 ;
        RECT 4.400 134.280 2196.000 135.680 ;
        RECT 4.000 132.960 2196.000 134.280 ;
        RECT 4.400 131.560 2196.000 132.960 ;
        RECT 4.000 130.240 2196.000 131.560 ;
        RECT 4.400 128.840 2196.000 130.240 ;
        RECT 4.000 127.520 2196.000 128.840 ;
        RECT 4.400 126.120 2196.000 127.520 ;
        RECT 4.000 124.800 2196.000 126.120 ;
        RECT 4.400 123.400 2196.000 124.800 ;
        RECT 4.000 122.080 2196.000 123.400 ;
        RECT 4.400 120.680 2196.000 122.080 ;
        RECT 4.000 119.360 2196.000 120.680 ;
        RECT 4.400 117.960 2196.000 119.360 ;
        RECT 4.000 116.640 2196.000 117.960 ;
        RECT 4.400 115.240 2196.000 116.640 ;
        RECT 4.000 113.920 2196.000 115.240 ;
        RECT 4.400 112.520 2196.000 113.920 ;
        RECT 4.000 111.200 2196.000 112.520 ;
        RECT 4.400 109.800 2196.000 111.200 ;
        RECT 4.000 108.480 2196.000 109.800 ;
        RECT 4.400 107.080 2196.000 108.480 ;
        RECT 4.000 105.760 2196.000 107.080 ;
        RECT 4.400 104.360 2196.000 105.760 ;
        RECT 4.000 103.040 2196.000 104.360 ;
        RECT 4.400 101.640 2196.000 103.040 ;
        RECT 4.000 100.320 2196.000 101.640 ;
        RECT 4.400 98.920 2196.000 100.320 ;
        RECT 4.000 97.600 2196.000 98.920 ;
        RECT 4.400 96.200 2196.000 97.600 ;
        RECT 4.000 94.880 2196.000 96.200 ;
        RECT 4.400 93.480 2196.000 94.880 ;
        RECT 4.000 92.160 2196.000 93.480 ;
        RECT 4.400 90.760 2196.000 92.160 ;
        RECT 4.000 89.440 2196.000 90.760 ;
        RECT 4.400 88.040 2196.000 89.440 ;
        RECT 4.000 86.720 2196.000 88.040 ;
        RECT 4.400 85.320 2196.000 86.720 ;
        RECT 4.000 84.000 2196.000 85.320 ;
        RECT 4.400 82.600 2196.000 84.000 ;
        RECT 4.000 81.280 2196.000 82.600 ;
        RECT 4.400 79.880 2196.000 81.280 ;
        RECT 4.000 78.560 2196.000 79.880 ;
        RECT 4.400 77.160 2196.000 78.560 ;
        RECT 4.000 75.840 2196.000 77.160 ;
        RECT 4.400 74.440 2196.000 75.840 ;
        RECT 4.000 73.120 2196.000 74.440 ;
        RECT 4.400 71.720 2196.000 73.120 ;
        RECT 4.000 70.400 2196.000 71.720 ;
        RECT 4.400 69.000 2196.000 70.400 ;
        RECT 4.000 67.680 2196.000 69.000 ;
        RECT 4.400 66.280 2196.000 67.680 ;
        RECT 4.000 64.960 2196.000 66.280 ;
        RECT 4.400 63.560 2196.000 64.960 ;
        RECT 4.000 62.240 2196.000 63.560 ;
        RECT 4.400 60.840 2196.000 62.240 ;
        RECT 4.000 59.520 2196.000 60.840 ;
        RECT 4.400 58.120 2196.000 59.520 ;
        RECT 4.000 56.800 2196.000 58.120 ;
        RECT 4.400 55.400 2196.000 56.800 ;
        RECT 4.000 54.080 2196.000 55.400 ;
        RECT 4.400 52.680 2196.000 54.080 ;
        RECT 4.000 51.360 2196.000 52.680 ;
        RECT 4.400 49.960 2196.000 51.360 ;
        RECT 4.000 48.640 2196.000 49.960 ;
        RECT 4.400 47.240 2196.000 48.640 ;
        RECT 4.000 45.920 2196.000 47.240 ;
        RECT 4.400 44.520 2196.000 45.920 ;
        RECT 4.000 43.200 2196.000 44.520 ;
        RECT 4.400 41.800 2196.000 43.200 ;
        RECT 4.000 40.480 2196.000 41.800 ;
        RECT 4.400 39.080 2196.000 40.480 ;
        RECT 4.000 37.760 2196.000 39.080 ;
        RECT 4.400 36.360 2196.000 37.760 ;
        RECT 4.000 35.040 2196.000 36.360 ;
        RECT 4.400 33.640 2196.000 35.040 ;
        RECT 4.000 32.320 2196.000 33.640 ;
        RECT 4.400 30.920 2196.000 32.320 ;
        RECT 4.000 29.600 2196.000 30.920 ;
        RECT 4.400 28.200 2196.000 29.600 ;
        RECT 4.000 26.880 2196.000 28.200 ;
        RECT 4.400 25.480 2196.000 26.880 ;
        RECT 4.000 24.160 2196.000 25.480 ;
        RECT 4.400 22.760 2196.000 24.160 ;
        RECT 4.000 21.440 2196.000 22.760 ;
        RECT 4.400 20.040 2196.000 21.440 ;
        RECT 4.000 18.720 2196.000 20.040 ;
        RECT 4.400 17.320 2196.000 18.720 ;
        RECT 4.000 16.000 2196.000 17.320 ;
        RECT 4.400 14.600 2196.000 16.000 ;
        RECT 4.000 13.280 2196.000 14.600 ;
        RECT 4.400 11.880 2196.000 13.280 ;
        RECT 4.000 10.560 2196.000 11.880 ;
        RECT 4.400 9.160 2196.000 10.560 ;
        RECT 4.000 7.840 2196.000 9.160 ;
        RECT 4.400 6.440 2196.000 7.840 ;
        RECT 4.000 5.120 2196.000 6.440 ;
        RECT 4.400 4.260 2196.000 5.120 ;
      LAYER met4 ;
        RECT 704.095 637.120 2180.105 649.905 ;
        RECT 704.095 10.240 711.840 637.120 ;
        RECT 714.240 10.240 788.640 637.120 ;
        RECT 791.040 10.240 865.440 637.120 ;
        RECT 867.840 10.240 942.240 637.120 ;
        RECT 944.640 10.240 1019.040 637.120 ;
        RECT 1021.440 10.240 1095.840 637.120 ;
        RECT 1098.240 10.240 1172.640 637.120 ;
        RECT 1175.040 10.240 1249.440 637.120 ;
        RECT 1251.840 10.240 1326.240 637.120 ;
        RECT 1328.640 10.240 1403.040 637.120 ;
        RECT 1405.440 10.240 1479.840 637.120 ;
        RECT 1482.240 10.240 1556.640 637.120 ;
        RECT 1559.040 10.240 1633.440 637.120 ;
        RECT 1635.840 10.240 1710.240 637.120 ;
        RECT 1712.640 10.240 1787.040 637.120 ;
        RECT 1789.440 10.240 1863.840 637.120 ;
        RECT 1866.240 10.240 1940.640 637.120 ;
        RECT 1943.040 10.240 2017.440 637.120 ;
        RECT 2019.840 10.240 2094.240 637.120 ;
        RECT 2096.640 10.240 2171.040 637.120 ;
        RECT 2173.440 10.240 2180.105 637.120 ;
        RECT 704.095 4.255 2180.105 10.240 ;
  END
END vliw
END LIBRARY

