magic
tech sky130B
magscale 1 2
timestamp 1716985692
<< obsli1 >>
rect 1104 2159 38824 197489
<< obsm1 >>
rect 14 2128 39914 197520
<< metal2 >>
rect 754 199200 810 200000
rect 1766 199200 1822 200000
rect 2778 199200 2834 200000
rect 3790 199200 3846 200000
rect 4802 199200 4858 200000
rect 5814 199200 5870 200000
rect 6826 199200 6882 200000
rect 7838 199200 7894 200000
rect 8850 199200 8906 200000
rect 9862 199200 9918 200000
rect 10874 199200 10930 200000
rect 11886 199200 11942 200000
rect 12898 199200 12954 200000
rect 13910 199200 13966 200000
rect 14922 199200 14978 200000
rect 15934 199200 15990 200000
rect 16946 199200 17002 200000
rect 17958 199200 18014 200000
rect 18970 199200 19026 200000
rect 19982 199200 20038 200000
rect 20994 199200 21050 200000
rect 22006 199200 22062 200000
rect 23018 199200 23074 200000
rect 24030 199200 24086 200000
rect 25042 199200 25098 200000
rect 26054 199200 26110 200000
rect 27066 199200 27122 200000
rect 28078 199200 28134 200000
rect 29090 199200 29146 200000
rect 30102 199200 30158 200000
rect 31114 199200 31170 200000
rect 32126 199200 32182 200000
rect 33138 199200 33194 200000
rect 34150 199200 34206 200000
rect 35162 199200 35218 200000
rect 36174 199200 36230 200000
rect 37186 199200 37242 200000
rect 38198 199200 38254 200000
rect 39210 199200 39266 200000
rect 1398 0 1454 800
rect 2594 0 2650 800
rect 3790 0 3846 800
rect 4986 0 5042 800
rect 6182 0 6238 800
rect 7378 0 7434 800
rect 8574 0 8630 800
rect 9770 0 9826 800
rect 10966 0 11022 800
rect 12162 0 12218 800
rect 13358 0 13414 800
rect 14554 0 14610 800
rect 15750 0 15806 800
rect 16946 0 17002 800
rect 18142 0 18198 800
rect 19338 0 19394 800
rect 20534 0 20590 800
rect 21730 0 21786 800
rect 22926 0 22982 800
rect 24122 0 24178 800
rect 25318 0 25374 800
rect 26514 0 26570 800
rect 27710 0 27766 800
rect 28906 0 28962 800
rect 30102 0 30158 800
rect 31298 0 31354 800
rect 32494 0 32550 800
rect 33690 0 33746 800
rect 34886 0 34942 800
rect 36082 0 36138 800
rect 37278 0 37334 800
rect 38474 0 38530 800
<< obsm2 >>
rect 20 199144 698 199322
rect 866 199144 1710 199322
rect 1878 199144 2722 199322
rect 2890 199144 3734 199322
rect 3902 199144 4746 199322
rect 4914 199144 5758 199322
rect 5926 199144 6770 199322
rect 6938 199144 7782 199322
rect 7950 199144 8794 199322
rect 8962 199144 9806 199322
rect 9974 199144 10818 199322
rect 10986 199144 11830 199322
rect 11998 199144 12842 199322
rect 13010 199144 13854 199322
rect 14022 199144 14866 199322
rect 15034 199144 15878 199322
rect 16046 199144 16890 199322
rect 17058 199144 17902 199322
rect 18070 199144 18914 199322
rect 19082 199144 19926 199322
rect 20094 199144 20938 199322
rect 21106 199144 21950 199322
rect 22118 199144 22962 199322
rect 23130 199144 23974 199322
rect 24142 199144 24986 199322
rect 25154 199144 25998 199322
rect 26166 199144 27010 199322
rect 27178 199144 28022 199322
rect 28190 199144 29034 199322
rect 29202 199144 30046 199322
rect 30214 199144 31058 199322
rect 31226 199144 32070 199322
rect 32238 199144 33082 199322
rect 33250 199144 34094 199322
rect 34262 199144 35106 199322
rect 35274 199144 36118 199322
rect 36286 199144 37130 199322
rect 37298 199144 38142 199322
rect 38310 199144 39154 199322
rect 39322 199144 39988 199322
rect 20 856 39988 199144
rect 20 800 1342 856
rect 1510 800 2538 856
rect 2706 800 3734 856
rect 3902 800 4930 856
rect 5098 800 6126 856
rect 6294 800 7322 856
rect 7490 800 8518 856
rect 8686 800 9714 856
rect 9882 800 10910 856
rect 11078 800 12106 856
rect 12274 800 13302 856
rect 13470 800 14498 856
rect 14666 800 15694 856
rect 15862 800 16890 856
rect 17058 800 18086 856
rect 18254 800 19282 856
rect 19450 800 20478 856
rect 20646 800 21674 856
rect 21842 800 22870 856
rect 23038 800 24066 856
rect 24234 800 25262 856
rect 25430 800 26458 856
rect 26626 800 27654 856
rect 27822 800 28850 856
rect 29018 800 30046 856
rect 30214 800 31242 856
rect 31410 800 32438 856
rect 32606 800 33634 856
rect 33802 800 34830 856
rect 34998 800 36026 856
rect 36194 800 37222 856
rect 37390 800 38418 856
rect 38586 800 39988 856
<< metal3 >>
rect 39200 198296 40000 198416
rect 39200 196936 40000 197056
rect 39200 195576 40000 195696
rect 39200 194216 40000 194336
rect 39200 192856 40000 192976
rect 39200 191496 40000 191616
rect 39200 190136 40000 190256
rect 39200 188776 40000 188896
rect 39200 187416 40000 187536
rect 39200 186056 40000 186176
rect 39200 184696 40000 184816
rect 39200 183336 40000 183456
rect 39200 181976 40000 182096
rect 39200 180616 40000 180736
rect 39200 179256 40000 179376
rect 39200 177896 40000 178016
rect 39200 176536 40000 176656
rect 39200 175176 40000 175296
rect 39200 173816 40000 173936
rect 39200 172456 40000 172576
rect 39200 171096 40000 171216
rect 39200 169736 40000 169856
rect 0 168376 800 168496
rect 39200 168376 40000 168496
rect 0 167832 800 167952
rect 0 167288 800 167408
rect 39200 167016 40000 167136
rect 0 166744 800 166864
rect 0 166200 800 166320
rect 0 165656 800 165776
rect 39200 165656 40000 165776
rect 0 165112 800 165232
rect 0 164568 800 164688
rect 39200 164296 40000 164416
rect 0 164024 800 164144
rect 0 163480 800 163600
rect 0 162936 800 163056
rect 39200 162936 40000 163056
rect 0 162392 800 162512
rect 0 161848 800 161968
rect 39200 161576 40000 161696
rect 0 161304 800 161424
rect 0 160760 800 160880
rect 0 160216 800 160336
rect 39200 160216 40000 160336
rect 0 159672 800 159792
rect 0 159128 800 159248
rect 39200 158856 40000 158976
rect 0 158584 800 158704
rect 0 158040 800 158160
rect 0 157496 800 157616
rect 39200 157496 40000 157616
rect 0 156952 800 157072
rect 0 156408 800 156528
rect 39200 156136 40000 156256
rect 0 155864 800 155984
rect 0 155320 800 155440
rect 0 154776 800 154896
rect 39200 154776 40000 154896
rect 0 154232 800 154352
rect 0 153688 800 153808
rect 39200 153416 40000 153536
rect 0 153144 800 153264
rect 0 152600 800 152720
rect 0 152056 800 152176
rect 39200 152056 40000 152176
rect 0 151512 800 151632
rect 0 150968 800 151088
rect 39200 150696 40000 150816
rect 0 150424 800 150544
rect 0 149880 800 150000
rect 0 149336 800 149456
rect 39200 149336 40000 149456
rect 0 148792 800 148912
rect 0 148248 800 148368
rect 39200 147976 40000 148096
rect 0 147704 800 147824
rect 0 147160 800 147280
rect 0 146616 800 146736
rect 39200 146616 40000 146736
rect 0 146072 800 146192
rect 0 145528 800 145648
rect 39200 145256 40000 145376
rect 0 144984 800 145104
rect 0 144440 800 144560
rect 0 143896 800 144016
rect 39200 143896 40000 144016
rect 0 143352 800 143472
rect 0 142808 800 142928
rect 39200 142536 40000 142656
rect 0 142264 800 142384
rect 0 141720 800 141840
rect 0 141176 800 141296
rect 39200 141176 40000 141296
rect 0 140632 800 140752
rect 0 140088 800 140208
rect 39200 139816 40000 139936
rect 0 139544 800 139664
rect 0 139000 800 139120
rect 0 138456 800 138576
rect 39200 138456 40000 138576
rect 0 137912 800 138032
rect 0 137368 800 137488
rect 39200 137096 40000 137216
rect 0 136824 800 136944
rect 0 136280 800 136400
rect 0 135736 800 135856
rect 39200 135736 40000 135856
rect 0 135192 800 135312
rect 0 134648 800 134768
rect 39200 134376 40000 134496
rect 0 134104 800 134224
rect 0 133560 800 133680
rect 0 133016 800 133136
rect 39200 133016 40000 133136
rect 0 132472 800 132592
rect 0 131928 800 132048
rect 39200 131656 40000 131776
rect 0 131384 800 131504
rect 0 130840 800 130960
rect 0 130296 800 130416
rect 39200 130296 40000 130416
rect 0 129752 800 129872
rect 0 129208 800 129328
rect 39200 128936 40000 129056
rect 0 128664 800 128784
rect 0 128120 800 128240
rect 0 127576 800 127696
rect 39200 127576 40000 127696
rect 0 127032 800 127152
rect 0 126488 800 126608
rect 39200 126216 40000 126336
rect 0 125944 800 126064
rect 0 125400 800 125520
rect 0 124856 800 124976
rect 39200 124856 40000 124976
rect 0 124312 800 124432
rect 0 123768 800 123888
rect 39200 123496 40000 123616
rect 0 123224 800 123344
rect 0 122680 800 122800
rect 0 122136 800 122256
rect 39200 122136 40000 122256
rect 0 121592 800 121712
rect 0 121048 800 121168
rect 39200 120776 40000 120896
rect 0 120504 800 120624
rect 0 119960 800 120080
rect 0 119416 800 119536
rect 39200 119416 40000 119536
rect 0 118872 800 118992
rect 0 118328 800 118448
rect 39200 118056 40000 118176
rect 0 117784 800 117904
rect 0 117240 800 117360
rect 0 116696 800 116816
rect 39200 116696 40000 116816
rect 0 116152 800 116272
rect 0 115608 800 115728
rect 39200 115336 40000 115456
rect 0 115064 800 115184
rect 0 114520 800 114640
rect 0 113976 800 114096
rect 39200 113976 40000 114096
rect 0 113432 800 113552
rect 0 112888 800 113008
rect 39200 112616 40000 112736
rect 0 112344 800 112464
rect 0 111800 800 111920
rect 0 111256 800 111376
rect 39200 111256 40000 111376
rect 0 110712 800 110832
rect 0 110168 800 110288
rect 39200 109896 40000 110016
rect 0 109624 800 109744
rect 0 109080 800 109200
rect 0 108536 800 108656
rect 39200 108536 40000 108656
rect 0 107992 800 108112
rect 0 107448 800 107568
rect 39200 107176 40000 107296
rect 0 106904 800 107024
rect 0 106360 800 106480
rect 0 105816 800 105936
rect 39200 105816 40000 105936
rect 0 105272 800 105392
rect 0 104728 800 104848
rect 39200 104456 40000 104576
rect 0 104184 800 104304
rect 0 103640 800 103760
rect 0 103096 800 103216
rect 39200 103096 40000 103216
rect 0 102552 800 102672
rect 0 102008 800 102128
rect 39200 101736 40000 101856
rect 0 101464 800 101584
rect 0 100920 800 101040
rect 0 100376 800 100496
rect 39200 100376 40000 100496
rect 0 99832 800 99952
rect 0 99288 800 99408
rect 39200 99016 40000 99136
rect 0 98744 800 98864
rect 0 98200 800 98320
rect 0 97656 800 97776
rect 39200 97656 40000 97776
rect 0 97112 800 97232
rect 0 96568 800 96688
rect 39200 96296 40000 96416
rect 0 96024 800 96144
rect 0 95480 800 95600
rect 0 94936 800 95056
rect 39200 94936 40000 95056
rect 0 94392 800 94512
rect 0 93848 800 93968
rect 39200 93576 40000 93696
rect 0 93304 800 93424
rect 0 92760 800 92880
rect 0 92216 800 92336
rect 39200 92216 40000 92336
rect 0 91672 800 91792
rect 0 91128 800 91248
rect 39200 90856 40000 90976
rect 0 90584 800 90704
rect 0 90040 800 90160
rect 0 89496 800 89616
rect 39200 89496 40000 89616
rect 0 88952 800 89072
rect 0 88408 800 88528
rect 39200 88136 40000 88256
rect 0 87864 800 87984
rect 0 87320 800 87440
rect 0 86776 800 86896
rect 39200 86776 40000 86896
rect 0 86232 800 86352
rect 0 85688 800 85808
rect 39200 85416 40000 85536
rect 0 85144 800 85264
rect 0 84600 800 84720
rect 0 84056 800 84176
rect 39200 84056 40000 84176
rect 0 83512 800 83632
rect 0 82968 800 83088
rect 39200 82696 40000 82816
rect 0 82424 800 82544
rect 0 81880 800 82000
rect 0 81336 800 81456
rect 39200 81336 40000 81456
rect 0 80792 800 80912
rect 0 80248 800 80368
rect 39200 79976 40000 80096
rect 0 79704 800 79824
rect 0 79160 800 79280
rect 0 78616 800 78736
rect 39200 78616 40000 78736
rect 0 78072 800 78192
rect 0 77528 800 77648
rect 39200 77256 40000 77376
rect 0 76984 800 77104
rect 0 76440 800 76560
rect 0 75896 800 76016
rect 39200 75896 40000 76016
rect 0 75352 800 75472
rect 0 74808 800 74928
rect 39200 74536 40000 74656
rect 0 74264 800 74384
rect 0 73720 800 73840
rect 0 73176 800 73296
rect 39200 73176 40000 73296
rect 0 72632 800 72752
rect 0 72088 800 72208
rect 39200 71816 40000 71936
rect 0 71544 800 71664
rect 0 71000 800 71120
rect 0 70456 800 70576
rect 39200 70456 40000 70576
rect 0 69912 800 70032
rect 0 69368 800 69488
rect 39200 69096 40000 69216
rect 0 68824 800 68944
rect 0 68280 800 68400
rect 0 67736 800 67856
rect 39200 67736 40000 67856
rect 0 67192 800 67312
rect 0 66648 800 66768
rect 39200 66376 40000 66496
rect 0 66104 800 66224
rect 0 65560 800 65680
rect 0 65016 800 65136
rect 39200 65016 40000 65136
rect 0 64472 800 64592
rect 0 63928 800 64048
rect 39200 63656 40000 63776
rect 0 63384 800 63504
rect 0 62840 800 62960
rect 0 62296 800 62416
rect 39200 62296 40000 62416
rect 0 61752 800 61872
rect 0 61208 800 61328
rect 39200 60936 40000 61056
rect 0 60664 800 60784
rect 0 60120 800 60240
rect 0 59576 800 59696
rect 39200 59576 40000 59696
rect 0 59032 800 59152
rect 0 58488 800 58608
rect 39200 58216 40000 58336
rect 0 57944 800 58064
rect 0 57400 800 57520
rect 0 56856 800 56976
rect 39200 56856 40000 56976
rect 0 56312 800 56432
rect 0 55768 800 55888
rect 39200 55496 40000 55616
rect 0 55224 800 55344
rect 0 54680 800 54800
rect 0 54136 800 54256
rect 39200 54136 40000 54256
rect 0 53592 800 53712
rect 0 53048 800 53168
rect 39200 52776 40000 52896
rect 0 52504 800 52624
rect 0 51960 800 52080
rect 0 51416 800 51536
rect 39200 51416 40000 51536
rect 0 50872 800 50992
rect 0 50328 800 50448
rect 39200 50056 40000 50176
rect 0 49784 800 49904
rect 0 49240 800 49360
rect 0 48696 800 48816
rect 39200 48696 40000 48816
rect 0 48152 800 48272
rect 0 47608 800 47728
rect 39200 47336 40000 47456
rect 0 47064 800 47184
rect 0 46520 800 46640
rect 0 45976 800 46096
rect 39200 45976 40000 46096
rect 0 45432 800 45552
rect 0 44888 800 45008
rect 39200 44616 40000 44736
rect 0 44344 800 44464
rect 0 43800 800 43920
rect 0 43256 800 43376
rect 39200 43256 40000 43376
rect 0 42712 800 42832
rect 0 42168 800 42288
rect 39200 41896 40000 42016
rect 0 41624 800 41744
rect 0 41080 800 41200
rect 0 40536 800 40656
rect 39200 40536 40000 40656
rect 0 39992 800 40112
rect 0 39448 800 39568
rect 39200 39176 40000 39296
rect 0 38904 800 39024
rect 0 38360 800 38480
rect 0 37816 800 37936
rect 39200 37816 40000 37936
rect 0 37272 800 37392
rect 0 36728 800 36848
rect 39200 36456 40000 36576
rect 0 36184 800 36304
rect 0 35640 800 35760
rect 0 35096 800 35216
rect 39200 35096 40000 35216
rect 0 34552 800 34672
rect 0 34008 800 34128
rect 39200 33736 40000 33856
rect 0 33464 800 33584
rect 0 32920 800 33040
rect 0 32376 800 32496
rect 39200 32376 40000 32496
rect 0 31832 800 31952
rect 0 31288 800 31408
rect 39200 31016 40000 31136
rect 39200 29656 40000 29776
rect 39200 28296 40000 28416
rect 39200 26936 40000 27056
rect 39200 25576 40000 25696
rect 39200 24216 40000 24336
rect 39200 22856 40000 22976
rect 39200 21496 40000 21616
rect 39200 20136 40000 20256
rect 39200 18776 40000 18896
rect 39200 17416 40000 17536
rect 39200 16056 40000 16176
rect 39200 14696 40000 14816
rect 39200 13336 40000 13456
rect 39200 11976 40000 12096
rect 39200 10616 40000 10736
rect 39200 9256 40000 9376
rect 39200 7896 40000 8016
rect 39200 6536 40000 6656
rect 39200 5176 40000 5296
rect 39200 3816 40000 3936
rect 39200 2456 40000 2576
rect 39200 1096 40000 1216
<< obsm3 >>
rect 381 198216 39120 198389
rect 381 197136 39200 198216
rect 381 196856 39120 197136
rect 381 195776 39200 196856
rect 381 195496 39120 195776
rect 381 194416 39200 195496
rect 381 194136 39120 194416
rect 381 193056 39200 194136
rect 381 192776 39120 193056
rect 381 191696 39200 192776
rect 381 191416 39120 191696
rect 381 190336 39200 191416
rect 381 190056 39120 190336
rect 381 188976 39200 190056
rect 381 188696 39120 188976
rect 381 187616 39200 188696
rect 381 187336 39120 187616
rect 381 186256 39200 187336
rect 381 185976 39120 186256
rect 381 184896 39200 185976
rect 381 184616 39120 184896
rect 381 183536 39200 184616
rect 381 183256 39120 183536
rect 381 182176 39200 183256
rect 381 181896 39120 182176
rect 381 180816 39200 181896
rect 381 180536 39120 180816
rect 381 179456 39200 180536
rect 381 179176 39120 179456
rect 381 178096 39200 179176
rect 381 177816 39120 178096
rect 381 176736 39200 177816
rect 381 176456 39120 176736
rect 381 175376 39200 176456
rect 381 175096 39120 175376
rect 381 174016 39200 175096
rect 381 173736 39120 174016
rect 381 172656 39200 173736
rect 381 172376 39120 172656
rect 381 171296 39200 172376
rect 381 171016 39120 171296
rect 381 169936 39200 171016
rect 381 169656 39120 169936
rect 381 168576 39200 169656
rect 880 168296 39120 168576
rect 381 168032 39200 168296
rect 880 167752 39200 168032
rect 381 167488 39200 167752
rect 880 167216 39200 167488
rect 880 167208 39120 167216
rect 381 166944 39120 167208
rect 880 166936 39120 166944
rect 880 166664 39200 166936
rect 381 166400 39200 166664
rect 880 166120 39200 166400
rect 381 165856 39200 166120
rect 880 165576 39120 165856
rect 381 165312 39200 165576
rect 880 165032 39200 165312
rect 381 164768 39200 165032
rect 880 164496 39200 164768
rect 880 164488 39120 164496
rect 381 164224 39120 164488
rect 880 164216 39120 164224
rect 880 163944 39200 164216
rect 381 163680 39200 163944
rect 880 163400 39200 163680
rect 381 163136 39200 163400
rect 880 162856 39120 163136
rect 381 162592 39200 162856
rect 880 162312 39200 162592
rect 381 162048 39200 162312
rect 880 161776 39200 162048
rect 880 161768 39120 161776
rect 381 161504 39120 161768
rect 880 161496 39120 161504
rect 880 161224 39200 161496
rect 381 160960 39200 161224
rect 880 160680 39200 160960
rect 381 160416 39200 160680
rect 880 160136 39120 160416
rect 381 159872 39200 160136
rect 880 159592 39200 159872
rect 381 159328 39200 159592
rect 880 159056 39200 159328
rect 880 159048 39120 159056
rect 381 158784 39120 159048
rect 880 158776 39120 158784
rect 880 158504 39200 158776
rect 381 158240 39200 158504
rect 880 157960 39200 158240
rect 381 157696 39200 157960
rect 880 157416 39120 157696
rect 381 157152 39200 157416
rect 880 156872 39200 157152
rect 381 156608 39200 156872
rect 880 156336 39200 156608
rect 880 156328 39120 156336
rect 381 156064 39120 156328
rect 880 156056 39120 156064
rect 880 155784 39200 156056
rect 381 155520 39200 155784
rect 880 155240 39200 155520
rect 381 154976 39200 155240
rect 880 154696 39120 154976
rect 381 154432 39200 154696
rect 880 154152 39200 154432
rect 381 153888 39200 154152
rect 880 153616 39200 153888
rect 880 153608 39120 153616
rect 381 153344 39120 153608
rect 880 153336 39120 153344
rect 880 153064 39200 153336
rect 381 152800 39200 153064
rect 880 152520 39200 152800
rect 381 152256 39200 152520
rect 880 151976 39120 152256
rect 381 151712 39200 151976
rect 880 151432 39200 151712
rect 381 151168 39200 151432
rect 880 150896 39200 151168
rect 880 150888 39120 150896
rect 381 150624 39120 150888
rect 880 150616 39120 150624
rect 880 150344 39200 150616
rect 381 150080 39200 150344
rect 880 149800 39200 150080
rect 381 149536 39200 149800
rect 880 149256 39120 149536
rect 381 148992 39200 149256
rect 880 148712 39200 148992
rect 381 148448 39200 148712
rect 880 148176 39200 148448
rect 880 148168 39120 148176
rect 381 147904 39120 148168
rect 880 147896 39120 147904
rect 880 147624 39200 147896
rect 381 147360 39200 147624
rect 880 147080 39200 147360
rect 381 146816 39200 147080
rect 880 146536 39120 146816
rect 381 146272 39200 146536
rect 880 145992 39200 146272
rect 381 145728 39200 145992
rect 880 145456 39200 145728
rect 880 145448 39120 145456
rect 381 145184 39120 145448
rect 880 145176 39120 145184
rect 880 144904 39200 145176
rect 381 144640 39200 144904
rect 880 144360 39200 144640
rect 381 144096 39200 144360
rect 880 143816 39120 144096
rect 381 143552 39200 143816
rect 880 143272 39200 143552
rect 381 143008 39200 143272
rect 880 142736 39200 143008
rect 880 142728 39120 142736
rect 381 142464 39120 142728
rect 880 142456 39120 142464
rect 880 142184 39200 142456
rect 381 141920 39200 142184
rect 880 141640 39200 141920
rect 381 141376 39200 141640
rect 880 141096 39120 141376
rect 381 140832 39200 141096
rect 880 140552 39200 140832
rect 381 140288 39200 140552
rect 880 140016 39200 140288
rect 880 140008 39120 140016
rect 381 139744 39120 140008
rect 880 139736 39120 139744
rect 880 139464 39200 139736
rect 381 139200 39200 139464
rect 880 138920 39200 139200
rect 381 138656 39200 138920
rect 880 138376 39120 138656
rect 381 138112 39200 138376
rect 880 137832 39200 138112
rect 381 137568 39200 137832
rect 880 137296 39200 137568
rect 880 137288 39120 137296
rect 381 137024 39120 137288
rect 880 137016 39120 137024
rect 880 136744 39200 137016
rect 381 136480 39200 136744
rect 880 136200 39200 136480
rect 381 135936 39200 136200
rect 880 135656 39120 135936
rect 381 135392 39200 135656
rect 880 135112 39200 135392
rect 381 134848 39200 135112
rect 880 134576 39200 134848
rect 880 134568 39120 134576
rect 381 134304 39120 134568
rect 880 134296 39120 134304
rect 880 134024 39200 134296
rect 381 133760 39200 134024
rect 880 133480 39200 133760
rect 381 133216 39200 133480
rect 880 132936 39120 133216
rect 381 132672 39200 132936
rect 880 132392 39200 132672
rect 381 132128 39200 132392
rect 880 131856 39200 132128
rect 880 131848 39120 131856
rect 381 131584 39120 131848
rect 880 131576 39120 131584
rect 880 131304 39200 131576
rect 381 131040 39200 131304
rect 880 130760 39200 131040
rect 381 130496 39200 130760
rect 880 130216 39120 130496
rect 381 129952 39200 130216
rect 880 129672 39200 129952
rect 381 129408 39200 129672
rect 880 129136 39200 129408
rect 880 129128 39120 129136
rect 381 128864 39120 129128
rect 880 128856 39120 128864
rect 880 128584 39200 128856
rect 381 128320 39200 128584
rect 880 128040 39200 128320
rect 381 127776 39200 128040
rect 880 127496 39120 127776
rect 381 127232 39200 127496
rect 880 126952 39200 127232
rect 381 126688 39200 126952
rect 880 126416 39200 126688
rect 880 126408 39120 126416
rect 381 126144 39120 126408
rect 880 126136 39120 126144
rect 880 125864 39200 126136
rect 381 125600 39200 125864
rect 880 125320 39200 125600
rect 381 125056 39200 125320
rect 880 124776 39120 125056
rect 381 124512 39200 124776
rect 880 124232 39200 124512
rect 381 123968 39200 124232
rect 880 123696 39200 123968
rect 880 123688 39120 123696
rect 381 123424 39120 123688
rect 880 123416 39120 123424
rect 880 123144 39200 123416
rect 381 122880 39200 123144
rect 880 122600 39200 122880
rect 381 122336 39200 122600
rect 880 122056 39120 122336
rect 381 121792 39200 122056
rect 880 121512 39200 121792
rect 381 121248 39200 121512
rect 880 120976 39200 121248
rect 880 120968 39120 120976
rect 381 120704 39120 120968
rect 880 120696 39120 120704
rect 880 120424 39200 120696
rect 381 120160 39200 120424
rect 880 119880 39200 120160
rect 381 119616 39200 119880
rect 880 119336 39120 119616
rect 381 119072 39200 119336
rect 880 118792 39200 119072
rect 381 118528 39200 118792
rect 880 118256 39200 118528
rect 880 118248 39120 118256
rect 381 117984 39120 118248
rect 880 117976 39120 117984
rect 880 117704 39200 117976
rect 381 117440 39200 117704
rect 880 117160 39200 117440
rect 381 116896 39200 117160
rect 880 116616 39120 116896
rect 381 116352 39200 116616
rect 880 116072 39200 116352
rect 381 115808 39200 116072
rect 880 115536 39200 115808
rect 880 115528 39120 115536
rect 381 115264 39120 115528
rect 880 115256 39120 115264
rect 880 114984 39200 115256
rect 381 114720 39200 114984
rect 880 114440 39200 114720
rect 381 114176 39200 114440
rect 880 113896 39120 114176
rect 381 113632 39200 113896
rect 880 113352 39200 113632
rect 381 113088 39200 113352
rect 880 112816 39200 113088
rect 880 112808 39120 112816
rect 381 112544 39120 112808
rect 880 112536 39120 112544
rect 880 112264 39200 112536
rect 381 112000 39200 112264
rect 880 111720 39200 112000
rect 381 111456 39200 111720
rect 880 111176 39120 111456
rect 381 110912 39200 111176
rect 880 110632 39200 110912
rect 381 110368 39200 110632
rect 880 110096 39200 110368
rect 880 110088 39120 110096
rect 381 109824 39120 110088
rect 880 109816 39120 109824
rect 880 109544 39200 109816
rect 381 109280 39200 109544
rect 880 109000 39200 109280
rect 381 108736 39200 109000
rect 880 108456 39120 108736
rect 381 108192 39200 108456
rect 880 107912 39200 108192
rect 381 107648 39200 107912
rect 880 107376 39200 107648
rect 880 107368 39120 107376
rect 381 107104 39120 107368
rect 880 107096 39120 107104
rect 880 106824 39200 107096
rect 381 106560 39200 106824
rect 880 106280 39200 106560
rect 381 106016 39200 106280
rect 880 105736 39120 106016
rect 381 105472 39200 105736
rect 880 105192 39200 105472
rect 381 104928 39200 105192
rect 880 104656 39200 104928
rect 880 104648 39120 104656
rect 381 104384 39120 104648
rect 880 104376 39120 104384
rect 880 104104 39200 104376
rect 381 103840 39200 104104
rect 880 103560 39200 103840
rect 381 103296 39200 103560
rect 880 103016 39120 103296
rect 381 102752 39200 103016
rect 880 102472 39200 102752
rect 381 102208 39200 102472
rect 880 101936 39200 102208
rect 880 101928 39120 101936
rect 381 101664 39120 101928
rect 880 101656 39120 101664
rect 880 101384 39200 101656
rect 381 101120 39200 101384
rect 880 100840 39200 101120
rect 381 100576 39200 100840
rect 880 100296 39120 100576
rect 381 100032 39200 100296
rect 880 99752 39200 100032
rect 381 99488 39200 99752
rect 880 99216 39200 99488
rect 880 99208 39120 99216
rect 381 98944 39120 99208
rect 880 98936 39120 98944
rect 880 98664 39200 98936
rect 381 98400 39200 98664
rect 880 98120 39200 98400
rect 381 97856 39200 98120
rect 880 97576 39120 97856
rect 381 97312 39200 97576
rect 880 97032 39200 97312
rect 381 96768 39200 97032
rect 880 96496 39200 96768
rect 880 96488 39120 96496
rect 381 96224 39120 96488
rect 880 96216 39120 96224
rect 880 95944 39200 96216
rect 381 95680 39200 95944
rect 880 95400 39200 95680
rect 381 95136 39200 95400
rect 880 94856 39120 95136
rect 381 94592 39200 94856
rect 880 94312 39200 94592
rect 381 94048 39200 94312
rect 880 93776 39200 94048
rect 880 93768 39120 93776
rect 381 93504 39120 93768
rect 880 93496 39120 93504
rect 880 93224 39200 93496
rect 381 92960 39200 93224
rect 880 92680 39200 92960
rect 381 92416 39200 92680
rect 880 92136 39120 92416
rect 381 91872 39200 92136
rect 880 91592 39200 91872
rect 381 91328 39200 91592
rect 880 91056 39200 91328
rect 880 91048 39120 91056
rect 381 90784 39120 91048
rect 880 90776 39120 90784
rect 880 90504 39200 90776
rect 381 90240 39200 90504
rect 880 89960 39200 90240
rect 381 89696 39200 89960
rect 880 89416 39120 89696
rect 381 89152 39200 89416
rect 880 88872 39200 89152
rect 381 88608 39200 88872
rect 880 88336 39200 88608
rect 880 88328 39120 88336
rect 381 88064 39120 88328
rect 880 88056 39120 88064
rect 880 87784 39200 88056
rect 381 87520 39200 87784
rect 880 87240 39200 87520
rect 381 86976 39200 87240
rect 880 86696 39120 86976
rect 381 86432 39200 86696
rect 880 86152 39200 86432
rect 381 85888 39200 86152
rect 880 85616 39200 85888
rect 880 85608 39120 85616
rect 381 85344 39120 85608
rect 880 85336 39120 85344
rect 880 85064 39200 85336
rect 381 84800 39200 85064
rect 880 84520 39200 84800
rect 381 84256 39200 84520
rect 880 83976 39120 84256
rect 381 83712 39200 83976
rect 880 83432 39200 83712
rect 381 83168 39200 83432
rect 880 82896 39200 83168
rect 880 82888 39120 82896
rect 381 82624 39120 82888
rect 880 82616 39120 82624
rect 880 82344 39200 82616
rect 381 82080 39200 82344
rect 880 81800 39200 82080
rect 381 81536 39200 81800
rect 880 81256 39120 81536
rect 381 80992 39200 81256
rect 880 80712 39200 80992
rect 381 80448 39200 80712
rect 880 80176 39200 80448
rect 880 80168 39120 80176
rect 381 79904 39120 80168
rect 880 79896 39120 79904
rect 880 79624 39200 79896
rect 381 79360 39200 79624
rect 880 79080 39200 79360
rect 381 78816 39200 79080
rect 880 78536 39120 78816
rect 381 78272 39200 78536
rect 880 77992 39200 78272
rect 381 77728 39200 77992
rect 880 77456 39200 77728
rect 880 77448 39120 77456
rect 381 77184 39120 77448
rect 880 77176 39120 77184
rect 880 76904 39200 77176
rect 381 76640 39200 76904
rect 880 76360 39200 76640
rect 381 76096 39200 76360
rect 880 75816 39120 76096
rect 381 75552 39200 75816
rect 880 75272 39200 75552
rect 381 75008 39200 75272
rect 880 74736 39200 75008
rect 880 74728 39120 74736
rect 381 74464 39120 74728
rect 880 74456 39120 74464
rect 880 74184 39200 74456
rect 381 73920 39200 74184
rect 880 73640 39200 73920
rect 381 73376 39200 73640
rect 880 73096 39120 73376
rect 381 72832 39200 73096
rect 880 72552 39200 72832
rect 381 72288 39200 72552
rect 880 72016 39200 72288
rect 880 72008 39120 72016
rect 381 71744 39120 72008
rect 880 71736 39120 71744
rect 880 71464 39200 71736
rect 381 71200 39200 71464
rect 880 70920 39200 71200
rect 381 70656 39200 70920
rect 880 70376 39120 70656
rect 381 70112 39200 70376
rect 880 69832 39200 70112
rect 381 69568 39200 69832
rect 880 69296 39200 69568
rect 880 69288 39120 69296
rect 381 69024 39120 69288
rect 880 69016 39120 69024
rect 880 68744 39200 69016
rect 381 68480 39200 68744
rect 880 68200 39200 68480
rect 381 67936 39200 68200
rect 880 67656 39120 67936
rect 381 67392 39200 67656
rect 880 67112 39200 67392
rect 381 66848 39200 67112
rect 880 66576 39200 66848
rect 880 66568 39120 66576
rect 381 66304 39120 66568
rect 880 66296 39120 66304
rect 880 66024 39200 66296
rect 381 65760 39200 66024
rect 880 65480 39200 65760
rect 381 65216 39200 65480
rect 880 64936 39120 65216
rect 381 64672 39200 64936
rect 880 64392 39200 64672
rect 381 64128 39200 64392
rect 880 63856 39200 64128
rect 880 63848 39120 63856
rect 381 63584 39120 63848
rect 880 63576 39120 63584
rect 880 63304 39200 63576
rect 381 63040 39200 63304
rect 880 62760 39200 63040
rect 381 62496 39200 62760
rect 880 62216 39120 62496
rect 381 61952 39200 62216
rect 880 61672 39200 61952
rect 381 61408 39200 61672
rect 880 61136 39200 61408
rect 880 61128 39120 61136
rect 381 60864 39120 61128
rect 880 60856 39120 60864
rect 880 60584 39200 60856
rect 381 60320 39200 60584
rect 880 60040 39200 60320
rect 381 59776 39200 60040
rect 880 59496 39120 59776
rect 381 59232 39200 59496
rect 880 58952 39200 59232
rect 381 58688 39200 58952
rect 880 58416 39200 58688
rect 880 58408 39120 58416
rect 381 58144 39120 58408
rect 880 58136 39120 58144
rect 880 57864 39200 58136
rect 381 57600 39200 57864
rect 880 57320 39200 57600
rect 381 57056 39200 57320
rect 880 56776 39120 57056
rect 381 56512 39200 56776
rect 880 56232 39200 56512
rect 381 55968 39200 56232
rect 880 55696 39200 55968
rect 880 55688 39120 55696
rect 381 55424 39120 55688
rect 880 55416 39120 55424
rect 880 55144 39200 55416
rect 381 54880 39200 55144
rect 880 54600 39200 54880
rect 381 54336 39200 54600
rect 880 54056 39120 54336
rect 381 53792 39200 54056
rect 880 53512 39200 53792
rect 381 53248 39200 53512
rect 880 52976 39200 53248
rect 880 52968 39120 52976
rect 381 52704 39120 52968
rect 880 52696 39120 52704
rect 880 52424 39200 52696
rect 381 52160 39200 52424
rect 880 51880 39200 52160
rect 381 51616 39200 51880
rect 880 51336 39120 51616
rect 381 51072 39200 51336
rect 880 50792 39200 51072
rect 381 50528 39200 50792
rect 880 50256 39200 50528
rect 880 50248 39120 50256
rect 381 49984 39120 50248
rect 880 49976 39120 49984
rect 880 49704 39200 49976
rect 381 49440 39200 49704
rect 880 49160 39200 49440
rect 381 48896 39200 49160
rect 880 48616 39120 48896
rect 381 48352 39200 48616
rect 880 48072 39200 48352
rect 381 47808 39200 48072
rect 880 47536 39200 47808
rect 880 47528 39120 47536
rect 381 47264 39120 47528
rect 880 47256 39120 47264
rect 880 46984 39200 47256
rect 381 46720 39200 46984
rect 880 46440 39200 46720
rect 381 46176 39200 46440
rect 880 45896 39120 46176
rect 381 45632 39200 45896
rect 880 45352 39200 45632
rect 381 45088 39200 45352
rect 880 44816 39200 45088
rect 880 44808 39120 44816
rect 381 44544 39120 44808
rect 880 44536 39120 44544
rect 880 44264 39200 44536
rect 381 44000 39200 44264
rect 880 43720 39200 44000
rect 381 43456 39200 43720
rect 880 43176 39120 43456
rect 381 42912 39200 43176
rect 880 42632 39200 42912
rect 381 42368 39200 42632
rect 880 42096 39200 42368
rect 880 42088 39120 42096
rect 381 41824 39120 42088
rect 880 41816 39120 41824
rect 880 41544 39200 41816
rect 381 41280 39200 41544
rect 880 41000 39200 41280
rect 381 40736 39200 41000
rect 880 40456 39120 40736
rect 381 40192 39200 40456
rect 880 39912 39200 40192
rect 381 39648 39200 39912
rect 880 39376 39200 39648
rect 880 39368 39120 39376
rect 381 39104 39120 39368
rect 880 39096 39120 39104
rect 880 38824 39200 39096
rect 381 38560 39200 38824
rect 880 38280 39200 38560
rect 381 38016 39200 38280
rect 880 37736 39120 38016
rect 381 37472 39200 37736
rect 880 37192 39200 37472
rect 381 36928 39200 37192
rect 880 36656 39200 36928
rect 880 36648 39120 36656
rect 381 36384 39120 36648
rect 880 36376 39120 36384
rect 880 36104 39200 36376
rect 381 35840 39200 36104
rect 880 35560 39200 35840
rect 381 35296 39200 35560
rect 880 35016 39120 35296
rect 381 34752 39200 35016
rect 880 34472 39200 34752
rect 381 34208 39200 34472
rect 880 33936 39200 34208
rect 880 33928 39120 33936
rect 381 33664 39120 33928
rect 880 33656 39120 33664
rect 880 33384 39200 33656
rect 381 33120 39200 33384
rect 880 32840 39200 33120
rect 381 32576 39200 32840
rect 880 32296 39120 32576
rect 381 32032 39200 32296
rect 880 31752 39200 32032
rect 381 31488 39200 31752
rect 880 31216 39200 31488
rect 880 31208 39120 31216
rect 381 30936 39120 31208
rect 381 29856 39200 30936
rect 381 29576 39120 29856
rect 381 28496 39200 29576
rect 381 28216 39120 28496
rect 381 27136 39200 28216
rect 381 26856 39120 27136
rect 381 25776 39200 26856
rect 381 25496 39120 25776
rect 381 24416 39200 25496
rect 381 24136 39120 24416
rect 381 23056 39200 24136
rect 381 22776 39120 23056
rect 381 21696 39200 22776
rect 381 21416 39120 21696
rect 381 20336 39200 21416
rect 381 20056 39120 20336
rect 381 18976 39200 20056
rect 381 18696 39120 18976
rect 381 17616 39200 18696
rect 381 17336 39120 17616
rect 381 16256 39200 17336
rect 381 15976 39120 16256
rect 381 14896 39200 15976
rect 381 14616 39120 14896
rect 381 13536 39200 14616
rect 381 13256 39120 13536
rect 381 12176 39200 13256
rect 381 11896 39120 12176
rect 381 10816 39200 11896
rect 381 10536 39120 10816
rect 381 9456 39200 10536
rect 381 9176 39120 9456
rect 381 8096 39200 9176
rect 381 7816 39120 8096
rect 381 6736 39200 7816
rect 381 6456 39120 6736
rect 381 5376 39200 6456
rect 381 5096 39120 5376
rect 381 4016 39200 5096
rect 381 3736 39120 4016
rect 381 2656 39200 3736
rect 381 2376 39120 2656
rect 381 1296 39200 2376
rect 381 1123 39120 1296
<< metal4 >>
rect 4208 2128 4528 197520
rect 19568 2128 19888 197520
rect 34928 2128 35248 197520
<< obsm4 >>
rect 611 3435 4128 160173
rect 4608 3435 19488 160173
rect 19968 3435 34848 160173
rect 35328 3435 37109 160173
<< labels >>
rlabel metal3 s 0 31288 800 31408 6 custom_settings[0]
port 1 nsew signal output
rlabel metal3 s 0 36728 800 36848 6 custom_settings[10]
port 2 nsew signal output
rlabel metal3 s 0 37272 800 37392 6 custom_settings[11]
port 3 nsew signal output
rlabel metal3 s 0 37816 800 37936 6 custom_settings[12]
port 4 nsew signal output
rlabel metal3 s 0 38360 800 38480 6 custom_settings[13]
port 5 nsew signal output
rlabel metal3 s 0 38904 800 39024 6 custom_settings[14]
port 6 nsew signal output
rlabel metal3 s 0 39448 800 39568 6 custom_settings[15]
port 7 nsew signal output
rlabel metal3 s 0 39992 800 40112 6 custom_settings[16]
port 8 nsew signal output
rlabel metal3 s 0 40536 800 40656 6 custom_settings[17]
port 9 nsew signal output
rlabel metal3 s 0 41080 800 41200 6 custom_settings[18]
port 10 nsew signal output
rlabel metal3 s 0 41624 800 41744 6 custom_settings[19]
port 11 nsew signal output
rlabel metal3 s 0 31832 800 31952 6 custom_settings[1]
port 12 nsew signal output
rlabel metal3 s 0 42168 800 42288 6 custom_settings[20]
port 13 nsew signal output
rlabel metal3 s 0 42712 800 42832 6 custom_settings[21]
port 14 nsew signal output
rlabel metal3 s 0 43256 800 43376 6 custom_settings[22]
port 15 nsew signal output
rlabel metal3 s 0 43800 800 43920 6 custom_settings[23]
port 16 nsew signal output
rlabel metal3 s 0 44344 800 44464 6 custom_settings[24]
port 17 nsew signal output
rlabel metal3 s 0 44888 800 45008 6 custom_settings[25]
port 18 nsew signal output
rlabel metal3 s 0 45432 800 45552 6 custom_settings[26]
port 19 nsew signal output
rlabel metal3 s 0 45976 800 46096 6 custom_settings[27]
port 20 nsew signal output
rlabel metal3 s 0 46520 800 46640 6 custom_settings[28]
port 21 nsew signal output
rlabel metal3 s 0 47064 800 47184 6 custom_settings[29]
port 22 nsew signal output
rlabel metal3 s 0 32376 800 32496 6 custom_settings[2]
port 23 nsew signal output
rlabel metal3 s 0 47608 800 47728 6 custom_settings[30]
port 24 nsew signal output
rlabel metal3 s 0 48152 800 48272 6 custom_settings[31]
port 25 nsew signal output
rlabel metal3 s 0 32920 800 33040 6 custom_settings[3]
port 26 nsew signal output
rlabel metal3 s 0 33464 800 33584 6 custom_settings[4]
port 27 nsew signal output
rlabel metal3 s 0 34008 800 34128 6 custom_settings[5]
port 28 nsew signal output
rlabel metal3 s 0 34552 800 34672 6 custom_settings[6]
port 29 nsew signal output
rlabel metal3 s 0 35096 800 35216 6 custom_settings[7]
port 30 nsew signal output
rlabel metal3 s 0 35640 800 35760 6 custom_settings[8]
port 31 nsew signal output
rlabel metal3 s 0 36184 800 36304 6 custom_settings[9]
port 32 nsew signal output
rlabel metal2 s 754 199200 810 200000 6 io_in_0
port 33 nsew signal input
rlabel metal3 s 0 48696 800 48816 6 io_oeb[0]
port 34 nsew signal output
rlabel metal3 s 0 54136 800 54256 6 io_oeb[10]
port 35 nsew signal output
rlabel metal3 s 0 54680 800 54800 6 io_oeb[11]
port 36 nsew signal output
rlabel metal3 s 0 55224 800 55344 6 io_oeb[12]
port 37 nsew signal output
rlabel metal3 s 0 55768 800 55888 6 io_oeb[13]
port 38 nsew signal output
rlabel metal3 s 0 56312 800 56432 6 io_oeb[14]
port 39 nsew signal output
rlabel metal3 s 0 56856 800 56976 6 io_oeb[15]
port 40 nsew signal output
rlabel metal3 s 0 57400 800 57520 6 io_oeb[16]
port 41 nsew signal output
rlabel metal3 s 0 57944 800 58064 6 io_oeb[17]
port 42 nsew signal output
rlabel metal3 s 0 58488 800 58608 6 io_oeb[18]
port 43 nsew signal output
rlabel metal3 s 0 59032 800 59152 6 io_oeb[19]
port 44 nsew signal output
rlabel metal3 s 0 49240 800 49360 6 io_oeb[1]
port 45 nsew signal output
rlabel metal3 s 0 59576 800 59696 6 io_oeb[20]
port 46 nsew signal output
rlabel metal3 s 0 60120 800 60240 6 io_oeb[21]
port 47 nsew signal output
rlabel metal3 s 0 60664 800 60784 6 io_oeb[22]
port 48 nsew signal output
rlabel metal3 s 0 61208 800 61328 6 io_oeb[23]
port 49 nsew signal output
rlabel metal3 s 0 61752 800 61872 6 io_oeb[24]
port 50 nsew signal output
rlabel metal3 s 0 62296 800 62416 6 io_oeb[25]
port 51 nsew signal output
rlabel metal3 s 0 62840 800 62960 6 io_oeb[26]
port 52 nsew signal output
rlabel metal3 s 0 63384 800 63504 6 io_oeb[27]
port 53 nsew signal output
rlabel metal3 s 0 63928 800 64048 6 io_oeb[28]
port 54 nsew signal output
rlabel metal3 s 0 64472 800 64592 6 io_oeb[29]
port 55 nsew signal output
rlabel metal3 s 0 49784 800 49904 6 io_oeb[2]
port 56 nsew signal output
rlabel metal3 s 0 65016 800 65136 6 io_oeb[30]
port 57 nsew signal output
rlabel metal3 s 0 65560 800 65680 6 io_oeb[31]
port 58 nsew signal output
rlabel metal3 s 0 66104 800 66224 6 io_oeb[32]
port 59 nsew signal output
rlabel metal3 s 0 66648 800 66768 6 io_oeb[33]
port 60 nsew signal output
rlabel metal3 s 0 67192 800 67312 6 io_oeb[34]
port 61 nsew signal output
rlabel metal3 s 0 67736 800 67856 6 io_oeb[35]
port 62 nsew signal output
rlabel metal3 s 0 68280 800 68400 6 io_oeb[36]
port 63 nsew signal output
rlabel metal3 s 0 68824 800 68944 6 io_oeb[37]
port 64 nsew signal output
rlabel metal3 s 0 50328 800 50448 6 io_oeb[3]
port 65 nsew signal output
rlabel metal3 s 0 50872 800 50992 6 io_oeb[4]
port 66 nsew signal output
rlabel metal3 s 0 51416 800 51536 6 io_oeb[5]
port 67 nsew signal output
rlabel metal3 s 0 51960 800 52080 6 io_oeb[6]
port 68 nsew signal output
rlabel metal3 s 0 52504 800 52624 6 io_oeb[7]
port 69 nsew signal output
rlabel metal3 s 0 53048 800 53168 6 io_oeb[8]
port 70 nsew signal output
rlabel metal3 s 0 53592 800 53712 6 io_oeb[9]
port 71 nsew signal output
rlabel metal3 s 0 110168 800 110288 6 io_oeb_scrapcpu[0]
port 72 nsew signal input
rlabel metal3 s 0 115608 800 115728 6 io_oeb_scrapcpu[10]
port 73 nsew signal input
rlabel metal3 s 0 116152 800 116272 6 io_oeb_scrapcpu[11]
port 74 nsew signal input
rlabel metal3 s 0 116696 800 116816 6 io_oeb_scrapcpu[12]
port 75 nsew signal input
rlabel metal3 s 0 117240 800 117360 6 io_oeb_scrapcpu[13]
port 76 nsew signal input
rlabel metal3 s 0 117784 800 117904 6 io_oeb_scrapcpu[14]
port 77 nsew signal input
rlabel metal3 s 0 118328 800 118448 6 io_oeb_scrapcpu[15]
port 78 nsew signal input
rlabel metal3 s 0 118872 800 118992 6 io_oeb_scrapcpu[16]
port 79 nsew signal input
rlabel metal3 s 0 119416 800 119536 6 io_oeb_scrapcpu[17]
port 80 nsew signal input
rlabel metal3 s 0 119960 800 120080 6 io_oeb_scrapcpu[18]
port 81 nsew signal input
rlabel metal3 s 0 120504 800 120624 6 io_oeb_scrapcpu[19]
port 82 nsew signal input
rlabel metal3 s 0 110712 800 110832 6 io_oeb_scrapcpu[1]
port 83 nsew signal input
rlabel metal3 s 0 121048 800 121168 6 io_oeb_scrapcpu[20]
port 84 nsew signal input
rlabel metal3 s 0 121592 800 121712 6 io_oeb_scrapcpu[21]
port 85 nsew signal input
rlabel metal3 s 0 122136 800 122256 6 io_oeb_scrapcpu[22]
port 86 nsew signal input
rlabel metal3 s 0 122680 800 122800 6 io_oeb_scrapcpu[23]
port 87 nsew signal input
rlabel metal3 s 0 123224 800 123344 6 io_oeb_scrapcpu[24]
port 88 nsew signal input
rlabel metal3 s 0 123768 800 123888 6 io_oeb_scrapcpu[25]
port 89 nsew signal input
rlabel metal3 s 0 124312 800 124432 6 io_oeb_scrapcpu[26]
port 90 nsew signal input
rlabel metal3 s 0 124856 800 124976 6 io_oeb_scrapcpu[27]
port 91 nsew signal input
rlabel metal3 s 0 125400 800 125520 6 io_oeb_scrapcpu[28]
port 92 nsew signal input
rlabel metal3 s 0 125944 800 126064 6 io_oeb_scrapcpu[29]
port 93 nsew signal input
rlabel metal3 s 0 111256 800 111376 6 io_oeb_scrapcpu[2]
port 94 nsew signal input
rlabel metal3 s 0 126488 800 126608 6 io_oeb_scrapcpu[30]
port 95 nsew signal input
rlabel metal3 s 0 127032 800 127152 6 io_oeb_scrapcpu[31]
port 96 nsew signal input
rlabel metal3 s 0 127576 800 127696 6 io_oeb_scrapcpu[32]
port 97 nsew signal input
rlabel metal3 s 0 128120 800 128240 6 io_oeb_scrapcpu[33]
port 98 nsew signal input
rlabel metal3 s 0 128664 800 128784 6 io_oeb_scrapcpu[34]
port 99 nsew signal input
rlabel metal3 s 0 129208 800 129328 6 io_oeb_scrapcpu[35]
port 100 nsew signal input
rlabel metal3 s 0 111800 800 111920 6 io_oeb_scrapcpu[3]
port 101 nsew signal input
rlabel metal3 s 0 112344 800 112464 6 io_oeb_scrapcpu[4]
port 102 nsew signal input
rlabel metal3 s 0 112888 800 113008 6 io_oeb_scrapcpu[5]
port 103 nsew signal input
rlabel metal3 s 0 113432 800 113552 6 io_oeb_scrapcpu[6]
port 104 nsew signal input
rlabel metal3 s 0 113976 800 114096 6 io_oeb_scrapcpu[7]
port 105 nsew signal input
rlabel metal3 s 0 114520 800 114640 6 io_oeb_scrapcpu[8]
port 106 nsew signal input
rlabel metal3 s 0 115064 800 115184 6 io_oeb_scrapcpu[9]
port 107 nsew signal input
rlabel metal3 s 0 149336 800 149456 6 io_oeb_vliw[0]
port 108 nsew signal input
rlabel metal3 s 0 154776 800 154896 6 io_oeb_vliw[10]
port 109 nsew signal input
rlabel metal3 s 0 155320 800 155440 6 io_oeb_vliw[11]
port 110 nsew signal input
rlabel metal3 s 0 155864 800 155984 6 io_oeb_vliw[12]
port 111 nsew signal input
rlabel metal3 s 0 156408 800 156528 6 io_oeb_vliw[13]
port 112 nsew signal input
rlabel metal3 s 0 156952 800 157072 6 io_oeb_vliw[14]
port 113 nsew signal input
rlabel metal3 s 0 157496 800 157616 6 io_oeb_vliw[15]
port 114 nsew signal input
rlabel metal3 s 0 158040 800 158160 6 io_oeb_vliw[16]
port 115 nsew signal input
rlabel metal3 s 0 158584 800 158704 6 io_oeb_vliw[17]
port 116 nsew signal input
rlabel metal3 s 0 159128 800 159248 6 io_oeb_vliw[18]
port 117 nsew signal input
rlabel metal3 s 0 159672 800 159792 6 io_oeb_vliw[19]
port 118 nsew signal input
rlabel metal3 s 0 149880 800 150000 6 io_oeb_vliw[1]
port 119 nsew signal input
rlabel metal3 s 0 160216 800 160336 6 io_oeb_vliw[20]
port 120 nsew signal input
rlabel metal3 s 0 160760 800 160880 6 io_oeb_vliw[21]
port 121 nsew signal input
rlabel metal3 s 0 161304 800 161424 6 io_oeb_vliw[22]
port 122 nsew signal input
rlabel metal3 s 0 161848 800 161968 6 io_oeb_vliw[23]
port 123 nsew signal input
rlabel metal3 s 0 162392 800 162512 6 io_oeb_vliw[24]
port 124 nsew signal input
rlabel metal3 s 0 162936 800 163056 6 io_oeb_vliw[25]
port 125 nsew signal input
rlabel metal3 s 0 163480 800 163600 6 io_oeb_vliw[26]
port 126 nsew signal input
rlabel metal3 s 0 164024 800 164144 6 io_oeb_vliw[27]
port 127 nsew signal input
rlabel metal3 s 0 164568 800 164688 6 io_oeb_vliw[28]
port 128 nsew signal input
rlabel metal3 s 0 165112 800 165232 6 io_oeb_vliw[29]
port 129 nsew signal input
rlabel metal3 s 0 150424 800 150544 6 io_oeb_vliw[2]
port 130 nsew signal input
rlabel metal3 s 0 165656 800 165776 6 io_oeb_vliw[30]
port 131 nsew signal input
rlabel metal3 s 0 166200 800 166320 6 io_oeb_vliw[31]
port 132 nsew signal input
rlabel metal3 s 0 166744 800 166864 6 io_oeb_vliw[32]
port 133 nsew signal input
rlabel metal3 s 0 167288 800 167408 6 io_oeb_vliw[33]
port 134 nsew signal input
rlabel metal3 s 0 167832 800 167952 6 io_oeb_vliw[34]
port 135 nsew signal input
rlabel metal3 s 0 168376 800 168496 6 io_oeb_vliw[35]
port 136 nsew signal input
rlabel metal3 s 0 150968 800 151088 6 io_oeb_vliw[3]
port 137 nsew signal input
rlabel metal3 s 0 151512 800 151632 6 io_oeb_vliw[4]
port 138 nsew signal input
rlabel metal3 s 0 152056 800 152176 6 io_oeb_vliw[5]
port 139 nsew signal input
rlabel metal3 s 0 152600 800 152720 6 io_oeb_vliw[6]
port 140 nsew signal input
rlabel metal3 s 0 153144 800 153264 6 io_oeb_vliw[7]
port 141 nsew signal input
rlabel metal3 s 0 153688 800 153808 6 io_oeb_vliw[8]
port 142 nsew signal input
rlabel metal3 s 0 154232 800 154352 6 io_oeb_vliw[9]
port 143 nsew signal input
rlabel metal3 s 0 129752 800 129872 6 io_oeb_z80[0]
port 144 nsew signal input
rlabel metal3 s 0 135192 800 135312 6 io_oeb_z80[10]
port 145 nsew signal input
rlabel metal3 s 0 135736 800 135856 6 io_oeb_z80[11]
port 146 nsew signal input
rlabel metal3 s 0 136280 800 136400 6 io_oeb_z80[12]
port 147 nsew signal input
rlabel metal3 s 0 136824 800 136944 6 io_oeb_z80[13]
port 148 nsew signal input
rlabel metal3 s 0 137368 800 137488 6 io_oeb_z80[14]
port 149 nsew signal input
rlabel metal3 s 0 137912 800 138032 6 io_oeb_z80[15]
port 150 nsew signal input
rlabel metal3 s 0 138456 800 138576 6 io_oeb_z80[16]
port 151 nsew signal input
rlabel metal3 s 0 139000 800 139120 6 io_oeb_z80[17]
port 152 nsew signal input
rlabel metal3 s 0 139544 800 139664 6 io_oeb_z80[18]
port 153 nsew signal input
rlabel metal3 s 0 140088 800 140208 6 io_oeb_z80[19]
port 154 nsew signal input
rlabel metal3 s 0 130296 800 130416 6 io_oeb_z80[1]
port 155 nsew signal input
rlabel metal3 s 0 140632 800 140752 6 io_oeb_z80[20]
port 156 nsew signal input
rlabel metal3 s 0 141176 800 141296 6 io_oeb_z80[21]
port 157 nsew signal input
rlabel metal3 s 0 141720 800 141840 6 io_oeb_z80[22]
port 158 nsew signal input
rlabel metal3 s 0 142264 800 142384 6 io_oeb_z80[23]
port 159 nsew signal input
rlabel metal3 s 0 142808 800 142928 6 io_oeb_z80[24]
port 160 nsew signal input
rlabel metal3 s 0 143352 800 143472 6 io_oeb_z80[25]
port 161 nsew signal input
rlabel metal3 s 0 143896 800 144016 6 io_oeb_z80[26]
port 162 nsew signal input
rlabel metal3 s 0 144440 800 144560 6 io_oeb_z80[27]
port 163 nsew signal input
rlabel metal3 s 0 144984 800 145104 6 io_oeb_z80[28]
port 164 nsew signal input
rlabel metal3 s 0 145528 800 145648 6 io_oeb_z80[29]
port 165 nsew signal input
rlabel metal3 s 0 130840 800 130960 6 io_oeb_z80[2]
port 166 nsew signal input
rlabel metal3 s 0 146072 800 146192 6 io_oeb_z80[30]
port 167 nsew signal input
rlabel metal3 s 0 146616 800 146736 6 io_oeb_z80[31]
port 168 nsew signal input
rlabel metal3 s 0 147160 800 147280 6 io_oeb_z80[32]
port 169 nsew signal input
rlabel metal3 s 0 147704 800 147824 6 io_oeb_z80[33]
port 170 nsew signal input
rlabel metal3 s 0 148248 800 148368 6 io_oeb_z80[34]
port 171 nsew signal input
rlabel metal3 s 0 148792 800 148912 6 io_oeb_z80[35]
port 172 nsew signal input
rlabel metal3 s 0 131384 800 131504 6 io_oeb_z80[3]
port 173 nsew signal input
rlabel metal3 s 0 131928 800 132048 6 io_oeb_z80[4]
port 174 nsew signal input
rlabel metal3 s 0 132472 800 132592 6 io_oeb_z80[5]
port 175 nsew signal input
rlabel metal3 s 0 133016 800 133136 6 io_oeb_z80[6]
port 176 nsew signal input
rlabel metal3 s 0 133560 800 133680 6 io_oeb_z80[7]
port 177 nsew signal input
rlabel metal3 s 0 134104 800 134224 6 io_oeb_z80[8]
port 178 nsew signal input
rlabel metal3 s 0 134648 800 134768 6 io_oeb_z80[9]
port 179 nsew signal input
rlabel metal3 s 39200 1096 40000 1216 6 io_out[0]
port 180 nsew signal output
rlabel metal3 s 39200 14696 40000 14816 6 io_out[10]
port 181 nsew signal output
rlabel metal3 s 39200 16056 40000 16176 6 io_out[11]
port 182 nsew signal output
rlabel metal3 s 39200 17416 40000 17536 6 io_out[12]
port 183 nsew signal output
rlabel metal3 s 39200 18776 40000 18896 6 io_out[13]
port 184 nsew signal output
rlabel metal3 s 39200 20136 40000 20256 6 io_out[14]
port 185 nsew signal output
rlabel metal3 s 39200 21496 40000 21616 6 io_out[15]
port 186 nsew signal output
rlabel metal3 s 39200 22856 40000 22976 6 io_out[16]
port 187 nsew signal output
rlabel metal3 s 39200 24216 40000 24336 6 io_out[17]
port 188 nsew signal output
rlabel metal3 s 39200 25576 40000 25696 6 io_out[18]
port 189 nsew signal output
rlabel metal3 s 39200 26936 40000 27056 6 io_out[19]
port 190 nsew signal output
rlabel metal3 s 39200 2456 40000 2576 6 io_out[1]
port 191 nsew signal output
rlabel metal3 s 39200 28296 40000 28416 6 io_out[20]
port 192 nsew signal output
rlabel metal3 s 39200 29656 40000 29776 6 io_out[21]
port 193 nsew signal output
rlabel metal3 s 39200 31016 40000 31136 6 io_out[22]
port 194 nsew signal output
rlabel metal3 s 39200 32376 40000 32496 6 io_out[23]
port 195 nsew signal output
rlabel metal3 s 39200 33736 40000 33856 6 io_out[24]
port 196 nsew signal output
rlabel metal3 s 39200 35096 40000 35216 6 io_out[25]
port 197 nsew signal output
rlabel metal3 s 39200 36456 40000 36576 6 io_out[26]
port 198 nsew signal output
rlabel metal3 s 39200 37816 40000 37936 6 io_out[27]
port 199 nsew signal output
rlabel metal3 s 39200 39176 40000 39296 6 io_out[28]
port 200 nsew signal output
rlabel metal3 s 39200 40536 40000 40656 6 io_out[29]
port 201 nsew signal output
rlabel metal3 s 39200 3816 40000 3936 6 io_out[2]
port 202 nsew signal output
rlabel metal3 s 39200 41896 40000 42016 6 io_out[30]
port 203 nsew signal output
rlabel metal3 s 39200 43256 40000 43376 6 io_out[31]
port 204 nsew signal output
rlabel metal3 s 39200 44616 40000 44736 6 io_out[32]
port 205 nsew signal output
rlabel metal3 s 39200 45976 40000 46096 6 io_out[33]
port 206 nsew signal output
rlabel metal3 s 39200 47336 40000 47456 6 io_out[34]
port 207 nsew signal output
rlabel metal3 s 39200 48696 40000 48816 6 io_out[35]
port 208 nsew signal output
rlabel metal3 s 39200 50056 40000 50176 6 io_out[36]
port 209 nsew signal output
rlabel metal3 s 39200 51416 40000 51536 6 io_out[37]
port 210 nsew signal output
rlabel metal3 s 39200 5176 40000 5296 6 io_out[3]
port 211 nsew signal output
rlabel metal3 s 39200 6536 40000 6656 6 io_out[4]
port 212 nsew signal output
rlabel metal3 s 39200 7896 40000 8016 6 io_out[5]
port 213 nsew signal output
rlabel metal3 s 39200 9256 40000 9376 6 io_out[6]
port 214 nsew signal output
rlabel metal3 s 39200 10616 40000 10736 6 io_out[7]
port 215 nsew signal output
rlabel metal3 s 39200 11976 40000 12096 6 io_out[8]
port 216 nsew signal output
rlabel metal3 s 39200 13336 40000 13456 6 io_out[9]
port 217 nsew signal output
rlabel metal3 s 0 69912 800 70032 6 io_out_scrapcpu[0]
port 218 nsew signal input
rlabel metal3 s 0 75352 800 75472 6 io_out_scrapcpu[10]
port 219 nsew signal input
rlabel metal3 s 0 75896 800 76016 6 io_out_scrapcpu[11]
port 220 nsew signal input
rlabel metal3 s 0 76440 800 76560 6 io_out_scrapcpu[12]
port 221 nsew signal input
rlabel metal3 s 0 76984 800 77104 6 io_out_scrapcpu[13]
port 222 nsew signal input
rlabel metal3 s 0 77528 800 77648 6 io_out_scrapcpu[14]
port 223 nsew signal input
rlabel metal3 s 0 78072 800 78192 6 io_out_scrapcpu[15]
port 224 nsew signal input
rlabel metal3 s 0 78616 800 78736 6 io_out_scrapcpu[16]
port 225 nsew signal input
rlabel metal3 s 0 79160 800 79280 6 io_out_scrapcpu[17]
port 226 nsew signal input
rlabel metal3 s 0 79704 800 79824 6 io_out_scrapcpu[18]
port 227 nsew signal input
rlabel metal3 s 0 80248 800 80368 6 io_out_scrapcpu[19]
port 228 nsew signal input
rlabel metal3 s 0 70456 800 70576 6 io_out_scrapcpu[1]
port 229 nsew signal input
rlabel metal3 s 0 80792 800 80912 6 io_out_scrapcpu[20]
port 230 nsew signal input
rlabel metal3 s 0 81336 800 81456 6 io_out_scrapcpu[21]
port 231 nsew signal input
rlabel metal3 s 0 81880 800 82000 6 io_out_scrapcpu[22]
port 232 nsew signal input
rlabel metal3 s 0 82424 800 82544 6 io_out_scrapcpu[23]
port 233 nsew signal input
rlabel metal3 s 0 82968 800 83088 6 io_out_scrapcpu[24]
port 234 nsew signal input
rlabel metal3 s 0 83512 800 83632 6 io_out_scrapcpu[25]
port 235 nsew signal input
rlabel metal3 s 0 84056 800 84176 6 io_out_scrapcpu[26]
port 236 nsew signal input
rlabel metal3 s 0 84600 800 84720 6 io_out_scrapcpu[27]
port 237 nsew signal input
rlabel metal3 s 0 85144 800 85264 6 io_out_scrapcpu[28]
port 238 nsew signal input
rlabel metal3 s 0 85688 800 85808 6 io_out_scrapcpu[29]
port 239 nsew signal input
rlabel metal3 s 0 71000 800 71120 6 io_out_scrapcpu[2]
port 240 nsew signal input
rlabel metal3 s 0 86232 800 86352 6 io_out_scrapcpu[30]
port 241 nsew signal input
rlabel metal3 s 0 86776 800 86896 6 io_out_scrapcpu[31]
port 242 nsew signal input
rlabel metal3 s 0 87320 800 87440 6 io_out_scrapcpu[32]
port 243 nsew signal input
rlabel metal3 s 0 87864 800 87984 6 io_out_scrapcpu[33]
port 244 nsew signal input
rlabel metal3 s 0 88408 800 88528 6 io_out_scrapcpu[34]
port 245 nsew signal input
rlabel metal3 s 0 88952 800 89072 6 io_out_scrapcpu[35]
port 246 nsew signal input
rlabel metal3 s 0 71544 800 71664 6 io_out_scrapcpu[3]
port 247 nsew signal input
rlabel metal3 s 0 72088 800 72208 6 io_out_scrapcpu[4]
port 248 nsew signal input
rlabel metal3 s 0 72632 800 72752 6 io_out_scrapcpu[5]
port 249 nsew signal input
rlabel metal3 s 0 73176 800 73296 6 io_out_scrapcpu[6]
port 250 nsew signal input
rlabel metal3 s 0 73720 800 73840 6 io_out_scrapcpu[7]
port 251 nsew signal input
rlabel metal3 s 0 74264 800 74384 6 io_out_scrapcpu[8]
port 252 nsew signal input
rlabel metal3 s 0 74808 800 74928 6 io_out_scrapcpu[9]
port 253 nsew signal input
rlabel metal2 s 3790 199200 3846 200000 6 io_out_vliw[0]
port 254 nsew signal input
rlabel metal2 s 13910 199200 13966 200000 6 io_out_vliw[10]
port 255 nsew signal input
rlabel metal2 s 14922 199200 14978 200000 6 io_out_vliw[11]
port 256 nsew signal input
rlabel metal2 s 15934 199200 15990 200000 6 io_out_vliw[12]
port 257 nsew signal input
rlabel metal2 s 16946 199200 17002 200000 6 io_out_vliw[13]
port 258 nsew signal input
rlabel metal2 s 17958 199200 18014 200000 6 io_out_vliw[14]
port 259 nsew signal input
rlabel metal2 s 18970 199200 19026 200000 6 io_out_vliw[15]
port 260 nsew signal input
rlabel metal2 s 19982 199200 20038 200000 6 io_out_vliw[16]
port 261 nsew signal input
rlabel metal2 s 20994 199200 21050 200000 6 io_out_vliw[17]
port 262 nsew signal input
rlabel metal2 s 22006 199200 22062 200000 6 io_out_vliw[18]
port 263 nsew signal input
rlabel metal2 s 23018 199200 23074 200000 6 io_out_vliw[19]
port 264 nsew signal input
rlabel metal2 s 4802 199200 4858 200000 6 io_out_vliw[1]
port 265 nsew signal input
rlabel metal2 s 24030 199200 24086 200000 6 io_out_vliw[20]
port 266 nsew signal input
rlabel metal2 s 25042 199200 25098 200000 6 io_out_vliw[21]
port 267 nsew signal input
rlabel metal2 s 26054 199200 26110 200000 6 io_out_vliw[22]
port 268 nsew signal input
rlabel metal2 s 27066 199200 27122 200000 6 io_out_vliw[23]
port 269 nsew signal input
rlabel metal2 s 28078 199200 28134 200000 6 io_out_vliw[24]
port 270 nsew signal input
rlabel metal2 s 29090 199200 29146 200000 6 io_out_vliw[25]
port 271 nsew signal input
rlabel metal2 s 30102 199200 30158 200000 6 io_out_vliw[26]
port 272 nsew signal input
rlabel metal2 s 31114 199200 31170 200000 6 io_out_vliw[27]
port 273 nsew signal input
rlabel metal2 s 32126 199200 32182 200000 6 io_out_vliw[28]
port 274 nsew signal input
rlabel metal2 s 33138 199200 33194 200000 6 io_out_vliw[29]
port 275 nsew signal input
rlabel metal2 s 5814 199200 5870 200000 6 io_out_vliw[2]
port 276 nsew signal input
rlabel metal2 s 34150 199200 34206 200000 6 io_out_vliw[30]
port 277 nsew signal input
rlabel metal2 s 35162 199200 35218 200000 6 io_out_vliw[31]
port 278 nsew signal input
rlabel metal2 s 36174 199200 36230 200000 6 io_out_vliw[32]
port 279 nsew signal input
rlabel metal2 s 37186 199200 37242 200000 6 io_out_vliw[33]
port 280 nsew signal input
rlabel metal2 s 38198 199200 38254 200000 6 io_out_vliw[34]
port 281 nsew signal input
rlabel metal2 s 39210 199200 39266 200000 6 io_out_vliw[35]
port 282 nsew signal input
rlabel metal2 s 6826 199200 6882 200000 6 io_out_vliw[3]
port 283 nsew signal input
rlabel metal2 s 7838 199200 7894 200000 6 io_out_vliw[4]
port 284 nsew signal input
rlabel metal2 s 8850 199200 8906 200000 6 io_out_vliw[5]
port 285 nsew signal input
rlabel metal2 s 9862 199200 9918 200000 6 io_out_vliw[6]
port 286 nsew signal input
rlabel metal2 s 10874 199200 10930 200000 6 io_out_vliw[7]
port 287 nsew signal input
rlabel metal2 s 11886 199200 11942 200000 6 io_out_vliw[8]
port 288 nsew signal input
rlabel metal2 s 12898 199200 12954 200000 6 io_out_vliw[9]
port 289 nsew signal input
rlabel metal3 s 39200 150696 40000 150816 6 io_out_z80[0]
port 290 nsew signal input
rlabel metal3 s 39200 164296 40000 164416 6 io_out_z80[10]
port 291 nsew signal input
rlabel metal3 s 39200 165656 40000 165776 6 io_out_z80[11]
port 292 nsew signal input
rlabel metal3 s 39200 167016 40000 167136 6 io_out_z80[12]
port 293 nsew signal input
rlabel metal3 s 39200 168376 40000 168496 6 io_out_z80[13]
port 294 nsew signal input
rlabel metal3 s 39200 169736 40000 169856 6 io_out_z80[14]
port 295 nsew signal input
rlabel metal3 s 39200 171096 40000 171216 6 io_out_z80[15]
port 296 nsew signal input
rlabel metal3 s 39200 172456 40000 172576 6 io_out_z80[16]
port 297 nsew signal input
rlabel metal3 s 39200 173816 40000 173936 6 io_out_z80[17]
port 298 nsew signal input
rlabel metal3 s 39200 175176 40000 175296 6 io_out_z80[18]
port 299 nsew signal input
rlabel metal3 s 39200 176536 40000 176656 6 io_out_z80[19]
port 300 nsew signal input
rlabel metal3 s 39200 152056 40000 152176 6 io_out_z80[1]
port 301 nsew signal input
rlabel metal3 s 39200 177896 40000 178016 6 io_out_z80[20]
port 302 nsew signal input
rlabel metal3 s 39200 179256 40000 179376 6 io_out_z80[21]
port 303 nsew signal input
rlabel metal3 s 39200 180616 40000 180736 6 io_out_z80[22]
port 304 nsew signal input
rlabel metal3 s 39200 181976 40000 182096 6 io_out_z80[23]
port 305 nsew signal input
rlabel metal3 s 39200 183336 40000 183456 6 io_out_z80[24]
port 306 nsew signal input
rlabel metal3 s 39200 184696 40000 184816 6 io_out_z80[25]
port 307 nsew signal input
rlabel metal3 s 39200 186056 40000 186176 6 io_out_z80[26]
port 308 nsew signal input
rlabel metal3 s 39200 187416 40000 187536 6 io_out_z80[27]
port 309 nsew signal input
rlabel metal3 s 39200 188776 40000 188896 6 io_out_z80[28]
port 310 nsew signal input
rlabel metal3 s 39200 190136 40000 190256 6 io_out_z80[29]
port 311 nsew signal input
rlabel metal3 s 39200 153416 40000 153536 6 io_out_z80[2]
port 312 nsew signal input
rlabel metal3 s 39200 191496 40000 191616 6 io_out_z80[30]
port 313 nsew signal input
rlabel metal3 s 39200 192856 40000 192976 6 io_out_z80[31]
port 314 nsew signal input
rlabel metal3 s 39200 194216 40000 194336 6 io_out_z80[32]
port 315 nsew signal input
rlabel metal3 s 39200 195576 40000 195696 6 io_out_z80[33]
port 316 nsew signal input
rlabel metal3 s 39200 196936 40000 197056 6 io_out_z80[34]
port 317 nsew signal input
rlabel metal3 s 39200 198296 40000 198416 6 io_out_z80[35]
port 318 nsew signal input
rlabel metal3 s 39200 154776 40000 154896 6 io_out_z80[3]
port 319 nsew signal input
rlabel metal3 s 39200 156136 40000 156256 6 io_out_z80[4]
port 320 nsew signal input
rlabel metal3 s 39200 157496 40000 157616 6 io_out_z80[5]
port 321 nsew signal input
rlabel metal3 s 39200 158856 40000 158976 6 io_out_z80[6]
port 322 nsew signal input
rlabel metal3 s 39200 160216 40000 160336 6 io_out_z80[7]
port 323 nsew signal input
rlabel metal3 s 39200 161576 40000 161696 6 io_out_z80[8]
port 324 nsew signal input
rlabel metal3 s 39200 162936 40000 163056 6 io_out_z80[9]
port 325 nsew signal input
rlabel metal3 s 39200 96296 40000 96416 6 la_data_out[0]
port 326 nsew signal output
rlabel metal3 s 39200 109896 40000 110016 6 la_data_out[10]
port 327 nsew signal output
rlabel metal3 s 39200 111256 40000 111376 6 la_data_out[11]
port 328 nsew signal output
rlabel metal3 s 39200 112616 40000 112736 6 la_data_out[12]
port 329 nsew signal output
rlabel metal3 s 39200 113976 40000 114096 6 la_data_out[13]
port 330 nsew signal output
rlabel metal3 s 39200 115336 40000 115456 6 la_data_out[14]
port 331 nsew signal output
rlabel metal3 s 39200 116696 40000 116816 6 la_data_out[15]
port 332 nsew signal output
rlabel metal3 s 39200 118056 40000 118176 6 la_data_out[16]
port 333 nsew signal output
rlabel metal3 s 39200 119416 40000 119536 6 la_data_out[17]
port 334 nsew signal output
rlabel metal3 s 39200 120776 40000 120896 6 la_data_out[18]
port 335 nsew signal output
rlabel metal3 s 39200 122136 40000 122256 6 la_data_out[19]
port 336 nsew signal output
rlabel metal3 s 39200 97656 40000 97776 6 la_data_out[1]
port 337 nsew signal output
rlabel metal3 s 39200 123496 40000 123616 6 la_data_out[20]
port 338 nsew signal output
rlabel metal3 s 39200 124856 40000 124976 6 la_data_out[21]
port 339 nsew signal output
rlabel metal3 s 39200 126216 40000 126336 6 la_data_out[22]
port 340 nsew signal output
rlabel metal3 s 39200 127576 40000 127696 6 la_data_out[23]
port 341 nsew signal output
rlabel metal3 s 39200 128936 40000 129056 6 la_data_out[24]
port 342 nsew signal output
rlabel metal3 s 39200 130296 40000 130416 6 la_data_out[25]
port 343 nsew signal output
rlabel metal3 s 39200 131656 40000 131776 6 la_data_out[26]
port 344 nsew signal output
rlabel metal3 s 39200 133016 40000 133136 6 la_data_out[27]
port 345 nsew signal output
rlabel metal3 s 39200 134376 40000 134496 6 la_data_out[28]
port 346 nsew signal output
rlabel metal3 s 39200 135736 40000 135856 6 la_data_out[29]
port 347 nsew signal output
rlabel metal3 s 39200 99016 40000 99136 6 la_data_out[2]
port 348 nsew signal output
rlabel metal3 s 39200 137096 40000 137216 6 la_data_out[30]
port 349 nsew signal output
rlabel metal3 s 39200 138456 40000 138576 6 la_data_out[31]
port 350 nsew signal output
rlabel metal3 s 39200 139816 40000 139936 6 la_data_out[32]
port 351 nsew signal output
rlabel metal3 s 39200 141176 40000 141296 6 la_data_out[33]
port 352 nsew signal output
rlabel metal3 s 39200 142536 40000 142656 6 la_data_out[34]
port 353 nsew signal output
rlabel metal3 s 39200 143896 40000 144016 6 la_data_out[35]
port 354 nsew signal output
rlabel metal3 s 39200 145256 40000 145376 6 la_data_out[36]
port 355 nsew signal output
rlabel metal3 s 39200 146616 40000 146736 6 la_data_out[37]
port 356 nsew signal output
rlabel metal3 s 39200 147976 40000 148096 6 la_data_out[38]
port 357 nsew signal output
rlabel metal3 s 39200 149336 40000 149456 6 la_data_out[39]
port 358 nsew signal output
rlabel metal3 s 39200 100376 40000 100496 6 la_data_out[3]
port 359 nsew signal output
rlabel metal3 s 39200 101736 40000 101856 6 la_data_out[4]
port 360 nsew signal output
rlabel metal3 s 39200 103096 40000 103216 6 la_data_out[5]
port 361 nsew signal output
rlabel metal3 s 39200 104456 40000 104576 6 la_data_out[6]
port 362 nsew signal output
rlabel metal3 s 39200 105816 40000 105936 6 la_data_out[7]
port 363 nsew signal output
rlabel metal3 s 39200 107176 40000 107296 6 la_data_out[8]
port 364 nsew signal output
rlabel metal3 s 39200 108536 40000 108656 6 la_data_out[9]
port 365 nsew signal output
rlabel metal3 s 0 69368 800 69488 6 rst_scrapcpu
port 366 nsew signal output
rlabel metal2 s 1766 199200 1822 200000 6 rst_vliw
port 367 nsew signal output
rlabel metal2 s 2778 199200 2834 200000 6 rst_z80
port 368 nsew signal output
rlabel metal4 s 4208 2128 4528 197520 6 vccd1
port 369 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 197520 6 vccd1
port 369 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 197520 6 vssd1
port 370 nsew ground bidirectional
rlabel metal3 s 0 89496 800 89616 6 wb_clk_i
port 371 nsew signal input
rlabel metal3 s 0 90040 800 90160 6 wb_rst_i
port 372 nsew signal input
rlabel metal3 s 0 109624 800 109744 6 wbs_ack_o
port 373 nsew signal output
rlabel metal2 s 1398 0 1454 800 6 wbs_adr_i[0]
port 374 nsew signal input
rlabel metal2 s 13358 0 13414 800 6 wbs_adr_i[10]
port 375 nsew signal input
rlabel metal2 s 14554 0 14610 800 6 wbs_adr_i[11]
port 376 nsew signal input
rlabel metal2 s 15750 0 15806 800 6 wbs_adr_i[12]
port 377 nsew signal input
rlabel metal2 s 16946 0 17002 800 6 wbs_adr_i[13]
port 378 nsew signal input
rlabel metal2 s 18142 0 18198 800 6 wbs_adr_i[14]
port 379 nsew signal input
rlabel metal2 s 19338 0 19394 800 6 wbs_adr_i[15]
port 380 nsew signal input
rlabel metal2 s 20534 0 20590 800 6 wbs_adr_i[16]
port 381 nsew signal input
rlabel metal2 s 21730 0 21786 800 6 wbs_adr_i[17]
port 382 nsew signal input
rlabel metal2 s 22926 0 22982 800 6 wbs_adr_i[18]
port 383 nsew signal input
rlabel metal2 s 24122 0 24178 800 6 wbs_adr_i[19]
port 384 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 wbs_adr_i[1]
port 385 nsew signal input
rlabel metal2 s 25318 0 25374 800 6 wbs_adr_i[20]
port 386 nsew signal input
rlabel metal2 s 26514 0 26570 800 6 wbs_adr_i[21]
port 387 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 wbs_adr_i[22]
port 388 nsew signal input
rlabel metal2 s 28906 0 28962 800 6 wbs_adr_i[23]
port 389 nsew signal input
rlabel metal2 s 30102 0 30158 800 6 wbs_adr_i[24]
port 390 nsew signal input
rlabel metal2 s 31298 0 31354 800 6 wbs_adr_i[25]
port 391 nsew signal input
rlabel metal2 s 32494 0 32550 800 6 wbs_adr_i[26]
port 392 nsew signal input
rlabel metal2 s 33690 0 33746 800 6 wbs_adr_i[27]
port 393 nsew signal input
rlabel metal2 s 34886 0 34942 800 6 wbs_adr_i[28]
port 394 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 wbs_adr_i[29]
port 395 nsew signal input
rlabel metal2 s 3790 0 3846 800 6 wbs_adr_i[2]
port 396 nsew signal input
rlabel metal2 s 37278 0 37334 800 6 wbs_adr_i[30]
port 397 nsew signal input
rlabel metal2 s 38474 0 38530 800 6 wbs_adr_i[31]
port 398 nsew signal input
rlabel metal2 s 4986 0 5042 800 6 wbs_adr_i[3]
port 399 nsew signal input
rlabel metal2 s 6182 0 6238 800 6 wbs_adr_i[4]
port 400 nsew signal input
rlabel metal2 s 7378 0 7434 800 6 wbs_adr_i[5]
port 401 nsew signal input
rlabel metal2 s 8574 0 8630 800 6 wbs_adr_i[6]
port 402 nsew signal input
rlabel metal2 s 9770 0 9826 800 6 wbs_adr_i[7]
port 403 nsew signal input
rlabel metal2 s 10966 0 11022 800 6 wbs_adr_i[8]
port 404 nsew signal input
rlabel metal2 s 12162 0 12218 800 6 wbs_adr_i[9]
port 405 nsew signal input
rlabel metal3 s 0 108536 800 108656 6 wbs_cyc_i
port 406 nsew signal input
rlabel metal3 s 0 90584 800 90704 6 wbs_dat_i[0]
port 407 nsew signal input
rlabel metal3 s 0 96024 800 96144 6 wbs_dat_i[10]
port 408 nsew signal input
rlabel metal3 s 0 96568 800 96688 6 wbs_dat_i[11]
port 409 nsew signal input
rlabel metal3 s 0 97112 800 97232 6 wbs_dat_i[12]
port 410 nsew signal input
rlabel metal3 s 0 97656 800 97776 6 wbs_dat_i[13]
port 411 nsew signal input
rlabel metal3 s 0 98200 800 98320 6 wbs_dat_i[14]
port 412 nsew signal input
rlabel metal3 s 0 98744 800 98864 6 wbs_dat_i[15]
port 413 nsew signal input
rlabel metal3 s 0 99288 800 99408 6 wbs_dat_i[16]
port 414 nsew signal input
rlabel metal3 s 0 99832 800 99952 6 wbs_dat_i[17]
port 415 nsew signal input
rlabel metal3 s 0 100376 800 100496 6 wbs_dat_i[18]
port 416 nsew signal input
rlabel metal3 s 0 100920 800 101040 6 wbs_dat_i[19]
port 417 nsew signal input
rlabel metal3 s 0 91128 800 91248 6 wbs_dat_i[1]
port 418 nsew signal input
rlabel metal3 s 0 101464 800 101584 6 wbs_dat_i[20]
port 419 nsew signal input
rlabel metal3 s 0 102008 800 102128 6 wbs_dat_i[21]
port 420 nsew signal input
rlabel metal3 s 0 102552 800 102672 6 wbs_dat_i[22]
port 421 nsew signal input
rlabel metal3 s 0 103096 800 103216 6 wbs_dat_i[23]
port 422 nsew signal input
rlabel metal3 s 0 103640 800 103760 6 wbs_dat_i[24]
port 423 nsew signal input
rlabel metal3 s 0 104184 800 104304 6 wbs_dat_i[25]
port 424 nsew signal input
rlabel metal3 s 0 104728 800 104848 6 wbs_dat_i[26]
port 425 nsew signal input
rlabel metal3 s 0 105272 800 105392 6 wbs_dat_i[27]
port 426 nsew signal input
rlabel metal3 s 0 105816 800 105936 6 wbs_dat_i[28]
port 427 nsew signal input
rlabel metal3 s 0 106360 800 106480 6 wbs_dat_i[29]
port 428 nsew signal input
rlabel metal3 s 0 91672 800 91792 6 wbs_dat_i[2]
port 429 nsew signal input
rlabel metal3 s 0 106904 800 107024 6 wbs_dat_i[30]
port 430 nsew signal input
rlabel metal3 s 0 107448 800 107568 6 wbs_dat_i[31]
port 431 nsew signal input
rlabel metal3 s 0 92216 800 92336 6 wbs_dat_i[3]
port 432 nsew signal input
rlabel metal3 s 0 92760 800 92880 6 wbs_dat_i[4]
port 433 nsew signal input
rlabel metal3 s 0 93304 800 93424 6 wbs_dat_i[5]
port 434 nsew signal input
rlabel metal3 s 0 93848 800 93968 6 wbs_dat_i[6]
port 435 nsew signal input
rlabel metal3 s 0 94392 800 94512 6 wbs_dat_i[7]
port 436 nsew signal input
rlabel metal3 s 0 94936 800 95056 6 wbs_dat_i[8]
port 437 nsew signal input
rlabel metal3 s 0 95480 800 95600 6 wbs_dat_i[9]
port 438 nsew signal input
rlabel metal3 s 39200 52776 40000 52896 6 wbs_dat_o[0]
port 439 nsew signal output
rlabel metal3 s 39200 66376 40000 66496 6 wbs_dat_o[10]
port 440 nsew signal output
rlabel metal3 s 39200 67736 40000 67856 6 wbs_dat_o[11]
port 441 nsew signal output
rlabel metal3 s 39200 69096 40000 69216 6 wbs_dat_o[12]
port 442 nsew signal output
rlabel metal3 s 39200 70456 40000 70576 6 wbs_dat_o[13]
port 443 nsew signal output
rlabel metal3 s 39200 71816 40000 71936 6 wbs_dat_o[14]
port 444 nsew signal output
rlabel metal3 s 39200 73176 40000 73296 6 wbs_dat_o[15]
port 445 nsew signal output
rlabel metal3 s 39200 74536 40000 74656 6 wbs_dat_o[16]
port 446 nsew signal output
rlabel metal3 s 39200 75896 40000 76016 6 wbs_dat_o[17]
port 447 nsew signal output
rlabel metal3 s 39200 77256 40000 77376 6 wbs_dat_o[18]
port 448 nsew signal output
rlabel metal3 s 39200 78616 40000 78736 6 wbs_dat_o[19]
port 449 nsew signal output
rlabel metal3 s 39200 54136 40000 54256 6 wbs_dat_o[1]
port 450 nsew signal output
rlabel metal3 s 39200 79976 40000 80096 6 wbs_dat_o[20]
port 451 nsew signal output
rlabel metal3 s 39200 81336 40000 81456 6 wbs_dat_o[21]
port 452 nsew signal output
rlabel metal3 s 39200 82696 40000 82816 6 wbs_dat_o[22]
port 453 nsew signal output
rlabel metal3 s 39200 84056 40000 84176 6 wbs_dat_o[23]
port 454 nsew signal output
rlabel metal3 s 39200 85416 40000 85536 6 wbs_dat_o[24]
port 455 nsew signal output
rlabel metal3 s 39200 86776 40000 86896 6 wbs_dat_o[25]
port 456 nsew signal output
rlabel metal3 s 39200 88136 40000 88256 6 wbs_dat_o[26]
port 457 nsew signal output
rlabel metal3 s 39200 89496 40000 89616 6 wbs_dat_o[27]
port 458 nsew signal output
rlabel metal3 s 39200 90856 40000 90976 6 wbs_dat_o[28]
port 459 nsew signal output
rlabel metal3 s 39200 92216 40000 92336 6 wbs_dat_o[29]
port 460 nsew signal output
rlabel metal3 s 39200 55496 40000 55616 6 wbs_dat_o[2]
port 461 nsew signal output
rlabel metal3 s 39200 93576 40000 93696 6 wbs_dat_o[30]
port 462 nsew signal output
rlabel metal3 s 39200 94936 40000 95056 6 wbs_dat_o[31]
port 463 nsew signal output
rlabel metal3 s 39200 56856 40000 56976 6 wbs_dat_o[3]
port 464 nsew signal output
rlabel metal3 s 39200 58216 40000 58336 6 wbs_dat_o[4]
port 465 nsew signal output
rlabel metal3 s 39200 59576 40000 59696 6 wbs_dat_o[5]
port 466 nsew signal output
rlabel metal3 s 39200 60936 40000 61056 6 wbs_dat_o[6]
port 467 nsew signal output
rlabel metal3 s 39200 62296 40000 62416 6 wbs_dat_o[7]
port 468 nsew signal output
rlabel metal3 s 39200 63656 40000 63776 6 wbs_dat_o[8]
port 469 nsew signal output
rlabel metal3 s 39200 65016 40000 65136 6 wbs_dat_o[9]
port 470 nsew signal output
rlabel metal3 s 0 109080 800 109200 6 wbs_stb_i
port 471 nsew signal input
rlabel metal3 s 0 107992 800 108112 6 wbs_we_i
port 472 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 40000 200000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 6242796
string GDS_FILE /media/lucah/8a6b8802-051e-45a8-8492-771202e4c08a/ci2406-rej-pommedeterrible-tholin/openlane/Multiplexer/runs/24_05_29_14_23/results/signoff/multiplexer.magic.gds
string GDS_START 405032
<< end >>

