* NGSPICE file created from ci2406_z80.ext - technology: sky130B

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_4 abstract view
.subckt sky130_fd_sc_hd__a311o_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_4 abstract view
.subckt sky130_fd_sc_hd__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_2 abstract view
.subckt sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_1 abstract view
.subckt sky130_fd_sc_hd__o41ai_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_4 abstract view
.subckt sky130_fd_sc_hd__and2b_4 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_2 abstract view
.subckt sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_2 abstract view
.subckt sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

.subckt ci2406_z80 custom_settings[0] custom_settings[1] custom_settings[2] custom_settings[3]
+ custom_settings[4] io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15]
+ io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22] io_in[23]
+ io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30] io_in[31]
+ io_in[32] io_in[33] io_in[34] io_in[35] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14]
+ io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21]
+ io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29]
+ io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[3]
+ io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9] io_out[0] io_out[10]
+ io_out[11] io_out[12] io_out[13] io_out[14] io_out[15] io_out[16] io_out[17] io_out[18]
+ io_out[19] io_out[1] io_out[20] io_out[21] io_out[22] io_out[23] io_out[24] io_out[25]
+ io_out[26] io_out[27] io_out[28] io_out[29] io_out[2] io_out[30] io_out[31] io_out[32]
+ io_out[33] io_out[34] io_out[35] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ io_out[8] io_out[9] rst_n vccd1 vssd1 wb_clk_i
XFILLER_0_94_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3676__C1 _5387_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3155_ _3414_/B _3161_/B vssd1 vssd1 vccd1 vccd1 _4360_/B sky130_fd_sc_hd__nor2_1
X_3086_ _6458_/Q vssd1 vssd1 vccd1 vccd1 _5411_/B sky130_fd_sc_hd__inv_2
XFILLER_0_27_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3988_ _4223_/A _3987_/B _3987_/Y _3759_/Y vssd1 vssd1 vccd1 vccd1 _3988_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_91_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5727_ _4300_/A _3083_/A _5611_/Y _5726_/X vssd1 vssd1 vccd1 vccd1 _5727_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_45_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5658_ _5732_/A _5656_/X _5657_/X _5655_/X vssd1 vssd1 vccd1 vccd1 _5658_/X sky130_fd_sc_hd__o31a_1
XFILLER_0_32_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5589_ hold531/X _5588_/X _6070_/A vssd1 vssd1 vccd1 vccd1 _5589_/X sky130_fd_sc_hd__mux2_1
X_4609_ hold417/X _4604_/X _4605_/X hold444/X _4608_/X vssd1 vssd1 vccd1 vccd1 _4609_/X
+ sky130_fd_sc_hd__a221o_1
Xhold340 _6319_/Q vssd1 vssd1 vccd1 vccd1 hold340/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold362 _5758_/X vssd1 vssd1 vccd1 vccd1 _6402_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold351 _6322_/Q vssd1 vssd1 vccd1 vccd1 hold351/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold395 _6121_/Q vssd1 vssd1 vccd1 vccd1 _4296_/A sky130_fd_sc_hd__buf_1
Xhold373 _6369_/Q vssd1 vssd1 vccd1 vccd1 _5521_/A sky130_fd_sc_hd__buf_1
Xhold384 _4958_/X vssd1 vssd1 vccd1 vccd1 _6324_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5440__S _5593_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold639_A _6314_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4631__A1 _4131_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5895__B1 _5771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3122__A1 _3530_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4870__B2 _4863_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4960_ _6259_/Q _6218_/Q _6194_/Q _6111_/Q _5100_/S1 _5100_/S0 vssd1 vssd1 vccd1
+ vccd1 _4960_/X sky130_fd_sc_hd__mux4_1
XANTENNA__4622__B2 _6312_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4622__A1 _6461_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_48_wb_clk_i_A clkbuf_leaf_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_3911_ _3904_/X _3905_/X _3910_/X _4441_/S vssd1 vssd1 vccd1 vccd1 _3911_/X sky130_fd_sc_hd__a22o_2
X_4891_ _4885_/X _4888_/X _4889_/X _4890_/X vssd1 vssd1 vccd1 vccd1 _4891_/X sky130_fd_sc_hd__o31a_1
XFILLER_0_13_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3842_ _6174_/Q _6253_/Q _3865_/S vssd1 vssd1 vccd1 vccd1 _3842_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_27_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3773_ _3774_/A _3774_/B vssd1 vssd1 vccd1 vccd1 _3773_/Y sky130_fd_sc_hd__nor2_2
X_5512_ _6465_/Q _5511_/X _5512_/S vssd1 vssd1 vccd1 vccd1 _5512_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_13_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3537__C _5314_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4689__A1 _4713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5443_ _5443_/A _5443_/B vssd1 vssd1 vccd1 vccd1 _5445_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_42_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5374_ _6432_/Q _5374_/B _5374_/C vssd1 vssd1 vccd1 vccd1 _5374_/X sky130_fd_sc_hd__and3_1
X_4325_ _4325_/A _5387_/B _4325_/C vssd1 vssd1 vccd1 vccd1 _5605_/D sky130_fd_sc_hd__nor3_2
Xfanout105 _4263_/A vssd1 vssd1 vccd1 vccd1 _5146_/C sky130_fd_sc_hd__clkbuf_8
Xfanout127 _4300_/A vssd1 vssd1 vccd1 vccd1 _4715_/B2 sky130_fd_sc_hd__buf_4
Xfanout116 _5581_/S vssd1 vssd1 vccd1 vccd1 _5489_/S sky130_fd_sc_hd__buf_4
XFILLER_0_1_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout138 _5404_/A0 vssd1 vssd1 vccd1 vccd1 _5100_/S0 sky130_fd_sc_hd__buf_6
Xfanout149 _6297_/Q vssd1 vssd1 vccd1 vccd1 _4268_/A sky130_fd_sc_hd__buf_4
X_4256_ _5388_/A _4253_/Y _5388_/C _3511_/A vssd1 vssd1 vccd1 vccd1 _4256_/X sky130_fd_sc_hd__o31a_1
XANTENNA__4310__A0 _6313_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3207_ _3204_/X _3206_/Y _4273_/A _3326_/B vssd1 vssd1 vccd1 vccd1 _3221_/B sky130_fd_sc_hd__a211o_1
X_4187_ _6225_/Q _3804_/X _3807_/X _6141_/Q vssd1 vssd1 vccd1 vccd1 _4187_/X sky130_fd_sc_hd__a22o_1
X_3138_ _4268_/A _4273_/A _4248_/B vssd1 vssd1 vccd1 vccd1 _4357_/C sky130_fd_sc_hd__and3_1
XANTENNA__3664__A2 _6019_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3069_ _3480_/B vssd1 vssd1 vccd1 vccd1 _3785_/B sky130_fd_sc_hd__inv_2
XFILLER_0_77_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4613__A1 _6459_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4613__B2 _6310_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3744__A _6284_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold491_A _6436_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold170 _6010_/X vssd1 vssd1 vccd1 vccd1 _6455_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold192 _6133_/Q vssd1 vssd1 vccd1 vccd1 hold192/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold181 _6147_/Q vssd1 vssd1 vccd1 vccd1 hold181/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4301__A0 _6311_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3355__A_N _5600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4514__S _4518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3357__C _5315_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3343__A1 _6431_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4110_ _4162_/A _4210_/A _6334_/Q vssd1 vssd1 vccd1 vccd1 _4111_/B sky130_fd_sc_hd__mux2_1
XANTENNA__5096__A1 _5771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5090_ _5109_/A1 _5085_/X _5089_/X _4924_/C vssd1 vssd1 vccd1 vccd1 _5090_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_75_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4041_ hold147/X hold173/X hold165/X hold73/X _5721_/C1 _5721_/B1 vssd1 vssd1 vccd1
+ vccd1 _4041_/X sky130_fd_sc_hd__mux4_2
XANTENNA__5080__S _5101_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5992_ _3636_/C _3635_/Y _5991_/X _3636_/B hold472/X vssd1 vssd1 vccd1 vccd1 _5992_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA_clkbuf_leaf_4_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_59_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4943_ _6365_/Q _6366_/Q _6367_/Q _6368_/Q vssd1 vssd1 vccd1 vccd1 _4945_/A sky130_fd_sc_hd__and4_1
XFILLER_0_24_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4874_ _6364_/Q _5861_/S _5842_/B1 _4873_/X vssd1 vssd1 vccd1 vccd1 _4874_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_74_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3825_ hold51/A hold53/A _3865_/S vssd1 vssd1 vccd1 vccd1 _3825_/X sky130_fd_sc_hd__mux2_1
X_3756_ _5136_/A _6284_/Q _6378_/Q _4060_/B _3755_/X vssd1 vssd1 vccd1 vccd1 _5162_/A
+ sky130_fd_sc_hd__o41a_1
XANTENNA_fanout125_A _4715_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6475_ _6475_/CLK _6475_/D fanout175/X vssd1 vssd1 vccd1 vccd1 _6475_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_0_42_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3687_ _3682_/X _3684_/Y _4262_/B _3681_/X _5146_/C vssd1 vssd1 vccd1 vccd1 _3687_/X
+ sky130_fd_sc_hd__a32o_1
X_5426_ _5607_/B2 _3789_/X _3790_/X _3788_/Y _5478_/S vssd1 vssd1 vccd1 vccd1 _5492_/A
+ sky130_fd_sc_hd__a311o_4
X_5357_ _5600_/A _4249_/A _5356_/Y _4289_/C vssd1 vssd1 vccd1 vccd1 _5357_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_10_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5288_ _6340_/Q _6282_/Q _5288_/S vssd1 vssd1 vccd1 vccd1 _5288_/X sky130_fd_sc_hd__mux2_1
X_4308_ _5581_/S _4312_/A _4307_/X vssd1 vssd1 vccd1 vccd1 _4308_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_4_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4239_ _5732_/A _4236_/X _4237_/X _4238_/X vssd1 vssd1 vccd1 vccd1 _4239_/X sky130_fd_sc_hd__o31a_1
XANTENNA__3637__A2 _3506_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold504_A _6331_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4770__A0 _4227_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4289__B _4289_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4509__S _4509_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4825__B2 _6459_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3610_ _3610_/A _5523_/A vssd1 vssd1 vccd1 vccd1 _3611_/C sky130_fd_sc_hd__nor2_1
X_4590_ _4276_/A _4588_/X _4589_/Y _3205_/B vssd1 vssd1 vccd1 vccd1 _4590_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_9_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3541_ _3307_/A _3541_/B _3541_/C vssd1 vssd1 vccd1 vccd1 _3541_/X sky130_fd_sc_hd__and3b_1
XFILLER_0_24_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5075__S _5974_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3472_ _3530_/A _3472_/B vssd1 vssd1 vccd1 vccd1 _3487_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_51_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6260_ _6490_/CLK _6260_/D vssd1 vssd1 vccd1 vccd1 _6260_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5211_ _6465_/Q _6464_/Q vssd1 vssd1 vccd1 vccd1 _5213_/A sky130_fd_sc_hd__xor2_1
X_6191_ _6454_/CLK _6191_/D vssd1 vssd1 vccd1 vccd1 _6191_/Q sky130_fd_sc_hd__dfxtp_1
X_5142_ _3773_/Y _4203_/A _5138_/X _3774_/A _5141_/X vssd1 vssd1 vccd1 vccd1 _5142_/X
+ sky130_fd_sc_hd__a221o_1
X_5073_ _6374_/Q _5848_/S _5972_/B1 _5072_/X vssd1 vssd1 vccd1 vccd1 _5073_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_79_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4024_ _6381_/Q _4021_/X _4022_/X _3759_/Y _4020_/X vssd1 vssd1 vccd1 vccd1 _4024_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3550__C _5388_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6018__A0 input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4943__A _6365_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4662__B _4668_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5975_ _5974_/X _5969_/A _5975_/S vssd1 vssd1 vccd1 vccd1 _5975_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_47_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4926_ _4920_/B _4925_/X _4948_/S vssd1 vssd1 vccd1 vccd1 _4926_/X sky130_fd_sc_hd__mux2_1
X_4857_ _4361_/B _4844_/X _4776_/Y vssd1 vssd1 vccd1 vccd1 _4857_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_51_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3808_ _3884_/S _3811_/B vssd1 vssd1 vccd1 vccd1 _4400_/A sky130_fd_sc_hd__nand2_2
XANTENNA__4347__A3 _5388_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4788_ _6447_/Q _4788_/B vssd1 vssd1 vccd1 vccd1 _4789_/B sky130_fd_sc_hd__and2_2
XANTENNA__3555__B2 _4324_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3555__A1 _4363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6527_ _6529_/A vssd1 vssd1 vccd1 vccd1 _6527_/X sky130_fd_sc_hd__buf_1
XFILLER_0_15_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3294__A _5315_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3739_ _6346_/Q _5247_/S vssd1 vssd1 vccd1 vccd1 _3979_/A sky130_fd_sc_hd__nand2_4
X_6458_ _6465_/CLK _6458_/D fanout181/X vssd1 vssd1 vccd1 vccd1 _6458_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6101__C _6101_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5409_ _6430_/Q _4289_/C _5405_/Y _5408_/X _5600_/A vssd1 vssd1 vccd1 vccd1 _5410_/B
+ sky130_fd_sc_hd__a32o_1
X_6389_ _6452_/CLK hold34/X vssd1 vssd1 vccd1 vccd1 hold33/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3741__B _6378_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6257__RESET_B fanout181/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4556__C _4556_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5014__A _6460_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3460__C _5478_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5480__A1 _5492_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold621_A _6462_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5387__C _5387_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3849__A2 _3884_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5471__A1 _6365_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5760_ _6311_/Q hold403/X _5765_/S vssd1 vssd1 vccd1 vccd1 _5760_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_29_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4711_ _6385_/Q _6381_/Q _4711_/S vssd1 vssd1 vccd1 vccd1 _4711_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5691_ _6453_/Q _5721_/A2 _5721_/B1 _6230_/Q _5730_/C1 vssd1 vssd1 vccd1 vccd1 _5693_/A
+ sky130_fd_sc_hd__o221a_1
XANTENNA__4702__S _4711_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4642_ _4190_/B _4611_/B _4602_/Y _4641_/X vssd1 vssd1 vccd1 vccd1 _4642_/X sky130_fd_sc_hd__o211a_1
XANTENNA__5526__A2 _5485_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4573_ hold485/X _6338_/Q _4575_/S vssd1 vssd1 vccd1 vccd1 _4573_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_4_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4003__A _4150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3524_ _3570_/B _3410_/Y _3521_/Y _3522_/X _3541_/C vssd1 vssd1 vccd1 vccd1 _3524_/X
+ sky130_fd_sc_hd__o41a_1
X_6312_ _6312_/CLK _6312_/D fanout182/X vssd1 vssd1 vccd1 vccd1 _6312_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_0_4_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3455_ _5617_/A _3405_/B _3452_/Y vssd1 vssd1 vccd1 vccd1 _3456_/D sky130_fd_sc_hd__o21ai_1
X_6243_ _6439_/CLK hold40/X fanout177/X vssd1 vssd1 vccd1 vccd1 hold39/A sky130_fd_sc_hd__dfrtp_1
XANTENNA__3561__B _3619_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3386_ _3386_/A _4802_/D vssd1 vssd1 vccd1 vccd1 _3386_/Y sky130_fd_sc_hd__nand2_1
X_6174_ _6454_/CLK _6174_/D vssd1 vssd1 vccd1 vccd1 _6174_/Q sky130_fd_sc_hd__dfxtp_1
X_5125_ _5244_/S vssd1 vssd1 vccd1 vccd1 _5125_/Y sky130_fd_sc_hd__inv_2
XANTENNA__6350__RESET_B fanout176/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5056_ hold359/X _5055_/X _6070_/A vssd1 vssd1 vccd1 vccd1 _5056_/X sky130_fd_sc_hd__mux2_1
X_4007_ _4007_/A _4007_/B vssd1 vssd1 vccd1 vccd1 _4007_/X sky130_fd_sc_hd__or2_1
XANTENNA__4673__A _6076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5958_ _6427_/Q _5970_/A vssd1 vssd1 vccd1 vccd1 _5959_/B sky130_fd_sc_hd__nor2_1
XANTENNA__4422__C1 _5730_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4909_ _4905_/Y _4907_/X _4908_/X _4906_/X vssd1 vssd1 vccd1 vccd1 _4909_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_47_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5889_ _6421_/Q _5970_/A vssd1 vssd1 vccd1 vccd1 _5889_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_90_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3528__B2 _5398_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5951__B _5970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold41 hold41/A vssd1 vssd1 vccd1 vccd1 hold41/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold30 hold30/A vssd1 vssd1 vccd1 vccd1 hold30/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold63 hold63/A vssd1 vssd1 vccd1 vccd1 hold63/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 hold74/A vssd1 vssd1 vccd1 vccd1 hold74/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold52 hold52/A vssd1 vssd1 vccd1 vccd1 hold52/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold96 hold96/A vssd1 vssd1 vccd1 vccd1 hold96/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 hold85/A vssd1 vssd1 vccd1 vccd1 hold85/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_85_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3767__A1 _4716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4522__S _4527_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_14_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6474_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_5 _5411_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3240_ _3627_/B _3240_/B vssd1 vssd1 vccd1 vccd1 _3240_/X sky130_fd_sc_hd__and2_1
XFILLER_0_67_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3171_ _4273_/A _4784_/B _3609_/A _5346_/A vssd1 vssd1 vccd1 vccd1 _3186_/B sky130_fd_sc_hd__a211o_1
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4924__C _4924_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3207__B1 _4273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5812_ _5813_/A _5813_/B _5811_/X vssd1 vssd1 vccd1 vccd1 _5826_/B sky130_fd_sc_hd__o21ba_1
XFILLER_0_9_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5743_ hold29/X _3892_/B _5769_/S vssd1 vssd1 vccd1 vccd1 hold30/A sky130_fd_sc_hd__mux2_1
XFILLER_0_29_297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5674_ _5674_/A _5674_/B _5674_/C vssd1 vssd1 vccd1 vccd1 _5674_/X sky130_fd_sc_hd__or3_1
XANTENNA__4707__A0 _6384_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4625_ _5757_/B hold470/X _4582_/Y _4624_/X vssd1 vssd1 vccd1 vccd1 _4625_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_32_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4556_ _6159_/Q _5489_/S _4556_/C _4957_/S vssd1 vssd1 vccd1 vccd1 _4575_/S sky130_fd_sc_hd__and4_4
Xhold511 _4571_/X vssd1 vssd1 vccd1 vccd1 _6278_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold500 _6353_/Q vssd1 vssd1 vccd1 vccd1 _4670_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5380__B1 _6021_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold544 _3646_/X vssd1 vssd1 vccd1 vccd1 _3647_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3507_ _3699_/A _3527_/B vssd1 vssd1 vccd1 vccd1 _3638_/B sky130_fd_sc_hd__and2_1
XANTENNA__5771__B _5771_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold533 _6373_/Q vssd1 vssd1 vccd1 vccd1 _5567_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold522 _6486_/Q vssd1 vssd1 vccd1 vccd1 hold522/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4668__A _4668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold577 _6437_/Q vssd1 vssd1 vccd1 vccd1 _5995_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold566 _6431_/Q vssd1 vssd1 vccd1 vccd1 hold566/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold555 _5675_/X vssd1 vssd1 vccd1 vccd1 _6380_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4487_ _4042_/X hold147/X _4491_/S vssd1 vssd1 vccd1 vccd1 _4487_/X sky130_fd_sc_hd__mux2_1
Xhold588 _6421_/Q vssd1 vssd1 vccd1 vccd1 hold588/X sky130_fd_sc_hd__dlygate4sd3_1
X_3438_ _4358_/B _5369_/D vssd1 vssd1 vccd1 vccd1 _3456_/B sky130_fd_sc_hd__or2_1
Xhold599 _6130_/Q vssd1 vssd1 vccd1 vccd1 hold599/X sky130_fd_sc_hd__dlygate4sd3_1
X_6226_ _6449_/CLK _6226_/D vssd1 vssd1 vccd1 vccd1 _6226_/Q sky130_fd_sc_hd__dfxtp_1
X_3369_ _6339_/Q _4720_/C _3367_/X _3986_/A vssd1 vssd1 vccd1 vccd1 _3370_/C sky130_fd_sc_hd__a211o_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6157_ _6263_/CLK _6157_/D vssd1 vssd1 vccd1 vccd1 _6157_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5108_ _6465_/Q _5107_/X _5108_/S vssd1 vssd1 vccd1 vccd1 _5108_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5435__A1 _4656_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6088_ _6101_/A _6087_/X _6107_/S vssd1 vssd1 vccd1 vccd1 _6088_/X sky130_fd_sc_hd__o21a_1
X_5039_ _6263_/Q _6198_/Q _6222_/Q _6115_/Q _5100_/S0 _5078_/S1 vssd1 vssd1 vccd1
+ vccd1 _5039_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_95_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5438__S _5489_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4410__A2 _4406_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput42 _6304_/Q vssd1 vssd1 vccd1 vccd1 io_out[23] sky130_fd_sc_hd__buf_12
Xoutput20 _6524_/X vssd1 vssd1 vccd1 vccd1 io_oeb[23] sky130_fd_sc_hd__buf_12
Xoutput31 _6324_/Q vssd1 vssd1 vccd1 vccd1 io_out[13] sky130_fd_sc_hd__buf_12
Xoutput53 _6163_/Q vssd1 vssd1 vccd1 vccd1 io_out[3] sky130_fd_sc_hd__buf_12
XANTENNA__3632__D _3632_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5426__A1 _5607_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4517__S _4518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_38_wb_clk_i_A clkbuf_leaf_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_85_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4410_ _6450_/Q _4406_/B _4420_/S _6227_/Q _5730_/C1 vssd1 vssd1 vccd1 vccd1 _4410_/X
+ sky130_fd_sc_hd__o221a_1
X_5390_ _4261_/Y _4264_/X _5364_/C _5607_/B2 vssd1 vssd1 vccd1 vccd1 _5391_/C sky130_fd_sc_hd__o31a_1
XFILLER_0_1_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3392__A _3497_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4341_ _5607_/B2 _4329_/X _4340_/X vssd1 vssd1 vccd1 vccd1 _4341_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4272_ _4675_/A _3570_/B _4264_/C _4271_/X vssd1 vssd1 vccd1 vccd1 _4272_/X sky130_fd_sc_hd__a31o_1
XANTENNA__5114__A0 _6465_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3223_ _4359_/C _3205_/X _3222_/X _3639_/D vssd1 vssd1 vccd1 vccd1 _3235_/B sky130_fd_sc_hd__o2bb2a_1
X_6011_ _4463_/X hold300/X _6011_/S vssd1 vssd1 vccd1 vccd1 _6456_/D sky130_fd_sc_hd__mux2_1
XANTENNA__5665__A1 _6460_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4000__B _6381_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3676__B1 _5777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3154_ _3326_/B _3360_/B vssd1 vssd1 vccd1 vccd1 _3161_/B sky130_fd_sc_hd__or2_1
X_3085_ _6459_/Q vssd1 vssd1 vccd1 vccd1 _5427_/B sky130_fd_sc_hd__inv_2
XANTENNA__6090__A1 _4366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout155_A _3284_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3987_ _4168_/B _3987_/B vssd1 vssd1 vccd1 vccd1 _3987_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_9_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5726_ _5726_/A _5726_/B _5726_/C vssd1 vssd1 vccd1 vccd1 _5726_/X sky130_fd_sc_hd__or3_1
XANTENNA__3286__B _3489_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5657_ _6135_/Q _4406_/B _4235_/S _6179_/Q _5731_/C1 vssd1 vssd1 vccd1 vccd1 _5657_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_60_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5588_ hold531/X _5520_/B _5587_/X _5415_/X vssd1 vssd1 vccd1 vccd1 _5588_/X sky130_fd_sc_hd__a22o_1
X_4608_ _6458_/Q _4606_/X _4607_/X _6309_/Q _4603_/X vssd1 vssd1 vccd1 vccd1 _4608_/X
+ sky130_fd_sc_hd__a221o_1
Xhold330 _6308_/Q vssd1 vssd1 vccd1 vccd1 hold330/X sky130_fd_sc_hd__dlygate4sd3_1
X_4539_ hold79/X _4416_/X _4545_/S vssd1 vssd1 vccd1 vccd1 hold80/A sky130_fd_sc_hd__mux2_1
Xhold341 _4860_/X vssd1 vssd1 vccd1 vccd1 _6319_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold352 _4916_/X vssd1 vssd1 vccd1 vccd1 _6322_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold385 _6466_/Q vssd1 vssd1 vccd1 vccd1 _6025_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold396 _4299_/X vssd1 vssd1 vccd1 vccd1 _6121_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold363 _6485_/Q vssd1 vssd1 vccd1 vccd1 hold363/X sky130_fd_sc_hd__buf_1
Xhold374 _5528_/X vssd1 vssd1 vccd1 vccd1 _6369_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6209_ _6456_/CLK _6209_/D vssd1 vssd1 vccd1 vccd1 _6209_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3667__B1 _5146_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout68_A _5816_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5019__S0 _5100_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3627__D _3674_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4800__S _4800_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4101__A _6289_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3122__A2 _3497_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output49_A _3656_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6072__B2 _4366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4083__B1 _4463_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3910_ hold276/X hold220/X hold163/X hold109/X _4235_/S _5721_/C1 vssd1 vssd1 vccd1
+ vccd1 _3910_/X sky130_fd_sc_hd__mux4_2
X_4890_ _6417_/Q _4930_/B vssd1 vssd1 vccd1 vccd1 _4890_/X sky130_fd_sc_hd__or2_1
X_3841_ hold85/A _6190_/Q _3865_/S vssd1 vssd1 vccd1 vccd1 _3841_/X sky130_fd_sc_hd__mux2_1
X_3772_ _6345_/Q _3772_/B vssd1 vssd1 vccd1 vccd1 _3774_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_13_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3818__C _3818_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5511_ _5509_/Y _5510_/X _5567_/B vssd1 vssd1 vccd1 vccd1 _5511_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_42_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5442_ _5492_/A _5441_/B _5441_/C vssd1 vssd1 vccd1 vccd1 _5443_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__4138__B2 _4441_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5373_ _5373_/A _5373_/B vssd1 vssd1 vccd1 vccd1 _5376_/S sky130_fd_sc_hd__nor2_1
X_4324_ _4324_/A _4324_/B vssd1 vssd1 vccd1 vccd1 _4324_/X sky130_fd_sc_hd__or2_1
Xfanout128 hold526/X vssd1 vssd1 vccd1 vccd1 _4300_/A sky130_fd_sc_hd__buf_4
Xfanout106 _3276_/Y vssd1 vssd1 vccd1 vccd1 _5607_/B2 sky130_fd_sc_hd__buf_6
Xfanout117 _6108_/S vssd1 vssd1 vccd1 vccd1 _5581_/S sky130_fd_sc_hd__buf_4
XANTENNA__5638__A1 _5655_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4255_ _4255_/A vssd1 vssd1 vccd1 vccd1 _5388_/C sky130_fd_sc_hd__inv_2
Xfanout139 hold644/X vssd1 vssd1 vccd1 vccd1 _5404_/A0 sky130_fd_sc_hd__buf_8
XFILLER_0_10_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3206_ _3547_/B _3176_/Y _3205_/X vssd1 vssd1 vccd1 vccd1 _3206_/Y sky130_fd_sc_hd__a21oi_1
X_4186_ _6266_/Q _3793_/X _3795_/X _6201_/Q _4185_/X vssd1 vssd1 vccd1 vccd1 _4189_/A
+ sky130_fd_sc_hd__a221o_1
X_3137_ _3414_/B vssd1 vssd1 vccd1 vccd1 _4359_/B sky130_fd_sc_hd__inv_2
XFILLER_0_89_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5777__A _5777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3068_ _3501_/A vssd1 vssd1 vccd1 vccd1 _5295_/A sky130_fd_sc_hd__inv_4
XANTENNA__5810__A1 _5867_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4681__A _6081_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3821__B1 _3810_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3585__C1 _5605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5709_ _5709_/A _5709_/B vssd1 vssd1 vccd1 vccd1 _5709_/X sky130_fd_sc_hd__or2_1
XFILLER_0_18_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold160 _4503_/X vssd1 vssd1 vccd1 vccd1 _6211_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold171 _6203_/Q vssd1 vssd1 vccd1 vccd1 hold171/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold193 _3542_/X vssd1 vssd1 vccd1 vccd1 _6133_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold182 _4383_/X vssd1 vssd1 vccd1 vccd1 _6147_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5801__A1 _5867_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3935__A _6287_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4530__S _4536_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3670__A _4268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4040_ hold15/X _4462_/A2 _4463_/S vssd1 vssd1 vccd1 vccd1 _4040_/X sky130_fd_sc_hd__o21a_1
XANTENNA__6045__A1 _6101_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6045__B2 _6036_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5991_ _6437_/Q _6438_/Q _5980_/Y _3489_/B _5980_/A vssd1 vssd1 vccd1 vccd1 _5991_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_86_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4942_ _5102_/A _4942_/B vssd1 vssd1 vccd1 vccd1 _4942_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_59_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6375__RESET_B fanout172/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4873_ _6364_/Q _4872_/X _5892_/S vssd1 vssd1 vccd1 vccd1 _4873_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6304__RESET_B fanout183/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3824_ _6208_/Q _3793_/X _3795_/X hold89/A vssd1 vssd1 vccd1 vccd1 _3830_/A sky130_fd_sc_hd__a22o_1
X_3755_ _3749_/X _3750_/Y _4060_/B _3754_/X vssd1 vssd1 vccd1 vccd1 _3755_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_15_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3686_ _3682_/X _3684_/Y _4262_/B _3681_/X _5146_/C vssd1 vssd1 vccd1 vccd1 _5296_/B
+ sky130_fd_sc_hd__a32oi_4
X_6474_ _6474_/CLK _6474_/D fanout180/X vssd1 vssd1 vccd1 vccd1 _6474_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout118_A _5866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5425_ _5489_/S _5421_/X _5424_/X hold581/X vssd1 vssd1 vccd1 vccd1 _5425_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5859__B2 _5874_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5356_ _4248_/C _5360_/C _3457_/X vssd1 vssd1 vccd1 vccd1 _5356_/Y sky130_fd_sc_hd__a21oi_1
X_5287_ _6340_/Q _5202_/A _5286_/X _4216_/Y _4223_/X vssd1 vssd1 vccd1 vccd1 _5287_/X
+ sky130_fd_sc_hd__a2111o_1
X_4307_ _6312_/Q _4322_/B _4304_/X _4306_/X vssd1 vssd1 vccd1 vccd1 _4307_/X sky130_fd_sc_hd__a22o_1
X_4238_ _5730_/C1 _4235_/X _4234_/X _5655_/B vssd1 vssd1 vccd1 vccd1 _4238_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_4_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4169_ _6289_/Q _5268_/A _4716_/A vssd1 vssd1 vccd1 vccd1 _5263_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_97_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4047__B1 _3795_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4598__A1 _3172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5795__B1 _5784_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5970__A _5970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3956__S0 _5721_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_39_wb_clk_i clkbuf_leaf_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6481_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_45_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4525__S _4527_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5210__A _6459_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3540_ _3574_/B _3539_/Y _5384_/A vssd1 vssd1 vccd1 vccd1 _3540_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__4761__A1 _6315_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4761__B2 _4957_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3471_ _4800_/S _3471_/B vssd1 vssd1 vccd1 vccd1 _3472_/B sky130_fd_sc_hd__nand2_4
X_5210_ _6459_/Q _6458_/Q vssd1 vssd1 vccd1 vccd1 _5214_/A sky130_fd_sc_hd__xor2_1
X_6190_ _6456_/CLK _6190_/D vssd1 vssd1 vccd1 vccd1 _6190_/Q sky130_fd_sc_hd__dfxtp_1
X_5141_ _4115_/A _5140_/X _5290_/S hold306/X _5139_/X vssd1 vssd1 vccd1 vccd1 _5141_/X
+ sky130_fd_sc_hd__a2111o_1
X_5072_ _6407_/Q _5071_/X _5971_/S vssd1 vssd1 vccd1 vccd1 _5072_/X sky130_fd_sc_hd__mux2_1
X_4023_ _5260_/A _5175_/B _5267_/D _3770_/A vssd1 vssd1 vccd1 vccd1 _4023_/X sky130_fd_sc_hd__a2bb2o_1
XANTENNA__4816__A2 _6070_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4943__B _6366_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5974_ _6465_/Q _5973_/X _5974_/S vssd1 vssd1 vccd1 vccd1 _5974_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_19_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4925_ _6419_/Q _6367_/Q _5105_/S vssd1 vssd1 vccd1 vccd1 _4925_/X sky130_fd_sc_hd__mux2_1
X_4856_ _5817_/A _4856_/B vssd1 vssd1 vccd1 vccd1 _4856_/Y sky130_fd_sc_hd__nand2_1
X_3807_ _3852_/A _3883_/S _3884_/S vssd1 vssd1 vccd1 vccd1 _3807_/X sky130_fd_sc_hd__and3_4
XANTENNA__3575__A _5605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4787_ _5422_/B _4787_/B vssd1 vssd1 vccd1 vccd1 _5816_/S sky130_fd_sc_hd__nand2_2
X_6526_ _6529_/A vssd1 vssd1 vccd1 vccd1 _6526_/X sky130_fd_sc_hd__buf_1
XFILLER_0_15_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3738_ _6346_/Q _5247_/S vssd1 vssd1 vccd1 vccd1 _3738_/X sky130_fd_sc_hd__and2_1
XFILLER_0_15_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6334__SET_B fanout183/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3669_ _3557_/B _3668_/Y _5522_/A vssd1 vssd1 vccd1 vccd1 _3669_/Y sky130_fd_sc_hd__o21ai_2
X_6457_ _6474_/CLK _6457_/D fanout179/X vssd1 vssd1 vccd1 vccd1 _6457_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_0_30_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5408_ _3444_/Y _3522_/X _5407_/X _4335_/B vssd1 vssd1 vccd1 vccd1 _5408_/X sky130_fd_sc_hd__a22o_1
X_6388_ _6452_/CLK hold30/X vssd1 vssd1 vccd1 vccd1 hold29/A sky130_fd_sc_hd__dfxtp_1
X_5339_ _5323_/B _3420_/Y _5338_/X _5364_/B _5605_/B vssd1 vssd1 vccd1 vccd1 _5339_/X
+ sky130_fd_sc_hd__o32a_1
XANTENNA__4556__D _4957_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5014__B _5771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5949__B _5970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4853__B _4930_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4991__B2 _4924_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4991__A1 _5109_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4743__A1 _6312_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4743__B2 _4957_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3218__A_N _4273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5759__A0 _6310_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3234__A1 _5124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4710_ _4715_/B2 _4706_/Y _4709_/X hold312/X _4672_/Y vssd1 vssd1 vccd1 vccd1 _4710_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_0_29_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5690_ _6337_/Q _5628_/X _5643_/X _6425_/Q vssd1 vssd1 vccd1 vccd1 _5700_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_56_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4641_ _4641_/A _4641_/B vssd1 vssd1 vccd1 vccd1 _4641_/X sky130_fd_sc_hd__or2_1
X_4572_ hold450/X _6337_/Q _4575_/S vssd1 vssd1 vccd1 vccd1 _4572_/X sky130_fd_sc_hd__mux2_1
X_3523_ _5322_/A _5384_/A vssd1 vssd1 vccd1 vccd1 _3541_/C sky130_fd_sc_hd__nor2_2
X_6311_ _6336_/CLK _6311_/D fanout182/X vssd1 vssd1 vccd1 vccd1 _6311_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_0_12_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3454_ _4253_/A _3412_/Y _3434_/Y _3409_/Y _3453_/X vssd1 vssd1 vccd1 vccd1 _3456_/C
+ sky130_fd_sc_hd__o221ai_1
X_6242_ _6242_/CLK hold36/X fanout180/X vssd1 vssd1 vccd1 vccd1 hold35/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5695__C1 _5721_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4938__B _5101_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3385_ _4324_/B _4792_/A _3384_/X vssd1 vssd1 vccd1 vccd1 _4802_/D sky130_fd_sc_hd__or3b_4
X_6173_ _6237_/CLK _6173_/D vssd1 vssd1 vccd1 vccd1 _6173_/Q sky130_fd_sc_hd__dfxtp_1
X_5124_ _5124_/A _5322_/A _5124_/C vssd1 vssd1 vccd1 vccd1 _5244_/S sky130_fd_sc_hd__or3_4
XANTENNA_fanout185_A input18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5055_ _6462_/Q _5054_/X _5974_/S vssd1 vssd1 vccd1 vccd1 _5055_/X sky130_fd_sc_hd__mux2_1
X_4006_ _3975_/A _3975_/B _3973_/A vssd1 vssd1 vccd1 vccd1 _4007_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_27_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4673__B _4714_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_338 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3289__B _5777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5957_ _6427_/Q _5970_/A vssd1 vssd1 vccd1 vccd1 _5959_/A sky130_fd_sc_hd__and2_1
X_4908_ _6463_/Q _4963_/B _4904_/X _5109_/A1 vssd1 vssd1 vccd1 vccd1 _4908_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_90_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5888_ hold518/X _5887_/X _5977_/S vssd1 vssd1 vccd1 vccd1 _5888_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_35_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4839_ _4957_/S _4836_/X _4837_/X _4838_/X vssd1 vssd1 vccd1 vccd1 _4839_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3736__C _5314_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3104__C_N _4273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold564_A _6285_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold20 hold20/A vssd1 vssd1 vccd1 vccd1 hold20/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 hold31/A vssd1 vssd1 vccd1 vccd1 hold31/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 hold42/A vssd1 vssd1 vccd1 vccd1 hold42/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 hold64/A vssd1 vssd1 vccd1 vccd1 hold64/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 hold53/A vssd1 vssd1 vccd1 vccd1 hold53/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 hold75/A vssd1 vssd1 vccd1 vccd1 hold75/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold86 hold86/A vssd1 vssd1 vccd1 vccd1 hold86/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 hold97/A vssd1 vssd1 vccd1 vccd1 hold97/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_28_wb_clk_i_A clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_78_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4964__B2 _4962_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4104__A _6333_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_6 _6444_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3170_ _5344_/B _4556_/C vssd1 vssd1 vccd1 vccd1 _3609_/A sky130_fd_sc_hd__or2_1
XANTENNA__5692__A2 _5721_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xci2406_z80_210 vssd1 vssd1 vccd1 vccd1 ci2406_z80_210/HI io_out[4] sky130_fd_sc_hd__conb_1
XFILLER_0_88_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5811_ _5826_/A _5811_/B vssd1 vssd1 vccd1 vccd1 _5811_/X sky130_fd_sc_hd__or2_1
XFILLER_0_91_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5742_ _5742_/A vssd1 vssd1 vccd1 vccd1 _6387_/D sky130_fd_sc_hd__inv_2
XFILLER_0_29_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5673_ hold493/X _5629_/X _5653_/X hold363/X _5672_/X vssd1 vssd1 vccd1 vccd1 _5674_/C
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4014__A _6285_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4707__A1 _6380_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4624_ _4602_/Y _4621_/X _4623_/X vssd1 vssd1 vccd1 vccd1 _4624_/X sky130_fd_sc_hd__a21o_1
X_4555_ _6159_/Q _4556_/C vssd1 vssd1 vccd1 vccd1 _4555_/Y sky130_fd_sc_hd__nand2_2
Xhold501 _5392_/X vssd1 vssd1 vccd1 vccd1 _6353_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5380__A1 _5767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4949__A _5064_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold545 _3647_/X vssd1 vssd1 vccd1 vccd1 _6473_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3506_ _5769_/S _3506_/B vssd1 vssd1 vccd1 vccd1 _5400_/B sky130_fd_sc_hd__nand2_1
XANTENNA__3391__B1 _4948_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold534 _5570_/X vssd1 vssd1 vccd1 vccd1 _6373_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold512 _6408_/Q vssd1 vssd1 vccd1 vccd1 hold512/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold523 _6090_/X vssd1 vssd1 vccd1 vccd1 _6486_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout100_A _5567_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4668__B _4668_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold567 _5990_/X vssd1 vssd1 vccd1 vccd1 _6431_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4486_ _3998_/X hold141/X _4491_/S vssd1 vssd1 vccd1 vccd1 _4486_/X sky130_fd_sc_hd__mux2_1
Xhold556 _6372_/Q vssd1 vssd1 vccd1 vccd1 hold556/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5668__C1 _5731_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold578 _6482_/Q vssd1 vssd1 vccd1 vccd1 hold578/X sky130_fd_sc_hd__buf_1
X_3437_ _4335_/B _3668_/B _4588_/A vssd1 vssd1 vccd1 vccd1 _3437_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_0_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold589 _5900_/X vssd1 vssd1 vccd1 vccd1 _6421_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6225_ _6393_/CLK _6225_/D vssd1 vssd1 vccd1 vccd1 _6225_/Q sky130_fd_sc_hd__dfxtp_1
X_3368_ _4720_/C _5757_/C _3368_/S vssd1 vssd1 vccd1 vccd1 _3512_/B sky130_fd_sc_hd__mux2_1
XANTENNA__3694__A1 _5607_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6156_ _6265_/CLK _6156_/D vssd1 vssd1 vccd1 vccd1 _6156_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5107_ _6376_/Q _5107_/B vssd1 vssd1 vccd1 vccd1 _5107_/X sky130_fd_sc_hd__xor2_1
XANTENNA__3999__S _4241_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3299_ _3183_/A _5387_/B _4248_/C _4248_/B vssd1 vssd1 vccd1 vccd1 _3300_/D sky130_fd_sc_hd__a2bb2o_1
X_6087_ _6101_/B _5021_/B _5554_/Y _6036_/X vssd1 vssd1 vccd1 vccd1 _6087_/X sky130_fd_sc_hd__o22a_1
X_5038_ _6155_/Q _6146_/Q _6138_/Q _6182_/Q _5404_/A0 _5078_/S1 vssd1 vssd1 vccd1
+ vccd1 _5038_/X sky130_fd_sc_hd__mux4_1
XANTENNA__3997__A2 _4462_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4946__A1 _6368_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3747__B _4150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput43 _6306_/Q vssd1 vssd1 vccd1 vccd1 io_out[24] sky130_fd_sc_hd__buf_12
Xoutput21 _6525_/X vssd1 vssd1 vccd1 vccd1 io_oeb[24] sky130_fd_sc_hd__buf_12
Xoutput32 _6325_/Q vssd1 vssd1 vccd1 vccd1 io_out[14] sky130_fd_sc_hd__buf_12
XFILLER_0_101_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput54 _6283_/Q vssd1 vssd1 vccd1 vccd1 io_out[5] sky130_fd_sc_hd__buf_12
XANTENNA__4882__B1 _5771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4533__S _4536_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4340_ _4249_/B _5362_/D _4337_/X _4339_/X _5522_/A vssd1 vssd1 vccd1 vccd1 _4340_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_1_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4271_ _4335_/B _3443_/B _4588_/A vssd1 vssd1 vccd1 vccd1 _4271_/X sky130_fd_sc_hd__o21a_1
X_3222_ _3168_/B _3204_/X _3193_/X vssd1 vssd1 vccd1 vccd1 _3222_/X sky130_fd_sc_hd__o21a_1
X_6010_ _4456_/X hold169/X _6011_/S vssd1 vssd1 vccd1 vccd1 _6010_/X sky130_fd_sc_hd__mux2_1
X_3153_ _3326_/B _3360_/B vssd1 vssd1 vccd1 vccd1 _4359_/C sky130_fd_sc_hd__nor2_2
XANTENNA__4873__A0 _6364_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4708__S _4712_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3084_ _6354_/Q vssd1 vssd1 vccd1 vccd1 _5284_/S sky130_fd_sc_hd__inv_2
XFILLER_0_27_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout148_A _4268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3986_ _3986_/A _4273_/B vssd1 vssd1 vccd1 vccd1 _3987_/B sky130_fd_sc_hd__nor2_1
XANTENNA__4670__C _4670_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4928__A1 _6464_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4928__B2 _5109_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5725_ _6315_/Q _5630_/X _5653_/X _6489_/Q _5724_/X vssd1 vssd1 vccd1 vccd1 _5726_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_94_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5656_ _6219_/Q _4406_/B _4235_/S _6112_/Q _5730_/C1 vssd1 vssd1 vccd1 vccd1 _5656_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_32_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5353__A1 _5600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4607_ _4611_/B _4607_/B vssd1 vssd1 vccd1 vccd1 _4607_/X sky130_fd_sc_hd__and2_2
XANTENNA__5353__B2 hold604/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold320 _6305_/Q vssd1 vssd1 vccd1 vccd1 hold320/X sky130_fd_sc_hd__dlygate4sd3_1
X_5587_ _5587_/A _5587_/B vssd1 vssd1 vccd1 vccd1 _5587_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_13_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold331 _4715_/X vssd1 vssd1 vccd1 vccd1 _6308_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold353 hold660/X vssd1 vssd1 vccd1 vccd1 _3594_/A sky130_fd_sc_hd__clkbuf_2
X_4538_ hold87/X _4404_/X _4545_/S vssd1 vssd1 vccd1 vccd1 hold88/A sky130_fd_sc_hd__mux2_1
Xhold342 _6387_/Q vssd1 vssd1 vccd1 vccd1 _3097_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold386 _3637_/X vssd1 vssd1 vccd1 vccd1 _6457_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4469_ hold236/X _4042_/X _4473_/S vssd1 vssd1 vccd1 vccd1 _6181_/D sky130_fd_sc_hd__mux2_1
Xhold364 _6086_/X vssd1 vssd1 vccd1 vccd1 _6485_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold375 _6416_/Q vssd1 vssd1 vccd1 vccd1 hold375/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold397 _6415_/Q vssd1 vssd1 vccd1 vccd1 hold397/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5656__A2 _4406_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6208_ _6455_/CLK _6208_/D vssd1 vssd1 vccd1 vccd1 _6208_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6139_ _6223_/CLK _6139_/D vssd1 vssd1 vccd1 vccd1 _6139_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5957__B _5970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5019__S1 _5100_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4778__S0 _5078_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5867__B _5867_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3668__A _3668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3291__C1 _3352_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3840_ _6206_/Q _3793_/X _3795_/X _6214_/Q vssd1 vssd1 vccd1 vccd1 _3846_/A sky130_fd_sc_hd__a22o_1
X_3771_ _6378_/Q _6382_/Q _6343_/Q vssd1 vssd1 vccd1 vccd1 _5267_/A sky130_fd_sc_hd__mux2_1
X_5510_ hold592/X _4668_/A _5510_/S vssd1 vssd1 vccd1 vccd1 _5510_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_6_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6490_ _6490_/CLK _6490_/D fanout176/X vssd1 vssd1 vccd1 vccd1 _6490_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA__5335__A1 _5757_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5441_ _5492_/A _5441_/B _5441_/C vssd1 vssd1 vccd1 vccd1 _5443_/A sky130_fd_sc_hd__and3_1
X_5372_ _5372_/A _5372_/B _5523_/C _5372_/D vssd1 vssd1 vccd1 vccd1 _5373_/B sky130_fd_sc_hd__or4_1
XFILLER_0_10_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4323_ _5581_/S _4320_/A _5766_/S _6315_/Q _4321_/X vssd1 vssd1 vccd1 vccd1 _4323_/X
+ sky130_fd_sc_hd__o221a_1
Xfanout118 _5866_/A vssd1 vssd1 vccd1 vccd1 _5322_/A sky130_fd_sc_hd__clkbuf_8
Xfanout107 _3276_/Y vssd1 vssd1 vccd1 vccd1 _4289_/C sky130_fd_sc_hd__clkbuf_4
Xfanout129 _4324_/A vssd1 vssd1 vccd1 vccd1 _5995_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4254_ _4313_/A _5387_/C _4267_/B _3379_/A _4261_/A vssd1 vssd1 vccd1 vccd1 _4255_/A
+ sky130_fd_sc_hd__o32a_1
XANTENNA__4846__A0 _4844_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3205_ _3229_/A _3205_/B _3216_/B vssd1 vssd1 vccd1 vccd1 _3205_/X sky130_fd_sc_hd__and3_1
X_4185_ _6158_/Q _3799_/X _3801_/X _6149_/Q vssd1 vssd1 vccd1 vccd1 _4185_/X sky130_fd_sc_hd__a22o_1
X_3136_ _3323_/A _3229_/A _3205_/B _3168_/B vssd1 vssd1 vccd1 vccd1 _3414_/B sky130_fd_sc_hd__or4bb_4
X_3067_ _6467_/Q vssd1 vssd1 vccd1 vccd1 _5146_/A sky130_fd_sc_hd__inv_2
XANTENNA__4962__A _5102_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5777__B _5777_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4681__B _4714_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3297__B _3297_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3969_ _4150_/A _3969_/B vssd1 vssd1 vccd1 vccd1 _3972_/C sky130_fd_sc_hd__nor2_1
X_5708_ _6139_/Q _5721_/A2 _5721_/B1 _6183_/Q _5721_/C1 vssd1 vssd1 vccd1 vccd1 _5709_/B
+ sky130_fd_sc_hd__o221a_1
X_5639_ _5655_/B _5639_/B _5639_/C vssd1 vssd1 vccd1 vccd1 _5639_/X sky130_fd_sc_hd__and3_1
Xhold150 _4520_/X vssd1 vssd1 vccd1 vccd1 _6226_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold161 _6152_/Q vssd1 vssd1 vccd1 vccd1 hold161/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold194 _6221_/Q vssd1 vssd1 vccd1 vccd1 hold194/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold183 _6141_/Q vssd1 vssd1 vccd1 vccd1 hold183/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 _4494_/X vssd1 vssd1 vccd1 vccd1 _6203_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3760__B _4557_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5907__S _5974_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4999__S0 _5404_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3935__B _6337_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3591__A3 _3673_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5208__A _6463_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4782__A _4782_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5990_ _3489_/B _3636_/B _3635_/Y _5989_/X vssd1 vssd1 vccd1 vccd1 _5990_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_91_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4941_ _4949_/B vssd1 vssd1 vccd1 vccd1 _4942_/B sky130_fd_sc_hd__inv_2
XANTENNA__5005__A0 _6423_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4872_ _6416_/Q _4930_/B _4870_/X _4871_/X vssd1 vssd1 vccd1 vccd1 _4872_/X sky130_fd_sc_hd__o22a_1
XANTENNA__5100__S0 _5100_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3823_ _4052_/A _4641_/A vssd1 vssd1 vccd1 vccd1 _4460_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3754_ _5136_/B _3743_/X _3750_/A _3753_/X vssd1 vssd1 vccd1 vccd1 _3754_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_9_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6467_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_42_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5308__A1 _5369_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3685_ _3685_/A _4386_/B vssd1 vssd1 vccd1 vccd1 _4262_/B sky130_fd_sc_hd__or2_2
X_6473_ _6474_/CLK _6473_/D fanout179/X vssd1 vssd1 vccd1 vccd1 _6473_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__4022__A _6381_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5424_ _4957_/S _5512_/S _5520_/B _4300_/A vssd1 vssd1 vccd1 vccd1 _5424_/X sky130_fd_sc_hd__a31o_1
XANTENNA__5859__A2 _5785_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5355_ _5393_/A1 hold612/X _5320_/X _5368_/S vssd1 vssd1 vccd1 vccd1 _6345_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_57_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5286_ _3774_/A _5284_/X _5285_/X _4115_/A vssd1 vssd1 vccd1 vccd1 _5286_/X sky130_fd_sc_hd__a22o_1
X_4306_ _4310_/S _4309_/B _4300_/A vssd1 vssd1 vccd1 vccd1 _4306_/X sky130_fd_sc_hd__a21o_1
XANTENNA__3580__B _3619_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4237_ hold242/X _4406_/B _4235_/S hold234/X _5730_/C1 vssd1 vssd1 vccd1 vccd1 _4237_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_97_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4168_ _4332_/B _4168_/B vssd1 vssd1 vccd1 vccd1 _4168_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_65_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3119_ _3323_/A _3168_/B _3326_/A vssd1 vssd1 vccd1 vccd1 _3167_/B sky130_fd_sc_hd__and3_1
X_4099_ _4199_/A _6289_/Q _6383_/Q _4060_/B _4098_/X vssd1 vssd1 vccd1 vccd1 _5257_/B
+ sky130_fd_sc_hd__o41a_2
XANTENNA__5244__A0 _6314_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4598__A2 _4324_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4631__S _4641_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4867__A _4924_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4589__A2 _5777_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5210__B _6458_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4541__S _4545_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3470_ _3636_/B vssd1 vssd1 vccd1 vccd1 _3471_/B sky130_fd_sc_hd__inv_2
X_5140_ _5605_/A _5268_/A _4217_/X vssd1 vssd1 vccd1 vccd1 _5140_/X sky130_fd_sc_hd__a21o_1
XANTENNA__3721__B1 _4441_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5071_ _6426_/Q _4793_/Y _5065_/X _5070_/X vssd1 vssd1 vccd1 vccd1 _5071_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_19_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4022_ _6381_/Q _4022_/B vssd1 vssd1 vccd1 vccd1 _4022_/X sky130_fd_sc_hd__or2_1
XANTENNA__5226__A0 _6381_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4943__C _6367_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5973_ _5964_/A _5972_/X _5102_/Y vssd1 vssd1 vccd1 vccd1 _5973_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_87_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4924_ _4922_/X _4924_/B _4924_/C vssd1 vssd1 vccd1 vccd1 _4929_/A sky130_fd_sc_hd__and3b_1
XANTENNA__4044__A4 _4036_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4855_ _4854_/X _6363_/Q _5861_/S vssd1 vssd1 vccd1 vccd1 _4856_/B sky130_fd_sc_hd__mux2_1
XANTENNA__5547__S _6070_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5529__A1 _4982_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4786_ _5322_/A _4786_/B _4786_/C _5523_/B vssd1 vssd1 vccd1 vccd1 _4787_/B sky130_fd_sc_hd__or4_2
XFILLER_0_7_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3806_ _3816_/B _3885_/A vssd1 vssd1 vccd1 vccd1 _3811_/B sky130_fd_sc_hd__nor2_1
X_3737_ _4087_/B vssd1 vssd1 vccd1 vccd1 _4227_/S sky130_fd_sc_hd__inv_4
X_6525_ _6529_/A vssd1 vssd1 vccd1 vccd1 _6525_/X sky130_fd_sc_hd__buf_1
XFILLER_0_70_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3960__B1 _3810_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3668_ _3668_/A _3668_/B vssd1 vssd1 vccd1 vccd1 _3668_/Y sky130_fd_sc_hd__nor2_1
X_6456_ _6456_/CLK _6456_/D vssd1 vssd1 vccd1 vccd1 _6456_/Q sky130_fd_sc_hd__dfxtp_1
X_5407_ _5774_/B _5407_/B _5774_/C _3379_/B vssd1 vssd1 vccd1 vccd1 _5407_/X sky130_fd_sc_hd__or4b_1
X_3599_ _3699_/A _3597_/Y _3598_/Y _3602_/B vssd1 vssd1 vccd1 vccd1 _3603_/A sky130_fd_sc_hd__a211o_1
XANTENNA__5701__A1 _4300_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6387_ _6412_/CLK _6387_/D vssd1 vssd1 vccd1 vccd1 _6387_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5338_ _4675_/A _3590_/A _5387_/C _5323_/C vssd1 vssd1 vccd1 vccd1 _5338_/X sky130_fd_sc_hd__a31o_1
X_5269_ _3770_/Y _5267_/X _5268_/X _5200_/X _5202_/Y vssd1 vssd1 vccd1 vccd1 _5269_/X
+ sky130_fd_sc_hd__o311a_1
XANTENNA_clkbuf_leaf_18_wb_clk_i_A _6448_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4626__S _4641_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold607_A _6364_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4536__S _4536_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6340__SET_B fanout183/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4640_ _5393_/A1 hold548/X _4582_/Y _4639_/X vssd1 vssd1 vccd1 vccd1 _4640_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4571_ hold510/X _6336_/Q _4575_/S vssd1 vssd1 vccd1 vccd1 _4571_/X sky130_fd_sc_hd__mux2_1
X_6310_ _6316_/CLK _6310_/D fanout174/X vssd1 vssd1 vccd1 vccd1 _6310_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_0_12_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3522_ _6447_/Q _5309_/A _6442_/Q vssd1 vssd1 vccd1 vccd1 _3522_/X sky130_fd_sc_hd__and3b_2
XFILLER_0_97_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3453_ _3617_/A _3406_/Y _5619_/A _3674_/A vssd1 vssd1 vccd1 vccd1 _3453_/X sky130_fd_sc_hd__o22a_1
X_6241_ _6456_/CLK hold62/X vssd1 vssd1 vccd1 vccd1 hold61/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__4300__A _4300_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6172_ _6449_/CLK _6172_/D vssd1 vssd1 vccd1 vccd1 _6172_/Q sky130_fd_sc_hd__dfxtp_1
X_3384_ _3285_/Y _3353_/X _3355_/X _3383_/X _3342_/X vssd1 vssd1 vccd1 vccd1 _3384_/X
+ sky130_fd_sc_hd__a32o_1
X_5123_ _5123_/A vssd1 vssd1 vccd1 vccd1 _5123_/Y sky130_fd_sc_hd__inv_2
XANTENNA__5998__A1 _5995_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5054_ _5964_/A _5053_/X _5041_/Y vssd1 vssd1 vccd1 vccd1 _5054_/X sky130_fd_sc_hd__a21bo_1
X_4005_ _4005_/A _4005_/B vssd1 vssd1 vccd1 vccd1 _4007_/A sky130_fd_sc_hd__nor2_1
XANTENNA_fanout178_A fanout180/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5956_ _5951_/A _5785_/Y _5955_/X _5977_/S vssd1 vssd1 vccd1 vccd1 _5956_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_62_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5887_ _5879_/X _5886_/Y _5887_/S vssd1 vssd1 vccd1 vccd1 _5887_/X sky130_fd_sc_hd__mux2_1
X_4907_ _6366_/Q _4922_/C _4924_/C vssd1 vssd1 vccd1 vccd1 _4907_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_90_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4838_ _6121_/Q _5783_/A vssd1 vssd1 vccd1 vccd1 _4838_/X sky130_fd_sc_hd__and2_1
XFILLER_0_7_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4186__B1 _3795_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4769_ _4767_/X _4768_/X _5289_/S vssd1 vssd1 vccd1 vccd1 _4769_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_15_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3933__B1 _6287_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6439_ _6439_/CLK _6439_/D fanout178/X vssd1 vssd1 vccd1 vccd1 _6439_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold21 hold21/A vssd1 vssd1 vccd1 vccd1 hold21/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold10 hold10/A vssd1 vssd1 vccd1 vccd1 hold10/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 hold32/A vssd1 vssd1 vccd1 vccd1 hold32/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 hold43/A vssd1 vssd1 vccd1 vccd1 hold43/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 hold65/A vssd1 vssd1 vccd1 vccd1 hold65/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 hold54/A vssd1 vssd1 vccd1 vccd1 hold54/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4356__S _5769_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold87 hold87/A vssd1 vssd1 vccd1 vccd1 hold87/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 hold76/A vssd1 vssd1 vccd1 vccd1 hold76/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold98 hold98/A vssd1 vssd1 vccd1 vccd1 hold98/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5041__A _5102_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6476__SET_B fanout176/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_7 _6336_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_23_wb_clk_i _6448_/CLK vssd1 vssd1 vccd1 vccd1 _6383_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__6047__A _6081_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xci2406_z80_211 vssd1 vssd1 vccd1 vccd1 ci2406_z80_211/HI io_out[30] sky130_fd_sc_hd__conb_1
XFILLER_0_88_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xci2406_z80_200 vssd1 vssd1 vccd1 vccd1 ci2406_z80_200/HI io_oeb[15] sky130_fd_sc_hd__conb_1
XANTENNA__4790__A _6431_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5810_ _5867_/B _5809_/C _6415_/Q vssd1 vssd1 vccd1 vccd1 _5811_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_29_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4404__A1 _4418_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5741_ _3097_/Y _4611_/A _5769_/S vssd1 vssd1 vccd1 vccd1 _5742_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_44_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5097__S _6070_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5672_ _6311_/Q _5630_/X _5632_/Y _5671_/X vssd1 vssd1 vccd1 vccd1 _5672_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4014__B _6286_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5904__A1 _6422_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4623_ _6478_/Q _4604_/X _4605_/X _6486_/Q _4622_/X vssd1 vssd1 vccd1 vccd1 _4623_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3915__B1 _6285_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold502 _6407_/Q vssd1 vssd1 vccd1 vccd1 hold502/X sky130_fd_sc_hd__buf_1
X_4554_ _4240_/X hold153/X _4554_/S vssd1 vssd1 vccd1 vccd1 _4554_/X sky130_fd_sc_hd__mux2_1
X_3505_ _3665_/A _5769_/S _5418_/A vssd1 vssd1 vccd1 vccd1 _3527_/C sky130_fd_sc_hd__and3_1
XANTENNA__3391__A1 _5109_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold513 _5764_/X vssd1 vssd1 vccd1 vccd1 _6408_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold535 _6487_/Q vssd1 vssd1 vccd1 vccd1 hold535/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4949__B _4949_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold524 _6419_/Q vssd1 vssd1 vccd1 vccd1 hold524/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold579 _6424_/Q vssd1 vssd1 vccd1 vccd1 _5922_/A sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold546 _6427_/Q vssd1 vssd1 vccd1 vccd1 hold546/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold557 _5558_/X vssd1 vssd1 vccd1 vccd1 _6372_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6224_ _6265_/CLK _6224_/D vssd1 vssd1 vccd1 vccd1 _6224_/Q sky130_fd_sc_hd__dfxtp_1
X_4485_ _3954_/X hold226/X _4491_/S vssd1 vssd1 vccd1 vccd1 _4485_/X sky130_fd_sc_hd__mux2_1
Xhold568 _6422_/Q vssd1 vssd1 vccd1 vccd1 _5901_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3436_ _3477_/A _6433_/Q _3489_/B vssd1 vssd1 vccd1 vccd1 _3668_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3367_ _4217_/A _3511_/A _6339_/Q vssd1 vssd1 vccd1 vccd1 _3367_/X sky130_fd_sc_hd__o21ba_1
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6155_ _6263_/CLK _6155_/D vssd1 vssd1 vccd1 vccd1 _6155_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5106_ _5102_/B _5105_/X _5106_/S vssd1 vssd1 vccd1 vccd1 _5106_/X sky130_fd_sc_hd__mux2_1
X_6086_ _4366_/A _6084_/X _6085_/Y hold363/X _6077_/Y vssd1 vssd1 vccd1 vccd1 _6086_/X
+ sky130_fd_sc_hd__o32a_1
X_3298_ _4313_/A _5360_/A _3296_/Y _3297_/Y _5866_/A vssd1 vssd1 vccd1 vccd1 _3298_/X
+ sky130_fd_sc_hd__a41o_1
X_5037_ _5036_/X hold369/X _5098_/S vssd1 vssd1 vccd1 vccd1 _5037_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_79_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4643__A1 hold628/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4643__B2 hold629/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3851__C1 _3885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4904__S _4948_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5939_ _6373_/Q _5848_/S _5972_/B1 _5938_/X vssd1 vssd1 vccd1 vccd1 _5939_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_35_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput33 _6326_/Q vssd1 vssd1 vccd1 vccd1 io_out[15] sky130_fd_sc_hd__buf_12
Xoutput22 _6526_/X vssd1 vssd1 vccd1 vccd1 io_oeb[25] sky130_fd_sc_hd__buf_12
XFILLER_0_101_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput44 _6307_/Q vssd1 vssd1 vccd1 vccd1 io_out[25] sky130_fd_sc_hd__buf_12
XFILLER_0_9_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput55 _6321_/Q vssd1 vssd1 vccd1 vccd1 io_out[6] sky130_fd_sc_hd__buf_12
XFILLER_0_37_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3358__A_N _5605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4882__A1 _4361_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4594__B _4595_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4086__S _4241_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6084__B1 _6107_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3673__B _3673_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4270_ _4253_/Y _4269_/X _5605_/C vssd1 vssd1 vccd1 vccd1 _4270_/X sky130_fd_sc_hd__o21a_1
X_3221_ _3221_/A _3221_/B _3221_/C _3221_/D vssd1 vssd1 vccd1 vccd1 _3235_/A sky130_fd_sc_hd__and4_1
X_3152_ _5605_/B _5605_/C vssd1 vssd1 vccd1 vccd1 _3360_/B sky130_fd_sc_hd__nand2b_2
XANTENNA__6369__RESET_B fanout172/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6075__B1 _6107_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3083_ _3083_/A vssd1 vssd1 vccd1 vccd1 _3083_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4625__A1 _5757_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4625__B2 _4624_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3985_ _3770_/A _5267_/C _5262_/A _4115_/A _3979_/A vssd1 vssd1 vccd1 vccd1 _3985_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_9_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5050__B2 _4924_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5050__A1 _5109_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4928__A2 _4963_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5724_ _6464_/Q _5645_/X _5723_/X _5632_/Y vssd1 vssd1 vccd1 vccd1 _5724_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_45_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5655_ _5655_/A _5655_/B vssd1 vssd1 vccd1 vccd1 _5655_/X sky130_fd_sc_hd__or2_1
XFILLER_0_17_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3864__A _3883_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4606_ _4641_/B _4607_/B vssd1 vssd1 vccd1 vccd1 _4606_/X sky130_fd_sc_hd__and2_2
Xhold310 _6301_/Q vssd1 vssd1 vccd1 vccd1 hold310/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5586_ _5576_/A _5576_/B _5574_/A vssd1 vssd1 vccd1 vccd1 _5587_/B sky130_fd_sc_hd__o21ai_1
Xhold321 _4700_/X vssd1 vssd1 vccd1 vccd1 _6305_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold332 _6127_/Q vssd1 vssd1 vccd1 vccd1 hold332/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold343 _6386_/Q vssd1 vssd1 vccd1 vccd1 _3096_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4537_ _4537_/A _6003_/B vssd1 vssd1 vccd1 vccd1 _4545_/S sky130_fd_sc_hd__nor2_4
Xhold365 _6257_/Q vssd1 vssd1 vccd1 vccd1 hold365/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold354 _6027_/X vssd1 vssd1 vccd1 vccd1 _6468_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold387 _6327_/Q vssd1 vssd1 vccd1 vccd1 hold387/X sky130_fd_sc_hd__dlygate4sd3_1
X_4468_ hold214/X _3998_/X _4473_/S vssd1 vssd1 vccd1 vccd1 _6180_/D sky130_fd_sc_hd__mux2_1
Xhold376 _5833_/X vssd1 vssd1 vccd1 vccd1 _6416_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3419_ _3590_/A _3419_/B vssd1 vssd1 vccd1 vccd1 _5316_/B sky130_fd_sc_hd__or2_2
Xhold398 _5820_/X vssd1 vssd1 vccd1 vccd1 _6415_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6207_ _6455_/CLK _6207_/D vssd1 vssd1 vccd1 vccd1 hold99/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__3667__A2 _3352_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4399_ _3695_/Y _3717_/A _4398_/X _5384_/A vssd1 vssd1 vccd1 vccd1 _6003_/B sky130_fd_sc_hd__a31o_4
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6138_ _6400_/CLK _6138_/D vssd1 vssd1 vccd1 vccd1 _6138_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4864__A1 _5102_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6069_ _6100_/A _4949_/B _5508_/Y _6037_/B vssd1 vssd1 vccd1 vccd1 _6070_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_95_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3477__C _5387_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5465__S _5593_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4778__S1 _5404_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6462__RESET_B fanout181/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4083__A2 _4462_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4544__S _4545_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3291__B1 _3668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3770_ _3770_/A vssd1 vssd1 vccd1 vccd1 _3770_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_27_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5440_ _6477_/Q _4844_/X _5593_/S vssd1 vssd1 vccd1 vccd1 _5441_/C sky130_fd_sc_hd__mux2_1
XFILLER_0_89_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3346__A1 _4268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5371_ _5371_/A _5371_/B _5371_/C _5371_/D vssd1 vssd1 vccd1 vccd1 _5372_/D sky130_fd_sc_hd__or4_1
XFILLER_0_50_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4322_ _5581_/S _4322_/B vssd1 vssd1 vccd1 vccd1 _5766_/S sky130_fd_sc_hd__nand2_1
Xfanout108 _3514_/B vssd1 vssd1 vccd1 vccd1 _4325_/C sky130_fd_sc_hd__buf_4
X_4253_ _4253_/A _5336_/A vssd1 vssd1 vccd1 vccd1 _4253_/Y sky130_fd_sc_hd__nor2_1
Xfanout119 _3062_/Y vssd1 vssd1 vccd1 vccd1 _5866_/A sky130_fd_sc_hd__clkbuf_8
X_3204_ _3323_/A _3326_/A _3205_/B vssd1 vssd1 vccd1 vccd1 _3204_/X sky130_fd_sc_hd__or3_2
XFILLER_0_10_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4184_ _4149_/A _4149_/B _4147_/A vssd1 vssd1 vccd1 vccd1 _4191_/A sky130_fd_sc_hd__a21o_1
X_3135_ _3323_/A _3211_/B _4782_/B vssd1 vssd1 vccd1 vccd1 _5387_/B sky130_fd_sc_hd__or3_4
XFILLER_0_96_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3066_ _5593_/S vssd1 vssd1 vccd1 vccd1 _5757_/A sky130_fd_sc_hd__inv_4
XFILLER_0_54_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4962__B _4962_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout160_A _3172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3821__A2 _3731_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3968_ _5136_/A _6380_/Q vssd1 vssd1 vccd1 vccd1 _3972_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_18_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5707_ _6223_/Q _5721_/A2 _5721_/B1 _6116_/Q _5730_/C1 vssd1 vssd1 vccd1 vccd1 _5709_/A
+ sky130_fd_sc_hd__o221a_1
XANTENNA__5285__S _5866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3899_ _3839_/B _3847_/B _4190_/A vssd1 vssd1 vccd1 vccd1 _4451_/C sky130_fd_sc_hd__o21a_1
XFILLER_0_72_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5638_ _5655_/B _5633_/X _5634_/X _5637_/X vssd1 vssd1 vccd1 vccd1 _5638_/X sky130_fd_sc_hd__a31o_1
X_5569_ _6462_/Q _5598_/S _5568_/X vssd1 vssd1 vccd1 vccd1 _5569_/X sky130_fd_sc_hd__o21ba_1
XANTENNA__5731__C1 _5731_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold151 _6237_/Q vssd1 vssd1 vccd1 vccd1 hold151/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold162 _4391_/X vssd1 vssd1 vccd1 vccd1 _6152_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold140 _4397_/X vssd1 vssd1 vccd1 vccd1 _6158_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 _6145_/Q vssd1 vssd1 vccd1 vccd1 hold173/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 _6135_/Q vssd1 vssd1 vccd1 vccd1 hold195/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold184 _4376_/X vssd1 vssd1 vccd1 vccd1 _6141_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout73_A _3909_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5798__C1 _5771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold637_A _6315_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4999__S1 _5100_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5208__B _6462_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold1_A hold1/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4539__S _4545_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output54_A _6283_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4940_ _5101_/S _4939_/X _4938_/Y vssd1 vssd1 vccd1 vccd1 _4949_/B sky130_fd_sc_hd__o21ai_4
XANTENNA__6055__A _6089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4871_ _6461_/Q _4963_/B _4869_/X _3387_/Y _4867_/X vssd1 vssd1 vccd1 vccd1 _4871_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_74_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3822_ _3822_/A _3822_/B _3822_/C vssd1 vssd1 vccd1 vccd1 _4641_/A sky130_fd_sc_hd__or3_2
XFILLER_0_61_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5100__S1 _5100_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3753_ _6345_/Q _6343_/Q _5136_/A vssd1 vssd1 vccd1 vccd1 _3753_/X sky130_fd_sc_hd__and3_2
XFILLER_0_54_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5308__A2 _5757_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3684_ _3693_/A vssd1 vssd1 vccd1 vccd1 _3684_/Y sky130_fd_sc_hd__inv_2
X_6472_ _6472_/CLK hold78/X fanout177/X vssd1 vssd1 vccd1 vccd1 hold45/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5423_ _5485_/S _5484_/S vssd1 vssd1 vccd1 vccd1 _5520_/B sky130_fd_sc_hd__and2_4
X_5354_ _5757_/B _4150_/A _5368_/S hold605/X vssd1 vssd1 vccd1 vccd1 _5354_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_2_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4305_ _4312_/A _5783_/A _5418_/A _4312_/D vssd1 vssd1 vccd1 vccd1 _4309_/B sky130_fd_sc_hd__nand4_1
X_5285_ _6340_/Q _5263_/B _5866_/A vssd1 vssd1 vccd1 vccd1 _5285_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_10_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4449__S _4464_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4236_ hold183/X _4406_/B _4235_/S hold145/X _5731_/C1 vssd1 vssd1 vccd1 vccd1 _4236_/X
+ sky130_fd_sc_hd__o221a_1
X_4167_ _4163_/Y _4166_/Y _6334_/Q vssd1 vssd1 vccd1 vccd1 _5171_/A sky130_fd_sc_hd__mux2_2
X_3118_ _4268_/A _4273_/A _6300_/Q _6299_/Q vssd1 vssd1 vccd1 vccd1 _3614_/A sky130_fd_sc_hd__or4bb_4
XFILLER_0_65_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4098_ _4060_/B _4094_/Y _4095_/X _4097_/X vssd1 vssd1 vccd1 vccd1 _4098_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_97_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4047__A2 _3793_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5704__C1 _5730_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5743__S _5769_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_47_wb_clk_i_A clkbuf_leaf_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__4883__A _6364_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3499__A _5384_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_48_wb_clk_i clkbuf_leaf_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6265_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_83_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout90 _4361_/B vssd1 vssd1 vccd1 vccd1 _5102_/A sky130_fd_sc_hd__buf_4
XFILLER_0_101_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5070_ _5109_/A1 _5067_/X _5069_/X _4924_/C vssd1 vssd1 vccd1 vccd1 _5070_/X sky130_fd_sc_hd__a22o_1
X_4021_ _3762_/Y _4223_/A _4022_/B vssd1 vssd1 vccd1 vccd1 _4021_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4793__A _4930_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5889__A _6421_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5972_ _6376_/Q _5848_/S _5972_/B1 _5971_/X vssd1 vssd1 vccd1 vccd1 _5972_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4943__D _6368_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4985__A0 _6422_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4923_ _6366_/Q _4922_/C _6367_/Q vssd1 vssd1 vccd1 vccd1 _4924_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_47_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4732__S _4768_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4854_ _5892_/S _4852_/X _4853_/X _4841_/X vssd1 vssd1 vccd1 vccd1 _4854_/X sky130_fd_sc_hd__a31o_1
X_4785_ _4785_/A _4785_/B _4785_/C vssd1 vssd1 vccd1 vccd1 _5523_/B sky130_fd_sc_hd__or3_1
XFILLER_0_43_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3805_ _3852_/A _3885_/A _3865_/S vssd1 vssd1 vccd1 vccd1 _6003_/A sky130_fd_sc_hd__or3_1
X_3736_ _5600_/A _5360_/A _5314_/S _4338_/B vssd1 vssd1 vccd1 vccd1 _4087_/B sky130_fd_sc_hd__and4_2
XANTENNA__5129__A _6021_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout123_A _5384_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6524_ _6529_/A vssd1 vssd1 vccd1 vccd1 _6524_/X sky130_fd_sc_hd__buf_1
X_3667_ _3786_/A _3352_/B _5387_/C _5146_/D _5146_/B vssd1 vssd1 vccd1 vccd1 _3667_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_0_2_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6455_ _6455_/CLK _6455_/D vssd1 vssd1 vccd1 vccd1 _6455_/Q sky130_fd_sc_hd__dfxtp_1
X_5406_ _5777_/A _5406_/B vssd1 vssd1 vccd1 vccd1 _5407_/B sky130_fd_sc_hd__nor2_1
X_3598_ _4324_/B _3593_/X _6529_/A vssd1 vssd1 vccd1 vccd1 _3598_/Y sky130_fd_sc_hd__o21ai_1
X_6386_ _6412_/CLK _6386_/D vssd1 vssd1 vccd1 vccd1 _6386_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5337_ _3172_/A _4784_/D _5336_/X _3511_/A _3632_/D vssd1 vssd1 vccd1 vccd1 _5337_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_11_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5268_ _5268_/A _6288_/Q _6289_/Q _6290_/Q vssd1 vssd1 vccd1 vccd1 _5268_/X sky130_fd_sc_hd__or4_1
X_4219_ _6333_/Q _4022_/B _4116_/A _5268_/A _4218_/X vssd1 vssd1 vccd1 vccd1 _5263_/B
+ sky130_fd_sc_hd__a221o_2
XANTENNA__4899__S0 _5100_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5465__A1 _4881_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5799__A _5866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5199_ _5199_/A _5199_/B _5199_/C _4223_/A vssd1 vssd1 vccd1 vccd1 _5199_/X sky130_fd_sc_hd__or4b_1
XANTENNA__4976__A0 _6458_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold502_A _6407_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3400__B1 _4325_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_3_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__3782__A _6076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5000__S0 _5404_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4742__A1_N _6312_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4552__S _4554_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4570_ hold448/X _6335_/Q _4575_/S vssd1 vssd1 vccd1 vccd1 _4570_/X sky130_fd_sc_hd__mux2_1
X_3521_ _5617_/B _5522_/D _5617_/A vssd1 vssd1 vccd1 vccd1 _3521_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_40_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3452_ _3399_/X _3411_/Y _5777_/A vssd1 vssd1 vccd1 vccd1 _3452_/Y sky130_fd_sc_hd__o21ai_1
X_6240_ _6452_/CLK hold52/X vssd1 vssd1 vccd1 vccd1 hold51/A sky130_fd_sc_hd__dfxtp_1
X_3383_ _3317_/X _3372_/Y _3380_/X _3382_/Y vssd1 vssd1 vccd1 vccd1 _3383_/X sky130_fd_sc_hd__o211a_1
X_6171_ _6237_/CLK hold64/X vssd1 vssd1 vccd1 vccd1 hold63/A sky130_fd_sc_hd__dfxtp_1
X_5122_ _6021_/S wire92/X vssd1 vssd1 vccd1 vccd1 _5123_/A sky130_fd_sc_hd__or2_1
XANTENNA__5447__A1 _4658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4727__S _5289_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5053_ _6373_/Q _5848_/S _5972_/B1 _5052_/X vssd1 vssd1 vccd1 vccd1 _5053_/X sky130_fd_sc_hd__a22o_1
X_4004_ _6287_/Q _4004_/B _4004_/C vssd1 vssd1 vccd1 vccd1 _4005_/B sky130_fd_sc_hd__nor3_1
X_5955_ _5786_/Y _5948_/X _5954_/X _5976_/S vssd1 vssd1 vccd1 vccd1 _5955_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5558__S _6104_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4422__A2 _6355_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5886_ _5886_/A _5890_/B vssd1 vssd1 vccd1 vccd1 _5886_/Y sky130_fd_sc_hd__nor2_1
X_4906_ _6480_/Q _5104_/A2 _4796_/Y _4901_/B _4793_/Y vssd1 vssd1 vccd1 vccd1 _4906_/X
+ sky130_fd_sc_hd__a221o_1
X_4837_ _6362_/Q _5863_/S vssd1 vssd1 vccd1 vccd1 _4837_/X sky130_fd_sc_hd__or2_1
XANTENNA__5058__S0 _5100_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4768_ hold572/X hold274/X _4768_/S vssd1 vssd1 vccd1 vccd1 _4768_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3933__A1 _6285_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5293__S _5489_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4699_ _4713_/A _4698_/X _4714_/S vssd1 vssd1 vccd1 vccd1 _4699_/X sky130_fd_sc_hd__o21a_1
X_3719_ _3714_/X _3717_/Y _3718_/X vssd1 vssd1 vccd1 vccd1 _3852_/A sky130_fd_sc_hd__o21a_4
X_6438_ _6439_/CLK _6438_/D fanout178/X vssd1 vssd1 vccd1 vccd1 _6438_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5686__A1 _6312_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6369_ _6480_/CLK _6369_/D fanout172/X vssd1 vssd1 vccd1 vccd1 _6369_/Q sky130_fd_sc_hd__dfrtp_1
Xhold22 hold22/A vssd1 vssd1 vccd1 vccd1 hold22/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold11 hold11/A vssd1 vssd1 vccd1 vccd1 hold11/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 hold44/A vssd1 vssd1 vccd1 vccd1 hold44/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 hold55/A vssd1 vssd1 vccd1 vccd1 hold55/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 hold33/A vssd1 vssd1 vccd1 vccd1 hold33/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5322__A _5322_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold452_A _6284_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold77 hold77/A vssd1 vssd1 vccd1 vccd1 hold77/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 hold66/A vssd1 vssd1 vccd1 vccd1 hold66/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 hold88/A vssd1 vssd1 vccd1 vccd1 hold88/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 hold99/A vssd1 vssd1 vccd1 vccd1 hold99/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4661__A2 _4652_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5041__B _5041_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4372__S _4376_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_8 _4934_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5677__A1 _6336_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5677__B2 _6424_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5931__S _5977_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4547__S _4554_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xci2406_z80_212 vssd1 vssd1 vccd1 vccd1 ci2406_z80_212/HI io_out[31] sky130_fd_sc_hd__conb_1
Xci2406_z80_201 vssd1 vssd1 vccd1 vccd1 ci2406_z80_201/HI io_oeb[16] sky130_fd_sc_hd__conb_1
XFILLER_0_16_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4790__B _6442_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5740_ _5740_/A vssd1 vssd1 vccd1 vccd1 _6386_/D sky130_fd_sc_hd__inv_2
XANTENNA__6063__A _6097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5671_ _4424_/X _5670_/X _5734_/S vssd1 vssd1 vccd1 vccd1 _5671_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4014__C _6287_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4622_ _6461_/Q _4606_/X _4607_/X _6312_/Q vssd1 vssd1 vccd1 vccd1 _4622_/X sky130_fd_sc_hd__a22o_1
X_4553_ _4182_/X hold128/X _4554_/S vssd1 vssd1 vccd1 vccd1 _4553_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold514 _6275_/Q vssd1 vssd1 vccd1 vccd1 hold514/X sky130_fd_sc_hd__dlygate4sd3_1
X_3504_ _4325_/A _6019_/S vssd1 vssd1 vccd1 vccd1 _3506_/B sky130_fd_sc_hd__nor2_2
Xhold503 _5763_/X vssd1 vssd1 vccd1 vccd1 _6407_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4484_ _3911_/X hold276/X _4491_/S vssd1 vssd1 vccd1 vccd1 _6194_/D sky130_fd_sc_hd__mux2_1
Xhold536 _6094_/X vssd1 vssd1 vccd1 vccd1 _6487_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold525 _5874_/X vssd1 vssd1 vccd1 vccd1 _6419_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3435_ _3632_/D _3434_/B _3409_/Y vssd1 vssd1 vccd1 vccd1 _3440_/B sky130_fd_sc_hd__o21a_1
Xhold558 _6442_/Q vssd1 vssd1 vccd1 vccd1 _4653_/A sky130_fd_sc_hd__clkbuf_2
Xhold547 _5967_/X vssd1 vssd1 vccd1 vccd1 _6427_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6223_ _6223_/CLK _6223_/D vssd1 vssd1 vccd1 vccd1 _6223_/Q sky130_fd_sc_hd__dfxtp_1
Xhold569 _5909_/X vssd1 vssd1 vccd1 vccd1 _6422_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3366_ _4716_/A _5605_/B vssd1 vssd1 vccd1 vccd1 _5757_/C sky130_fd_sc_hd__or2_2
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6154_ _6239_/CLK hold74/X vssd1 vssd1 vccd1 vccd1 hold73/A sky130_fd_sc_hd__dfxtp_1
X_3297_ _3652_/B _3297_/B vssd1 vssd1 vccd1 vccd1 _3297_/Y sky130_fd_sc_hd__nand2_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5105_ _6428_/Q _6376_/Q _5105_/S vssd1 vssd1 vccd1 vccd1 _5105_/X sky130_fd_sc_hd__mux2_1
X_6085_ _6085_/A _6107_/S vssd1 vssd1 vccd1 vccd1 _6085_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__4457__S _4464_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5036_ _6405_/Q _5035_/X _6070_/A vssd1 vssd1 vccd1 vccd1 _5036_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_32_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6482__SET_B fanout176/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5938_ _6406_/Q _6425_/Q _5971_/S vssd1 vssd1 vccd1 vccd1 _5938_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_75_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5869_ _5867_/B _5867_/C _6419_/Q vssd1 vssd1 vccd1 vccd1 _5870_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_35_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5108__A0 _6465_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput34 _6327_/Q vssd1 vssd1 vccd1 vccd1 io_out[16] sky130_fd_sc_hd__buf_12
Xoutput23 _6527_/X vssd1 vssd1 vccd1 vccd1 io_oeb[26] sky130_fd_sc_hd__buf_12
Xoutput45 _6303_/Q vssd1 vssd1 vccd1 vccd1 io_out[26] sky130_fd_sc_hd__buf_12
Xoutput56 _6320_/Q vssd1 vssd1 vccd1 vccd1 io_out[7] sky130_fd_sc_hd__buf_12
XANTENNA__5751__S _6104_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4882__A2 _4881_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5831__A1 _6364_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4570__A1 _6335_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3392__D _5369_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4858__C1 _5783_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3220_ _3240_/B _3204_/X _3219_/Y vssd1 vssd1 vccd1 vccd1 _3221_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_94_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3151_ _5605_/B _5315_/A vssd1 vssd1 vccd1 vccd1 _5398_/A sky130_fd_sc_hd__nor2_4
XFILLER_0_27_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3082_ _6380_/Q vssd1 vssd1 vccd1 vccd1 _3969_/B sky130_fd_sc_hd__inv_2
XANTENNA__4181__S0 _5721_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3984_ _6285_/Q _6287_/Q _4716_/A vssd1 vssd1 vccd1 vccd1 _5262_/A sky130_fd_sc_hd__mux2_1
XANTENNA__3210__A _4675_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5723_ _4455_/X _5719_/X _4181_/X _5722_/X _5655_/B _5734_/S vssd1 vssd1 vccd1 vccd1
+ _5723_/X sky130_fd_sc_hd__mux4_2
XFILLER_0_45_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4740__S _4770_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5654_ _6422_/Q _5643_/X _5645_/X _6459_/Q vssd1 vssd1 vccd1 vccd1 _5654_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_72_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4605_ _5767_/A _4605_/B _4605_/C _4611_/B vssd1 vssd1 vccd1 vccd1 _4605_/X sky130_fd_sc_hd__and4_2
Xhold311 _4680_/X vssd1 vssd1 vccd1 vccd1 _6301_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4561__A1 _6310_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5585_ _5585_/A _5585_/B vssd1 vssd1 vccd1 vccd1 _5587_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold300 _6456_/Q vssd1 vssd1 vccd1 vccd1 hold300/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold333 _4356_/X vssd1 vssd1 vccd1 vccd1 _6127_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4536_ hold61/X _4463_/X _4536_/S vssd1 vssd1 vccd1 vccd1 hold62/A sky130_fd_sc_hd__mux2_1
Xhold344 _6125_/Q vssd1 vssd1 vccd1 vccd1 _4319_/B sky130_fd_sc_hd__clkbuf_2
Xhold322 _6356_/Q vssd1 vssd1 vccd1 vccd1 hold322/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold366 _3552_/X vssd1 vssd1 vccd1 vccd1 _6257_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold377 _6128_/Q vssd1 vssd1 vccd1 vccd1 _4919_/S sky130_fd_sc_hd__buf_2
X_4467_ hold136/X _3954_/X _4473_/S vssd1 vssd1 vccd1 vccd1 _4467_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5571__S _5593_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold355 _6320_/Q vssd1 vssd1 vccd1 vccd1 hold355/X sky130_fd_sc_hd__dlygate4sd3_1
X_3418_ _3284_/B _3268_/B _3587_/B vssd1 vssd1 vccd1 vccd1 _3419_/B sky130_fd_sc_hd__o21ai_1
Xhold399 _6384_/Q vssd1 vssd1 vccd1 vccd1 _3083_/A sky130_fd_sc_hd__buf_1
X_4398_ _5117_/A _4398_/B _4670_/C vssd1 vssd1 vccd1 vccd1 _4398_/X sky130_fd_sc_hd__or3b_2
Xhold388 _5017_/X vssd1 vssd1 vccd1 vccd1 _6327_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6206_ _6454_/CLK _6206_/D vssd1 vssd1 vccd1 vccd1 _6206_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3667__A3 _5387_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3349_ _3258_/B _3285_/D _4338_/A vssd1 vssd1 vccd1 vccd1 _3355_/D sky130_fd_sc_hd__a21o_1
X_6137_ _6223_/CLK _6137_/D vssd1 vssd1 vccd1 vccd1 _6137_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4864__A2 _4863_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4077__A0 _6462_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6068_ _4366_/A _6066_/X _6067_/Y hold440/X _6040_/Y vssd1 vssd1 vccd1 vccd1 _6068_/X
+ sky130_fd_sc_hd__o32a_1
XANTENNA__4915__S _5016_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5019_ _6262_/Q _6197_/Q _6221_/Q _6114_/Q _5100_/S0 _5100_/S1 vssd1 vssd1 vccd1
+ vccd1 _5019_/X sky130_fd_sc_hd__mux4_1
XANTENNA__3824__B1 _3795_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5600__A _5600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5746__S _6104_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4304__A1 _4313_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6057__A1 _6101_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6057__B2 _6036_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3291__B2 _3581_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5370_ _5774_/A _5370_/B _5370_/C _5370_/D vssd1 vssd1 vccd1 vccd1 _5371_/D sky130_fd_sc_hd__or4_1
X_4321_ _4318_/X _4320_/Y _4322_/B vssd1 vssd1 vccd1 vccd1 _4321_/X sky130_fd_sc_hd__a21o_1
XANTENNA__4796__A _5064_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout109 _5360_/A vssd1 vssd1 vccd1 vccd1 _5388_/A sky130_fd_sc_hd__buf_4
X_4252_ _4335_/C _5345_/C _3618_/B vssd1 vssd1 vccd1 vccd1 _4785_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_1_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3203_ _3614_/A _3193_/X _3196_/Y _3202_/X _3190_/X vssd1 vssd1 vccd1 vccd1 _3221_/A
+ sky130_fd_sc_hd__o2111a_1
XANTENNA__6048__A1 _5384_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4183_ _4182_/X hold217/X _4241_/S vssd1 vssd1 vccd1 vccd1 _6117_/D sky130_fd_sc_hd__mux2_1
X_3134_ _3614_/A _3240_/B vssd1 vssd1 vccd1 vccd1 _3305_/A sky130_fd_sc_hd__nor2_1
X_3065_ _6432_/Q vssd1 vssd1 vccd1 vccd1 _3477_/A sky130_fd_sc_hd__inv_2
XANTENNA__4735__S _5232_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5241__A1_N _6093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout153_A _4716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3967_ _3967_/A _3967_/B vssd1 vssd1 vccd1 vccd1 _5303_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_70_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4470__S _4473_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5706_ _5706_/A _5706_/B vssd1 vssd1 vccd1 vccd1 _5706_/X sky130_fd_sc_hd__or2_1
XFILLER_0_45_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3898_ _3898_/A _4444_/A _3898_/C vssd1 vssd1 vccd1 vccd1 _3901_/A sky130_fd_sc_hd__and3_1
XFILLER_0_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5637_ _5732_/A _5637_/B vssd1 vssd1 vccd1 vccd1 _5637_/X sky130_fd_sc_hd__and2_1
XFILLER_0_79_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5568_ _5567_/B _5566_/X _5567_/Y _5598_/S vssd1 vssd1 vccd1 vccd1 _5568_/X sky130_fd_sc_hd__o211a_1
Xhold152 _4532_/X vssd1 vssd1 vccd1 vccd1 _6237_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold141 _6196_/Q vssd1 vssd1 vccd1 vccd1 hold141/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_37_wb_clk_i_A clkbuf_leaf_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_4519_ _4519_/A _6003_/B vssd1 vssd1 vccd1 vccd1 _4527_/S sky130_fd_sc_hd__or2_4
Xhold130 _6204_/Q vssd1 vssd1 vccd1 vccd1 hold130/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold185 _6443_/Q vssd1 vssd1 vccd1 vccd1 hold185/X sky130_fd_sc_hd__dlygate4sd3_1
X_5499_ _5497_/X _5498_/X _5499_/S vssd1 vssd1 vccd1 vccd1 _5499_/X sky130_fd_sc_hd__mux2_1
Xhold174 _6137_/Q vssd1 vssd1 vccd1 vccd1 hold174/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold163 _6142_/Q vssd1 vssd1 vccd1 vccd1 hold163/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold196 _4370_/X vssd1 vssd1 vccd1 vccd1 _6135_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4773__A1 _3489_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4380__S _4385_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4870_ _6478_/Q _4794_/Y _4796_/Y _4863_/X _4793_/Y vssd1 vssd1 vccd1 vccd1 _4870_/X
+ sky130_fd_sc_hd__a221o_1
X_3821_ _6233_/Q _3731_/X _3810_/X _6256_/Q vssd1 vssd1 vccd1 vccd1 _3822_/C sky130_fd_sc_hd__a22o_1
XFILLER_0_39_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3752_ _6345_/Q _3752_/B vssd1 vssd1 vccd1 vccd1 _4060_/B sky130_fd_sc_hd__nand2_4
XFILLER_0_82_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3683_ _3258_/B _5146_/D _5607_/B2 vssd1 vssd1 vccd1 vccd1 _3693_/A sky130_fd_sc_hd__o21ai_1
X_6471_ _6472_/CLK _6471_/D fanout177/X vssd1 vssd1 vccd1 vccd1 hold77/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5422_ _6019_/S _5422_/B vssd1 vssd1 vccd1 vccd1 _5484_/S sky130_fd_sc_hd__or2_2
XFILLER_0_42_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5353_ _5600_/A _5337_/X _5352_/X hold604/X _5343_/X vssd1 vssd1 vccd1 vccd1 _5353_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_49_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5415__A _6434_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6010__S _6011_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4304_ _4313_/A _5418_/A _4312_/D _4312_/A vssd1 vssd1 vccd1 vccd1 _4304_/X sky130_fd_sc_hd__a31o_1
X_5284_ _6340_/Q _5160_/B _5284_/S vssd1 vssd1 vccd1 vccd1 _5284_/X sky130_fd_sc_hd__mux2_1
X_4235_ hold167/X hold153/X _4235_/S vssd1 vssd1 vccd1 vccd1 _4235_/X sky130_fd_sc_hd__mux2_1
X_4166_ _4210_/B _4166_/B vssd1 vssd1 vccd1 vccd1 _4166_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_4_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3117_ _3326_/B _4557_/C vssd1 vssd1 vccd1 vccd1 _3249_/A sky130_fd_sc_hd__nor2_1
X_4097_ _3753_/X _4095_/A _4096_/X _5136_/B vssd1 vssd1 vccd1 vccd1 _4097_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3589__B _5387_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4999_ hold93/A hold95/A _6136_/Q _6180_/Q _5404_/A0 _5100_/S1 vssd1 vssd1 vccd1
+ vccd1 _4999_/X sky130_fd_sc_hd__mux4_1
XANTENNA__4755__A1 _6314_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4755__B2 _4957_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5704__B1 _5721_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5133__A1_N _6333_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4375__S _4376_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4883__B _6365_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3499__B _5567_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout80 _3791_/X vssd1 vssd1 vccd1 vccd1 _4190_/A sky130_fd_sc_hd__buf_4
XFILLER_0_36_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4020_ _4115_/A _5262_/B vssd1 vssd1 vccd1 vccd1 _4020_/X sky130_fd_sc_hd__and2_1
XANTENNA__5889__B _5970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4682__A0 _6379_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3485__A1 _5995_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5971_ _6409_/Q _6428_/Q _5971_/S vssd1 vssd1 vccd1 vccd1 _5971_/X sky130_fd_sc_hd__mux2_1
X_4922_ _6366_/Q _6367_/Q _4922_/C vssd1 vssd1 vccd1 vccd1 _4922_/X sky130_fd_sc_hd__and3_1
XFILLER_0_59_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_30 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4853_ _6415_/Q _4930_/B vssd1 vssd1 vccd1 vccd1 _4853_/X sky130_fd_sc_hd__or2_1
X_4784_ _5346_/A _4784_/B _4784_/C _4784_/D vssd1 vssd1 vccd1 vccd1 _4785_/C sky130_fd_sc_hd__or4_1
XFILLER_0_62_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4737__A1 _6311_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4737__B2 _4957_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3804_ _3816_/B _3883_/S _3884_/S vssd1 vssd1 vccd1 vccd1 _3804_/X sky130_fd_sc_hd__and3_4
XFILLER_0_27_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6005__S _6011_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5129__B _5783_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6523_ _6529_/A vssd1 vssd1 vccd1 vccd1 _6523_/X sky130_fd_sc_hd__buf_1
X_3735_ _4438_/A vssd1 vssd1 vccd1 vccd1 _4414_/A sky130_fd_sc_hd__inv_2
XFILLER_0_42_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3960__A2 _3731_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6454_ _6454_/CLK _6454_/D vssd1 vssd1 vccd1 vccd1 _6454_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5405_ _5405_/A _5405_/B vssd1 vssd1 vccd1 vccd1 _5405_/Y sky130_fd_sc_hd__nand2_1
X_3666_ _3704_/B _6021_/S vssd1 vssd1 vccd1 vccd1 _6443_/D sky130_fd_sc_hd__and2_1
XANTENNA_fanout116_A _5581_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3173__A0 _4782_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3597_ _5362_/A _5866_/C vssd1 vssd1 vccd1 vccd1 _3597_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_62_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6385_ _6462_/CLK _6385_/D vssd1 vssd1 vccd1 vccd1 _6385_/Q sky130_fd_sc_hd__dfxtp_4
X_5336_ _5336_/A _5336_/B vssd1 vssd1 vccd1 vccd1 _5336_/X sky130_fd_sc_hd__or2_1
X_5267_ _5267_/A _5267_/B _5267_/C _5267_/D vssd1 vssd1 vccd1 vccd1 _5267_/X sky130_fd_sc_hd__or4_1
X_4218_ _5605_/A _6290_/Q _3115_/Y _4217_/X vssd1 vssd1 vccd1 vccd1 _4218_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4899__S1 _5100_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5799__B _6459_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5198_ _6384_/Q _4332_/B _4022_/B _6381_/Q vssd1 vssd1 vccd1 vccd1 _5199_/C sky130_fd_sc_hd__a22o_1
XFILLER_0_97_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4149_ _4149_/A _4149_/B vssd1 vssd1 vccd1 vccd1 _5304_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_97_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5754__S _6104_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6102__B1 _6107_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5000__S1 _5078_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5929__S _6021_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3520_ _5384_/A hold59/X _3519_/Y vssd1 vssd1 vccd1 vccd1 hold60/A sky130_fd_sc_hd__a21o_1
XFILLER_0_97_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4788__B _4788_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3942__A2 _6081_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3451_ _3431_/B _3441_/Y _3450_/X _5995_/C vssd1 vssd1 vccd1 vccd1 _3464_/C sky130_fd_sc_hd__a31o_1
XFILLER_0_12_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3382_ _3405_/A _3671_/B vssd1 vssd1 vccd1 vccd1 _3382_/Y sky130_fd_sc_hd__nand2_1
X_6170_ _6237_/CLK hold66/X vssd1 vssd1 vccd1 vccd1 hold65/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__5695__A2 _5721_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4804__A_N _5322_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5121_ _6347_/Q _5294_/B _4223_/A vssd1 vssd1 vccd1 vccd1 _5151_/B sky130_fd_sc_hd__a21o_2
XANTENNA__3912__S _4241_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3458__A1 _5607_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5052_ _6406_/Q _5051_/X _5971_/S vssd1 vssd1 vccd1 vccd1 _5052_/X sky130_fd_sc_hd__mux2_1
X_4003_ _4150_/A _4005_/A vssd1 vssd1 vccd1 vccd1 _4003_/X sky130_fd_sc_hd__or2_1
XFILLER_0_79_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3213__A _5605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4407__B1 _5731_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5954_ _5954_/A _5954_/B vssd1 vssd1 vccd1 vccd1 _5954_/X sky130_fd_sc_hd__xor2_1
XANTENNA__6524__A _6529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3630__A1 _3489_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5885_ _5884_/A _5884_/B _5884_/C vssd1 vssd1 vccd1 vccd1 _5890_/B sky130_fd_sc_hd__a21oi_1
X_4905_ _6366_/Q _4922_/C vssd1 vssd1 vccd1 vccd1 _4905_/Y sky130_fd_sc_hd__nand2_1
X_4836_ _5817_/A _4834_/X _4835_/Y _5771_/A vssd1 vssd1 vccd1 vccd1 _4836_/X sky130_fd_sc_hd__a211o_1
XANTENNA__5907__A0 _6459_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5058__S1 _5100_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4186__A2 _3793_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4767_ _6316_/Q _4719_/A _4766_/X _4957_/S vssd1 vssd1 vccd1 vccd1 _4767_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_7_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3933__A2 _6286_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4698_ _6284_/Q _4697_/X _4712_/S vssd1 vssd1 vccd1 vccd1 _4698_/X sky130_fd_sc_hd__mux2_1
X_3718_ _3717_/A _3717_/B _6377_/Q vssd1 vssd1 vccd1 vccd1 _3718_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_43_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5135__A1 _5268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6437_ _6439_/CLK _6437_/D fanout178/X vssd1 vssd1 vccd1 vccd1 _6437_/Q sky130_fd_sc_hd__dfrtp_1
X_3649_ _5295_/A _3640_/C hold622/X vssd1 vssd1 vccd1 vccd1 _3650_/C sky130_fd_sc_hd__o21ba_1
XFILLER_0_30_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6368_ _6475_/CLK _6368_/D fanout181/X vssd1 vssd1 vccd1 vccd1 _6368_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_87_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5319_ _5323_/B _3281_/X _5323_/C _5318_/X _5607_/B2 vssd1 vssd1 vccd1 vccd1 _5319_/X
+ sky130_fd_sc_hd__o41a_1
XFILLER_0_11_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6299_ _6446_/CLK _6299_/D fanout184/X vssd1 vssd1 vccd1 vccd1 _6299_/Q sky130_fd_sc_hd__dfrtp_4
Xhold23 hold23/A vssd1 vssd1 vccd1 vccd1 hold23/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold12 hold12/A vssd1 vssd1 vccd1 vccd1 hold12/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 hold45/A vssd1 vssd1 vccd1 vccd1 hold45/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 hold56/A vssd1 vssd1 vccd1 vccd1 hold56/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 hold34/A vssd1 vssd1 vccd1 vccd1 hold34/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 hold78/A vssd1 vssd1 vccd1 vccd1 hold78/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 hold67/A vssd1 vssd1 vccd1 vccd1 hold67/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold89 hold89/A vssd1 vssd1 vccd1 vccd1 hold89/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5749__S _6104_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3924__A2 _6285_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_9 _5317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5126__A1 _4716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_18 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4980__S0 _5100_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xci2406_z80_202 vssd1 vssd1 vccd1 vccd1 ci2406_z80_202/HI io_oeb[17] sky130_fd_sc_hd__conb_1
XFILLER_0_16_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xci2406_z80_213 vssd1 vssd1 vccd1 vccd1 ci2406_z80_213/HI io_out[35] sky130_fd_sc_hd__conb_1
XANTENNA__5659__S _5734_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3612__A1 _3205_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5670_ _3956_/X _5655_/B _5667_/X _5669_/X vssd1 vssd1 vccd1 vccd1 _5670_/X sky130_fd_sc_hd__o22a_1
Xclkbuf_leaf_32_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6409_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__5365__A1 _5600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4621_ _3859_/B _4036_/B _4641_/B vssd1 vssd1 vccd1 vccd1 _4621_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_37_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4552_ _4138_/X hold208/X _4554_/S vssd1 vssd1 vccd1 vccd1 _6264_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_25_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold526 _6444_/Q vssd1 vssd1 vccd1 vccd1 hold526/X sky130_fd_sc_hd__buf_2
Xhold515 _4568_/X vssd1 vssd1 vccd1 vccd1 _6275_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3503_ _3503_/A _3503_/B vssd1 vssd1 vccd1 vccd1 _3503_/Y sky130_fd_sc_hd__nand2_1
Xhold504 _6331_/Q vssd1 vssd1 vccd1 vccd1 hold504/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4483_ _4546_/A _4501_/A vssd1 vssd1 vccd1 vccd1 _4491_/S sky130_fd_sc_hd__or2_4
X_3434_ _3632_/D _3434_/B vssd1 vssd1 vccd1 vccd1 _3434_/Y sky130_fd_sc_hd__nor2_1
Xhold548 _6290_/Q vssd1 vssd1 vccd1 vccd1 hold548/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3208__A _3304_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold559 _6000_/X vssd1 vssd1 vccd1 vccd1 _6442_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold537 _6428_/Q vssd1 vssd1 vccd1 vccd1 _5969_/A sky130_fd_sc_hd__clkdlybuf4s25_1
X_6222_ _6263_/CLK _6222_/D vssd1 vssd1 vccd1 vccd1 _6222_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5668__A2 _5721_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4876__B1 _6070_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3365_ _4338_/B _3364_/Y _6340_/Q vssd1 vssd1 vccd1 vccd1 _3370_/B sky130_fd_sc_hd__mux2_1
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5423__A _5485_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6153_ _6490_/CLK hold94/X vssd1 vssd1 vccd1 vccd1 hold93/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4738__S _4768_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3296_ _5314_/S _4338_/B vssd1 vssd1 vccd1 vccd1 _3296_/Y sky130_fd_sc_hd__nand2_1
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6084_ _6101_/A _6083_/X _6107_/S vssd1 vssd1 vccd1 vccd1 _6084_/X sky130_fd_sc_hd__o21a_1
X_5104_ _6490_/Q _5104_/A2 _5103_/X vssd1 vssd1 vccd1 vccd1 _5104_/X sky130_fd_sc_hd__a21o_1
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5035_ _6461_/Q _5034_/X _5974_/S vssd1 vssd1 vccd1 vccd1 _5035_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_79_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout183_A fanout185/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4473__S _4473_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3597__B _5866_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5937_ _5937_/A _5937_/B vssd1 vssd1 vccd1 vccd1 _5937_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_75_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5868_ _5870_/A vssd1 vssd1 vccd1 vccd1 _5884_/A sky130_fd_sc_hd__inv_2
XANTENNA__4159__A2 _6290_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5356__A1 _4248_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4819_ hold83/A hold63/A _6187_/Q hold79/A _5078_/S1 _5404_/A0 vssd1 vssd1 vccd1
+ vccd1 _4819_/X sky130_fd_sc_hd__mux4_1
X_5799_ _5866_/A _6459_/Q _5866_/C vssd1 vssd1 vccd1 vccd1 _5800_/C sky130_fd_sc_hd__or3_1
XFILLER_0_7_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5317__B _5317_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3118__A _4268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput24 _6528_/X vssd1 vssd1 vccd1 vccd1 io_oeb[27] sky130_fd_sc_hd__buf_12
XFILLER_0_101_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput46 _6308_/Q vssd1 vssd1 vccd1 vccd1 io_out[27] sky130_fd_sc_hd__buf_12
XANTENNA_fanout96_A _3297_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput35 _6328_/Q vssd1 vssd1 vccd1 vccd1 io_out[17] sky130_fd_sc_hd__buf_12
Xoutput57 _6319_/Q vssd1 vssd1 vccd1 vccd1 io_out[8] sky130_fd_sc_hd__buf_12
XANTENNA__5292__A0 _4227_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5831__A2 _5974_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4383__S _4385_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5044__A0 _6425_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5347__A1 _4273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4131__B _4131_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5942__S _5975_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3150_ _5315_/A _3322_/C _3281_/A vssd1 vssd1 vccd1 vccd1 _4247_/A sky130_fd_sc_hd__and3_1
X_3081_ _3081_/A vssd1 vssd1 vccd1 vccd1 _3928_/A sky130_fd_sc_hd__inv_2
XFILLER_0_89_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3698__A _5478_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4181__S1 _5721_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5035__A0 _6461_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3983_ _6380_/Q _6384_/Q _6343_/Q vssd1 vssd1 vccd1 vccd1 _5267_/C sky130_fd_sc_hd__mux2_1
XFILLER_0_9_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5722_ _5722_/A _5722_/B vssd1 vssd1 vccd1 vccd1 _5722_/X sky130_fd_sc_hd__or2_1
XFILLER_0_84_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5338__A1 _4675_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5653_ _5653_/A _5653_/B vssd1 vssd1 vccd1 vccd1 _5653_/X sky130_fd_sc_hd__and2_2
XANTENNA__6307__RESET_B fanout183/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5418__A _5418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6013__S _6019_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5584_ _5594_/A _5584_/B vssd1 vssd1 vccd1 vccd1 _5585_/B sky130_fd_sc_hd__nor2_1
XANTENNA__4322__A _5581_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4604_ _5767_/A _4605_/B _4605_/C _4641_/B vssd1 vssd1 vccd1 vccd1 _4604_/X sky130_fd_sc_hd__and4_2
Xhold301 hold661/X vssd1 vssd1 vccd1 vccd1 _3493_/C sky130_fd_sc_hd__buf_1
X_4535_ hold51/X _4456_/X _4536_/S vssd1 vssd1 vccd1 vccd1 hold52/A sky130_fd_sc_hd__mux2_1
Xhold334 _6302_/Q vssd1 vssd1 vccd1 vccd1 hold334/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold312 _6307_/Q vssd1 vssd1 vccd1 vccd1 hold312/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_27_wb_clk_i_A clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold323 _5396_/X vssd1 vssd1 vccd1 vccd1 _6356_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold378 _4365_/X vssd1 vssd1 vccd1 vccd1 _6128_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4849__B1 _4924_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold345 _4317_/X vssd1 vssd1 vccd1 vccd1 _6125_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4466_ hold268/X _3911_/X _4473_/S vssd1 vssd1 vccd1 vccd1 _4466_/X sky130_fd_sc_hd__mux2_1
Xhold356 _4878_/X vssd1 vssd1 vccd1 vccd1 _6320_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold367 _6318_/Q vssd1 vssd1 vccd1 vccd1 hold367/X sky130_fd_sc_hd__dlygate4sd3_1
X_3417_ _3400_/X _3440_/A _3408_/X _3416_/X _5522_/A vssd1 vssd1 vccd1 vccd1 _3417_/X
+ sky130_fd_sc_hd__o41a_1
Xhold389 _6434_/Q vssd1 vssd1 vccd1 vccd1 _4363_/A sky130_fd_sc_hd__buf_2
XFILLER_0_68_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5510__A1 _4668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6205_ _6237_/CLK _6205_/D vssd1 vssd1 vccd1 vccd1 _6205_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4468__S _4473_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4397_ hold139/X _4240_/X _4397_/S vssd1 vssd1 vccd1 vccd1 _4397_/X sky130_fd_sc_hd__mux2_1
X_3348_ _4792_/A _4802_/C vssd1 vssd1 vccd1 vccd1 _3386_/A sky130_fd_sc_hd__or2_1
X_6136_ _6263_/CLK _6136_/D vssd1 vssd1 vccd1 vccd1 _6136_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3279_ _3639_/C _4325_/C vssd1 vssd1 vccd1 vccd1 _4264_/B sky130_fd_sc_hd__nor2_2
X_6067_ _6067_/A _6071_/S vssd1 vssd1 vccd1 vccd1 _6067_/Y sky130_fd_sc_hd__nor2_1
X_5018_ hold73/A _6145_/Q _6137_/Q _6181_/Q _5100_/S0 _5100_/S1 vssd1 vssd1 vccd1
+ vccd1 _5018_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_67_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3120__B _3172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5762__S _5765_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4304__A2 _5418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4378__S _4385_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5063__A _5102_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6057__A2 _4881_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3910__S1 _5721_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5568__A1 _5567_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4240__B2 _4441_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3981__A _6285_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4320_ _4320_/A _4320_/B vssd1 vssd1 vccd1 vccd1 _4320_/Y sky130_fd_sc_hd__nand2_1
X_4251_ _4338_/B _4251_/B vssd1 vssd1 vccd1 vccd1 _5336_/A sky130_fd_sc_hd__nor2_1
X_3202_ _6430_/Q _4325_/C _4248_/C _4338_/A _6435_/Q vssd1 vssd1 vccd1 vccd1 _3202_/X
+ sky130_fd_sc_hd__a311o_1
XANTENNA__3205__B _3205_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4182_ _4179_/X _4180_/X _4181_/X _4441_/S vssd1 vssd1 vccd1 vccd1 _4182_/X sky130_fd_sc_hd__a22o_2
X_3133_ _3205_/B _3639_/C vssd1 vssd1 vccd1 vccd1 _3240_/B sky130_fd_sc_hd__or2_2
X_3064_ _3064_/A vssd1 vssd1 vccd1 vccd1 _3368_/S sky130_fd_sc_hd__inv_2
XFILLER_0_54_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5008__A0 _6460_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6008__S _6011_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5559__A1 _5041_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4036__B _4036_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4751__S _5289_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3966_ _4045_/B _3966_/B _3966_/C vssd1 vssd1 vccd1 vccd1 _3967_/B sky130_fd_sc_hd__and3_1
XFILLER_0_57_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5705_ _6175_/Q _5721_/A2 _5721_/B1 _6254_/Q _5721_/C1 vssd1 vssd1 vccd1 vccd1 _5706_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_18_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5636_ _6178_/Q _5721_/A2 _4235_/S _6134_/Q _5730_/C1 vssd1 vssd1 vccd1 vccd1 _5639_/C
+ sky130_fd_sc_hd__a221o_1
X_3897_ _4444_/A _3898_/C vssd1 vssd1 vccd1 vccd1 _4451_/B sky130_fd_sc_hd__and2_1
XFILLER_0_60_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5582__S _5593_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5567_ _5567_/A _5567_/B vssd1 vssd1 vccd1 vccd1 _5567_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__3181__D_N _3168_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold120 hold659/X vssd1 vssd1 vccd1 vccd1 _3704_/B sky130_fd_sc_hd__buf_1
X_5498_ hold590/X input9/X _5510_/S vssd1 vssd1 vccd1 vccd1 _5498_/X sky130_fd_sc_hd__mux2_1
Xhold142 _4486_/X vssd1 vssd1 vccd1 vccd1 _6196_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold153 _6266_/Q vssd1 vssd1 vccd1 vccd1 hold153/X sky130_fd_sc_hd__dlygate4sd3_1
X_4518_ _4240_/X hold242/X _4518_/S vssd1 vssd1 vccd1 vccd1 _4518_/X sky130_fd_sc_hd__mux2_1
Xhold131 _4495_/X vssd1 vssd1 vccd1 vccd1 _6204_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold186 _3654_/X vssd1 vssd1 vccd1 vccd1 _3655_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold164 _4378_/X vssd1 vssd1 vccd1 vccd1 _6142_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold175 _4372_/X vssd1 vssd1 vccd1 vccd1 _6137_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4449_ hold263/X _4448_/X _4464_/S vssd1 vssd1 vccd1 vccd1 _6175_/D sky130_fd_sc_hd__mux2_1
XANTENNA__4298__A1 _6310_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold197 _6206_/Q vssd1 vssd1 vccd1 vccd1 hold197/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_95_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5247__A0 _6383_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6119_ _6412_/CLK hold6/X vssd1 vssd1 vccd1 vccd1 hold5/A sky130_fd_sc_hd__dfxtp_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4926__S _4948_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3131__A _3205_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3820_ _6456_/Q _3804_/X _3807_/X _6177_/Q vssd1 vssd1 vccd1 vccd1 _3822_/B sky130_fd_sc_hd__a22o_1
X_3751_ _6345_/Q _3752_/B vssd1 vssd1 vccd1 vccd1 _4156_/A sky130_fd_sc_hd__and2_2
XFILLER_0_82_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3682_ _3352_/B _3691_/B _5387_/C _3786_/A vssd1 vssd1 vccd1 vccd1 _3682_/X sky130_fd_sc_hd__a211o_1
X_6470_ _6470_/CLK _6470_/D fanout177/X vssd1 vssd1 vccd1 vccd1 _6470_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5421_ _6458_/Q _5420_/X _5512_/S vssd1 vssd1 vccd1 vccd1 _5421_/X sky130_fd_sc_hd__mux2_1
X_5352_ _6300_/Q _3428_/B _5314_/X _3511_/A _5351_/X vssd1 vssd1 vccd1 vccd1 _5352_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_2_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5415__B _6469_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4303_ _4303_/A _6121_/Q _4303_/C vssd1 vssd1 vccd1 vccd1 _4312_/D sky130_fd_sc_hd__and3_1
X_5283_ _3064_/A _5282_/Y _5489_/S vssd1 vssd1 vccd1 vccd1 _6339_/D sky130_fd_sc_hd__mux2_1
X_4234_ hold121/X _5721_/B1 _5721_/C1 _4233_/X vssd1 vssd1 vccd1 vccd1 _4234_/X sky130_fd_sc_hd__o211a_1
X_4165_ _4212_/A _4210_/A vssd1 vssd1 vccd1 vccd1 _4166_/B sky130_fd_sc_hd__nor2_1
XANTENNA__4746__S _4770_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6527__A _6529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3116_ _4268_/A _4273_/A vssd1 vssd1 vccd1 vccd1 _4557_/C sky130_fd_sc_hd__or2_4
X_4096_ _4150_/A _4096_/B vssd1 vssd1 vccd1 vccd1 _4096_/X sky130_fd_sc_hd__or2_1
XFILLER_0_77_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4481__S _4482_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4998_ _4997_/X hold336/X _5098_/S vssd1 vssd1 vccd1 vccd1 _4998_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_92_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3949_ _4052_/A _4600_/A _3902_/Y vssd1 vssd1 vccd1 vccd1 _3950_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_73_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5619_ _5619_/A _5619_/B vssd1 vssd1 vccd1 vccd1 _5619_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__3715__B1 _4948_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4140__B1 _3795_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold642_A _6312_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5341__A _5605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5487__S _5567_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4391__S _4397_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3796__A _3852_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout70 _3886_/S vssd1 vssd1 vccd1 vccd1 _3884_/S sky130_fd_sc_hd__clkbuf_8
Xfanout81 _3791_/X vssd1 vssd1 vccd1 vccd1 _3892_/A sky130_fd_sc_hd__buf_2
XFILLER_0_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4682__A1 _6285_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5970_ _5970_/A _5970_/B vssd1 vssd1 vccd1 vccd1 _5970_/Y sky130_fd_sc_hd__xnor2_1
X_4921_ _6367_/Q _4790_/X _4789_/B vssd1 vssd1 vccd1 vccd1 _4921_/X sky130_fd_sc_hd__a21o_1
XANTENNA__5631__B1 _5610_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4852_ _4852_/A _4852_/B _4852_/C vssd1 vssd1 vccd1 vccd1 _4852_/X sky130_fd_sc_hd__or3_1
XFILLER_0_19_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3803_ _6151_/Q _4528_/A _4474_/A _6142_/Q _3797_/X vssd1 vssd1 vccd1 vccd1 _3813_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_28_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4783_ _5322_/A _5146_/D _4803_/B _4782_/X vssd1 vssd1 vccd1 vccd1 _5422_/B sky130_fd_sc_hd__or4b_2
XFILLER_0_82_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3734_ _3665_/A _6468_/Q _3624_/Y _3694_/X vssd1 vssd1 vccd1 vccd1 _3734_/X sky130_fd_sc_hd__o211a_2
XFILLER_0_42_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3945__B1 _3807_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3665_ _3665_/A _3665_/B vssd1 vssd1 vccd1 vccd1 _6163_/D sky130_fd_sc_hd__or2_2
X_6453_ _6454_/CLK _6453_/D vssd1 vssd1 vccd1 vccd1 _6453_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__6021__S _6021_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5404_ _5404_/A0 _5403_/Y _5513_/S vssd1 vssd1 vccd1 vccd1 _6360_/D sky130_fd_sc_hd__mux2_1
X_3596_ _3632_/D _3561_/Y _3619_/C _3433_/B vssd1 vssd1 vccd1 vccd1 _5866_/C sky130_fd_sc_hd__o2bb2a_4
X_6384_ _6384_/CLK _6384_/D vssd1 vssd1 vccd1 vccd1 _6384_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_11_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5335_ _5757_/B hold619/X _5331_/X _5368_/S vssd1 vssd1 vccd1 vccd1 _6343_/D sky130_fd_sc_hd__a22o_1
X_5266_ _5322_/A _5264_/X _5265_/Y vssd1 vssd1 vccd1 vccd1 _5266_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_55_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4217_ _4217_/A _6284_/Q vssd1 vssd1 vccd1 vccd1 _4217_/X sky130_fd_sc_hd__and2_1
XFILLER_0_76_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4476__S _4482_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5799__C _5866_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5197_ _6383_/Q _4116_/A _3760_/Y _6378_/Q vssd1 vssd1 vccd1 vccd1 _5199_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_97_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4148_ _4132_/B _4134_/B _4130_/A vssd1 vssd1 vccd1 vccd1 _4149_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_78_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4079_ _4227_/S _4077_/X _4078_/X vssd1 vssd1 vccd1 vccd1 _6093_/A sky130_fd_sc_hd__a21oi_4
XFILLER_0_93_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5925__A1 _6424_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_hold592_A _6368_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3872__C1 _3852_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4416__A1 _4441_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5916__A1 _6423_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5392__A2 _6023_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4150__A _4150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3450_ _5146_/C _3450_/B vssd1 vssd1 vccd1 vccd1 _3450_/X sky130_fd_sc_hd__or2_1
X_3381_ _6431_/Q _3370_/A _3370_/B _3370_/C _3673_/B vssd1 vssd1 vccd1 vccd1 _3671_/B
+ sky130_fd_sc_hd__a41o_2
X_5120_ hold617/X _5294_/B _4223_/A vssd1 vssd1 vccd1 vccd1 _5290_/S sky130_fd_sc_hd__a21oi_4
XFILLER_0_20_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5051_ _6425_/Q _4793_/Y _5043_/X _5050_/X vssd1 vssd1 vccd1 vccd1 _5051_/X sky130_fd_sc_hd__a211o_1
XANTENNA__4655__A1 _3168_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4002_ _4004_/B _4004_/C _6287_/Q vssd1 vssd1 vccd1 vccd1 _4005_/A sky130_fd_sc_hd__o21a_1
XANTENNA__3213__B _3281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5953_ _5937_/A _5937_/B _5934_/A vssd1 vssd1 vccd1 vccd1 _5954_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_1_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4325__A _4325_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6016__S _6019_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4904_ _4901_/B _4903_/X _4948_/S vssd1 vssd1 vccd1 vccd1 _4904_/X sky130_fd_sc_hd__mux2_1
X_5884_ _5884_/A _5884_/B _5884_/C vssd1 vssd1 vccd1 vccd1 _5886_/A sky130_fd_sc_hd__and3_1
XFILLER_0_90_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4835_ _5817_/A _4835_/B vssd1 vssd1 vccd1 vccd1 _4835_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_7_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4766_ _6316_/Q _4720_/X _5224_/A2 hold434/X vssd1 vssd1 vccd1 vccd1 _4766_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_43_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3717_ _3717_/A _3717_/B vssd1 vssd1 vccd1 vccd1 _3717_/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_70_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4697_ _6382_/Q _6378_/Q _4711_/S vssd1 vssd1 vccd1 vccd1 _4697_/X sky130_fd_sc_hd__mux2_1
X_6436_ _6470_/CLK _6436_/D fanout178/X vssd1 vssd1 vccd1 vccd1 _6436_/Q sky130_fd_sc_hd__dfrtp_4
X_3648_ hold298/X _3648_/B _3648_/C vssd1 vssd1 vccd1 vccd1 _3650_/B sky130_fd_sc_hd__and3b_1
XFILLER_0_3_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3579_ _4263_/A _3573_/X _3574_/X _3578_/X vssd1 vssd1 vccd1 vccd1 _6529_/A sky130_fd_sc_hd__a31o_4
X_6367_ _6475_/CLK _6367_/D fanout175/X vssd1 vssd1 vccd1 vccd1 _6367_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_3_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5318_ _5323_/D _5316_/Y _5317_/Y _5605_/C vssd1 vssd1 vccd1 vccd1 _5318_/X sky130_fd_sc_hd__o31a_1
X_6298_ _6446_/CLK _6298_/D fanout184/X vssd1 vssd1 vccd1 vccd1 _6298_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__6096__B1 _6107_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold13 hold13/A vssd1 vssd1 vccd1 vccd1 hold13/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3404__A _5777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold35 hold35/A vssd1 vssd1 vccd1 vccd1 hold35/X sky130_fd_sc_hd__dlygate4sd3_1
X_5249_ _6338_/Q _5202_/A _5247_/X _3774_/A _5248_/X vssd1 vssd1 vccd1 vccd1 _5249_/X
+ sky130_fd_sc_hd__a221o_1
Xhold46 hold46/A vssd1 vssd1 vccd1 vccd1 hold46/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_2_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6449_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold24 hold24/A vssd1 vssd1 vccd1 vccd1 hold24/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold57 hold57/A vssd1 vssd1 vccd1 vccd1 hold57/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 hold79/A vssd1 vssd1 vccd1 vccd1 hold79/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold68 hold68/A vssd1 vssd1 vccd1 vccd1 hold68/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3123__B _3168_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5071__A1 _6426_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5765__S _5765_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3793__B _3885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3924__A3 _6379_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5126__A2 _6333_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4980__S1 _5100_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5005__S _5105_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4129__B _4131_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xci2406_z80_203 vssd1 vssd1 vccd1 vccd1 ci2406_z80_203/HI io_oeb[18] sky130_fd_sc_hd__conb_1
XANTENNA__4844__S _5101_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3968__B _6380_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xci2406_z80_214 vssd1 vssd1 vccd1 vccd1 io_oeb[4] ci2406_z80_214/LO sky130_fd_sc_hd__conb_1
XFILLER_0_69_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4620_ _5393_/A1 hold529/X _4582_/Y _4619_/X vssd1 vssd1 vccd1 vccd1 _4620_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_44_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4551_ _4085_/X hold204/X _4554_/S vssd1 vssd1 vccd1 vccd1 _4551_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_12_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold527 _6276_/Q vssd1 vssd1 vccd1 vccd1 hold527/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold516 _6469_/Q vssd1 vssd1 vccd1 vccd1 _5410_/A sky130_fd_sc_hd__clkbuf_2
X_3502_ _5567_/B _6019_/S hold526/X vssd1 vssd1 vccd1 vccd1 _3503_/B sky130_fd_sc_hd__a21oi_4
Xhold505 _5098_/X vssd1 vssd1 vccd1 vccd1 _6331_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4482_ hold215/X _4463_/X _4482_/S vssd1 vssd1 vccd1 vccd1 _4482_/X sky130_fd_sc_hd__mux2_1
X_3433_ _4344_/A _3433_/B vssd1 vssd1 vccd1 vccd1 _3434_/B sky130_fd_sc_hd__nand2_1
Xhold549 _4640_/X vssd1 vssd1 vccd1 vccd1 _6290_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold538 _5977_/X vssd1 vssd1 vccd1 vccd1 _6428_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6221_ _6223_/CLK _6221_/D vssd1 vssd1 vccd1 vccd1 _6221_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6152_ _6376_/CLK _6152_/D vssd1 vssd1 vccd1 vccd1 _6152_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4876__A1 _6364_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3364_ _4217_/A _3511_/A _3986_/A vssd1 vssd1 vccd1 vccd1 _3364_/Y sky130_fd_sc_hd__nand3_2
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5103_ _6316_/Q _4963_/B _5102_/B _4796_/Y vssd1 vssd1 vccd1 vccd1 _5103_/X sky130_fd_sc_hd__a22o_1
X_3295_ _4217_/A _3511_/A _3986_/A vssd1 vssd1 vccd1 vccd1 _4338_/B sky130_fd_sc_hd__nand3b_4
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6083_ _6101_/B _5002_/B _5545_/Y _6036_/X vssd1 vssd1 vccd1 vccd1 _6083_/X sky130_fd_sc_hd__o22a_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5034_ _5964_/A _5033_/X _5021_/Y vssd1 vssd1 vccd1 vccd1 _5034_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_73_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3851__A2 _3884_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout176_A input18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5936_ _5914_/A _5914_/C _5924_/A _5935_/Y vssd1 vssd1 vccd1 vccd1 _5937_/B sky130_fd_sc_hd__o31a_1
XFILLER_0_48_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5867_ _6419_/Q _5867_/B _5867_/C vssd1 vssd1 vccd1 vccd1 _5870_/A sky130_fd_sc_hd__and3_1
XANTENNA__4159__A3 _6384_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5356__A2 _5360_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5798_ _5817_/A _5797_/X _4835_/Y _5771_/A vssd1 vssd1 vccd1 vccd1 _5798_/X sky130_fd_sc_hd__a211o_1
X_4818_ _6362_/Q _4790_/X _4789_/B vssd1 vssd1 vccd1 vccd1 _4818_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_28_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4749_ _6313_/Q _4719_/A _4748_/X _4957_/S vssd1 vssd1 vccd1 vccd1 _4749_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_71_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3118__B _4273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput25 _6529_/X vssd1 vssd1 vccd1 vccd1 io_oeb[28] sky130_fd_sc_hd__buf_12
X_6419_ _6419_/CLK _6419_/D fanout173/X vssd1 vssd1 vccd1 vccd1 _6419_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_31_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput47 _6302_/Q vssd1 vssd1 vccd1 vccd1 io_out[28] sky130_fd_sc_hd__buf_12
Xoutput36 _6329_/Q vssd1 vssd1 vccd1 vccd1 io_out[18] sky130_fd_sc_hd__buf_12
Xoutput58 _6317_/Q vssd1 vssd1 vccd1 vccd1 io_out[9] sky130_fd_sc_hd__buf_12
XFILLER_0_31_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout89_A _4418_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3300__C _3632_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3080_ _6286_/Q vssd1 vssd1 vccd1 vccd1 _3080_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_89_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3982_ _3982_/A _3982_/B vssd1 vssd1 vccd1 vccd1 _5260_/B sky130_fd_sc_hd__xnor2_2
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5721_ _6140_/Q _5721_/A2 _5721_/B1 _6184_/Q _5721_/C1 vssd1 vssd1 vccd1 vccd1 _5722_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_72_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5652_ _5757_/B hold489/X _5611_/Y _5651_/X vssd1 vssd1 vccd1 vccd1 _5652_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_60_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5583_ _5594_/A _5584_/B vssd1 vssd1 vccd1 vccd1 _5585_/A sky130_fd_sc_hd__and2_1
XANTENNA__4322__B _4322_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4603_ _4401_/B _4641_/B _4600_/Y _4602_/Y vssd1 vssd1 vccd1 vccd1 _4603_/X sky130_fd_sc_hd__o211a_1
Xhold302 _3483_/X vssd1 vssd1 vccd1 vccd1 _6248_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4534_ hold132/X _4448_/X _4536_/S vssd1 vssd1 vccd1 vccd1 _4534_/X sky130_fd_sc_hd__mux2_1
Xhold335 _4685_/X vssd1 vssd1 vccd1 vccd1 _6302_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold313 _4710_/X vssd1 vssd1 vccd1 vccd1 _6307_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold324 _6122_/Q vssd1 vssd1 vccd1 vccd1 _4303_/C sky130_fd_sc_hd__buf_1
XFILLER_0_13_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold346 _6359_/Q vssd1 vssd1 vccd1 vccd1 hold346/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4465_ _4546_/A _4537_/A vssd1 vssd1 vccd1 vccd1 _4473_/S sky130_fd_sc_hd__nor2_4
Xhold357 _6418_/Q vssd1 vssd1 vccd1 vccd1 _5852_/A sky130_fd_sc_hd__buf_1
Xhold368 _4840_/X vssd1 vssd1 vccd1 vccd1 _6318_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3416_ _3409_/Y _3410_/Y _3411_/Y _3415_/X vssd1 vssd1 vccd1 vccd1 _3416_/X sky130_fd_sc_hd__a211o_1
X_4396_ hold116/X _4182_/X _4397_/S vssd1 vssd1 vccd1 vccd1 _4396_/X sky130_fd_sc_hd__mux2_1
X_6204_ _6456_/CLK _6204_/D vssd1 vssd1 vccd1 vccd1 _6204_/Q sky130_fd_sc_hd__dfxtp_1
Xhold379 _6417_/Q vssd1 vssd1 vccd1 vccd1 hold379/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3521__A1 _5617_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3347_ _3298_/X _3346_/X _3341_/X _3336_/A vssd1 vssd1 vccd1 vccd1 _4802_/C sky130_fd_sc_hd__o211a_2
X_6135_ _6399_/CLK _6135_/D vssd1 vssd1 vccd1 vccd1 _6135_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6066_ _6101_/A _6065_/X _6071_/S vssd1 vssd1 vccd1 vccd1 _6066_/X sky130_fd_sc_hd__o21a_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3278_ _3278_/A _3278_/B vssd1 vssd1 vccd1 vccd1 _3285_/B sky130_fd_sc_hd__nor2_1
X_5017_ _5016_/X hold387/X _5098_/S vssd1 vssd1 vccd1 vccd1 _5017_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4484__S _4491_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3824__A2 _3793_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3401__B _3489_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3120__C _4782_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5919_ _5002_/Y _5918_/Y _5771_/A vssd1 vssd1 vccd1 vccd1 _5919_/X sky130_fd_sc_hd__a21o_1
XANTENNA__4880__S0 _5100_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5609__A _5610_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4232__B _4463_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5265__A1 _5322_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3799__A _3884_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4394__S _4397_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3981__B _6286_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5864__B1_N _5887_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4250_ _5388_/B _5362_/C vssd1 vssd1 vccd1 vccd1 _4250_/X sky130_fd_sc_hd__or2_1
XFILLER_0_10_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3201_ _5995_/C _3786_/A vssd1 vssd1 vccd1 vccd1 _3426_/B sky130_fd_sc_hd__nor2_1
X_4181_ hold138/X hold114/X hold128/X hold116/X _5721_/C1 _5721_/B1 vssd1 vssd1 vccd1
+ vccd1 _4181_/X sky130_fd_sc_hd__mux4_2
X_3132_ _4675_/A _3639_/C vssd1 vssd1 vccd1 vccd1 _3642_/C sky130_fd_sc_hd__nor2_1
X_3063_ _4324_/B vssd1 vssd1 vccd1 vccd1 _5315_/B sky130_fd_sc_hd__inv_2
XANTENNA__6085__A _6085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3965_ _3966_/B _3966_/C _4045_/B vssd1 vssd1 vccd1 vccd1 _3967_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_70_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5429__A _5492_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4862__S0 _5404_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5704_ _6454_/Q _5721_/A2 _5721_/B1 _6231_/Q _5730_/C1 vssd1 vssd1 vccd1 vccd1 _5706_/A
+ sky130_fd_sc_hd__o221a_1
X_3896_ _4437_/B _4437_/A vssd1 vssd1 vccd1 vccd1 _3898_/C sky130_fd_sc_hd__and2b_1
XFILLER_0_45_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5635_ _6111_/Q _5721_/A2 _4235_/S _6218_/Q _5731_/C1 vssd1 vssd1 vccd1 vccd1 _5639_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_85_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5566_ _6373_/Q _5520_/B _5565_/Y _5485_/S vssd1 vssd1 vccd1 vccd1 _5566_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_13_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold110 _4390_/X vssd1 vssd1 vccd1 vccd1 _6151_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5731__A2 _4406_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold143 _6470_/Q vssd1 vssd1 vccd1 vccd1 _3700_/A sky130_fd_sc_hd__clkbuf_2
X_5497_ hold590/X _5520_/B _5496_/Y _5415_/X vssd1 vssd1 vccd1 vccd1 _5497_/X sky130_fd_sc_hd__a22o_1
X_4517_ _4182_/X hold240/X _4518_/S vssd1 vssd1 vccd1 vccd1 _4517_/X sky130_fd_sc_hd__mux2_1
Xhold132 _6239_/Q vssd1 vssd1 vccd1 vccd1 hold132/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold121 _6149_/Q vssd1 vssd1 vccd1 vccd1 hold121/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4479__S _4482_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold165 _6262_/Q vssd1 vssd1 vccd1 vccd1 hold165/X sky130_fd_sc_hd__dlygate4sd3_1
X_4448_ _4445_/X _4446_/X _4447_/X _4441_/S vssd1 vssd1 vccd1 vccd1 _4448_/X sky130_fd_sc_hd__a22o_2
Xhold176 _6191_/Q vssd1 vssd1 vccd1 vccd1 hold176/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold154 _4554_/X vssd1 vssd1 vccd1 vccd1 _6266_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold187 _6183_/Q vssd1 vssd1 vccd1 vccd1 hold187/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4298__A2 _4322_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold198 _4497_/X vssd1 vssd1 vccd1 vccd1 _6206_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4917__S1 _6129_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4379_ hold91/X _3954_/X _4385_/S vssd1 vssd1 vccd1 vccd1 hold92/A sky130_fd_sc_hd__mux2_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6118_ _6489_/CLK _6118_/D vssd1 vssd1 vccd1 vccd1 _6118_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6049_ _6101_/B _4844_/X _5445_/X _6036_/X vssd1 vssd1 vccd1 vccd1 _6049_/X sky130_fd_sc_hd__o22a_1
XANTENNA__3412__A _4313_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3785__C _5317_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5707__C1 _5730_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5486__A1 input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5789__A2 _5771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5948__S _5974_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3750_ _3750_/A _3750_/B vssd1 vssd1 vccd1 vccd1 _3750_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_27_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3681_ _3675_/X _3677_/X _3680_/Y _3669_/Y vssd1 vssd1 vccd1 vccd1 _3681_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5420_ _5414_/Y _5417_/Y _5419_/X _5567_/B vssd1 vssd1 vccd1 vccd1 _5420_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_40_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5351_ _5346_/X _5350_/Y _5341_/X vssd1 vssd1 vccd1 vccd1 _5351_/X sky130_fd_sc_hd__o21a_1
XANTENNA__4299__S _5232_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4921__B1 _4789_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4600__B _4641_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5282_ _5282_/A vssd1 vssd1 vccd1 vccd1 _5282_/Y sky130_fd_sc_hd__inv_2
X_4302_ _4303_/C _4301_/X _4302_/S vssd1 vssd1 vccd1 vccd1 _4302_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_2_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4233_ _6158_/Q _4406_/B _4441_/S vssd1 vssd1 vccd1 vccd1 _4233_/X sky130_fd_sc_hd__or3_1
X_4164_ _6290_/Q _4207_/C vssd1 vssd1 vccd1 vccd1 _4210_/B sky130_fd_sc_hd__xor2_1
X_4095_ _4095_/A _4095_/B vssd1 vssd1 vccd1 vccd1 _4095_/X sky130_fd_sc_hd__or2_1
X_3115_ _3511_/A _3986_/A vssd1 vssd1 vccd1 vccd1 _3115_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__6019__S _6019_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3232__A _4557_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4762__S _4768_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5401__A1 _5315_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4997_ _6403_/Q _4996_/X _5016_/S vssd1 vssd1 vccd1 vccd1 _4997_/X sky130_fd_sc_hd__mux2_1
X_3948_ _4190_/A _3948_/B vssd1 vssd1 vccd1 vccd1 _4045_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_73_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6362__RESET_B fanout181/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3879_ _3878_/B _3878_/C _3892_/A vssd1 vssd1 vccd1 vccd1 _3880_/B sky130_fd_sc_hd__a21o_1
XANTENNA__5593__S _5593_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5618_ _5374_/B _4332_/B _4344_/Y _5617_/Y vssd1 vssd1 vccd1 vccd1 _5618_/X sky130_fd_sc_hd__a211o_1
XANTENNA__5704__A2 _5721_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5549_ hold541/X _5548_/X _5581_/S vssd1 vssd1 vccd1 vccd1 _5549_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6488__SET_B fanout172/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3126__B _4557_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3142__A _3497_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5768__S _5769_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold635_A _6311_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5995__C _5995_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5079__S0 _5100_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3796__B _3883_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout60 _5975_/S vssd1 vssd1 vccd1 vccd1 _6021_/S sky130_fd_sc_hd__buf_8
Xfanout82 _4408_/S vssd1 vssd1 vccd1 vccd1 _5721_/B1 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_91_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3954__B2 _4441_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout93 _5016_/S vssd1 vssd1 vccd1 vccd1 _6070_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_101_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4701__A _6097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5156__A0 _6335_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5008__S _5108_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output52_A _3659_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_26_wb_clk_i _6448_/CLK vssd1 vssd1 vccd1 vccd1 _6475_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_35_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5631__A1 _5644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4920_ _5102_/A _4920_/B vssd1 vssd1 vccd1 vccd1 _4920_/X sky130_fd_sc_hd__and2_1
XFILLER_0_87_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4851_ _6460_/Q _4963_/B _4846_/X _5109_/A1 vssd1 vssd1 vccd1 vccd1 _4852_/C sky130_fd_sc_hd__a22o_1
XFILLER_0_28_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5395__A0 _4406_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3802_ _3865_/S _3818_/C vssd1 vssd1 vccd1 vccd1 _4474_/A sky130_fd_sc_hd__nand2_2
X_4782_ _4782_/A _4782_/B _6300_/Q vssd1 vssd1 vccd1 vccd1 _4782_/X sky130_fd_sc_hd__and3_1
XFILLER_0_27_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3733_ _4546_/A _4519_/A vssd1 vssd1 vccd1 vccd1 _4241_/S sky130_fd_sc_hd__or2_4
X_3664_ _5757_/A _6019_/S _4325_/A vssd1 vssd1 vccd1 vccd1 _6283_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6452_ _6452_/CLK _6452_/D vssd1 vssd1 vccd1 vccd1 _6452_/Q sky130_fd_sc_hd__dfxtp_1
X_5403_ _3386_/A _4363_/B _4362_/Y vssd1 vssd1 vccd1 vccd1 _5403_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_42_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5698__A1 _6462_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3595_ _5387_/C _5619_/A vssd1 vssd1 vccd1 vccd1 _5362_/A sky130_fd_sc_hd__nor2_2
X_6383_ _6383_/CLK _6383_/D vssd1 vssd1 vccd1 vccd1 _6383_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5334_ _5757_/B _5786_/A vssd1 vssd1 vccd1 vccd1 _5368_/S sky130_fd_sc_hd__nor2_2
XANTENNA__5145__C _6021_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5265_ _5322_/A _6339_/Q _4115_/A vssd1 vssd1 vccd1 vccd1 _5265_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__4757__S _5289_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4216_ _4216_/A vssd1 vssd1 vccd1 vccd1 _4216_/Y sky130_fd_sc_hd__inv_2
X_5196_ _6379_/Q _3927_/Y _3987_/B _6380_/Q vssd1 vssd1 vccd1 vccd1 _5196_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_48_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4147_ _4147_/A _4147_/B vssd1 vssd1 vccd1 vccd1 _4149_/A sky130_fd_sc_hd__nor2_1
X_4078_ _4078_/A _4087_/B vssd1 vssd1 vccd1 vccd1 _4078_/X sky130_fd_sc_hd__and2_1
XFILLER_0_92_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6102__A2 _6070_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4113__A1 _6289_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5861__A1 _6367_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3194__D_N _3168_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5613__A1 _5600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3600__A _4653_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4150__B _6384_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3380_ _4344_/A _3338_/X _3375_/X _3379_/X _3334_/B vssd1 vssd1 vccd1 vccd1 _3380_/X
+ sky130_fd_sc_hd__o2111a_1
XANTENNA__4352__A1 _5607_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5050_ _5109_/A1 _5045_/X _5049_/X _4924_/C vssd1 vssd1 vccd1 vccd1 _5050_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4655__A2 _4652_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4001_ _5136_/A _6381_/Q vssd1 vssd1 vccd1 vccd1 _4004_/C sky130_fd_sc_hd__and2_1
XANTENNA__5604__A1 _4595_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4407__A2 _4408_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5952_ _5952_/A _5952_/B vssd1 vssd1 vccd1 vccd1 _5954_/A sky130_fd_sc_hd__nand2_1
XANTENNA__6093__A _6093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4606__A _4641_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_46_wb_clk_i_A clkbuf_leaf_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_4903_ _6418_/Q _6366_/Q _5105_/S vssd1 vssd1 vccd1 vccd1 _4903_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_87_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5883_ _5890_/A _5883_/B vssd1 vssd1 vccd1 vccd1 _5884_/C sky130_fd_sc_hd__or2_1
XFILLER_0_75_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4834_ _4833_/X _6362_/Q _5861_/S vssd1 vssd1 vccd1 vccd1 _4834_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_7_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4765_ hold637/X _4764_/X _5232_/S vssd1 vssd1 vccd1 vccd1 _6315_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_7_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4040__B1 _4463_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4591__A1 _4675_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3656__S input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3716_ _5295_/A _3711_/Y _4948_/S vssd1 vssd1 vccd1 vccd1 _3717_/B sky130_fd_sc_hd__a21o_1
XANTENNA_fanout121_A _5478_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4696_ _6093_/A _4714_/S vssd1 vssd1 vccd1 vccd1 _4696_/Y sky130_fd_sc_hd__nor2_1
X_6435_ _6444_/CLK _6435_/D fanout177/X vssd1 vssd1 vccd1 vccd1 _6435_/Q sky130_fd_sc_hd__dfrtp_4
X_3647_ _3641_/X _3650_/A _3647_/C _3647_/D vssd1 vssd1 vccd1 vccd1 _3647_/X sky130_fd_sc_hd__and4bb_1
XFILLER_0_3_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4343__A1 _5398_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3578_ _3285_/B _5146_/D _3569_/X _3575_/Y _3577_/X vssd1 vssd1 vccd1 vccd1 _3578_/X
+ sky130_fd_sc_hd__o221a_1
X_6366_ _6462_/CLK _6366_/D fanout181/X vssd1 vssd1 vccd1 vccd1 _6366_/Q sky130_fd_sc_hd__dfrtp_4
X_5317_ _5317_/A _5317_/B vssd1 vssd1 vccd1 vccd1 _5317_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__4487__S _4491_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6297_ _6446_/CLK _6297_/D fanout184/X vssd1 vssd1 vccd1 vccd1 _6297_/Q sky130_fd_sc_hd__dfrtp_2
Xhold14 hold14/A vssd1 vssd1 vccd1 vccd1 hold14/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 hold36/A vssd1 vssd1 vccd1 vccd1 hold36/X sky130_fd_sc_hd__dlygate4sd3_1
X_5248_ _6383_/Q _5314_/S _4223_/A _4113_/X _4115_/X vssd1 vssd1 vccd1 vccd1 _5248_/X
+ sky130_fd_sc_hd__a311o_1
Xhold47 hold47/A vssd1 vssd1 vccd1 vccd1 hold47/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 hold25/A vssd1 vssd1 vccd1 vccd1 hold25/X sky130_fd_sc_hd__dlygate4sd3_1
X_5179_ _6334_/Q _4104_/B _4203_/A _5178_/Y vssd1 vssd1 vccd1 vccd1 _5180_/B sky130_fd_sc_hd__o211a_1
Xhold58 hold58/A vssd1 vssd1 vccd1 vccd1 hold58/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold69 hold69/A vssd1 vssd1 vccd1 vccd1 hold69/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5359__B1 _4313_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6020__A1 _4325_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4031__B1 _3795_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3793__C _3884_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4397__S _4397_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6087__A1 _6101_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6087__B2 _6036_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4637__A2 _4611_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3845__B1 _3804_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6465__RESET_B fanout181/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5598__A0 _6465_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xci2406_z80_204 vssd1 vssd1 vccd1 vccd1 ci2406_z80_204/HI io_oeb[19] sky130_fd_sc_hd__conb_1
Xci2406_z80_215 vssd1 vssd1 vccd1 vccd1 io_oeb[30] ci2406_z80_215/LO sky130_fd_sc_hd__conb_1
XANTENNA__4270__B1 _5605_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3612__A3 _3281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4573__A1 _6338_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4550_ _4042_/X hold165/X _4554_/S vssd1 vssd1 vccd1 vccd1 _4550_/X sky130_fd_sc_hd__mux2_1
Xhold506 _6289_/Q vssd1 vssd1 vccd1 vccd1 hold506/X sky130_fd_sc_hd__dlygate4sd3_1
X_3501_ _3501_/A _3501_/B vssd1 vssd1 vccd1 vccd1 _6019_/S sky130_fd_sc_hd__nand2_8
Xhold517 _6029_/X vssd1 vssd1 vccd1 vccd1 _6470_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4481_ hold53/X _4456_/X _4482_/S vssd1 vssd1 vccd1 vccd1 hold54/A sky130_fd_sc_hd__mux2_1
X_3432_ _3399_/X _3411_/Y _4325_/A vssd1 vssd1 vccd1 vccd1 _3432_/X sky130_fd_sc_hd__o21a_1
Xhold528 _4569_/X vssd1 vssd1 vccd1 vccd1 _6276_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6220_ _6263_/CLK _6220_/D vssd1 vssd1 vccd1 vccd1 _6220_/Q sky130_fd_sc_hd__dfxtp_1
Xhold539 _6376_/Q vssd1 vssd1 vccd1 vccd1 hold539/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3363_ _4716_/A _3511_/A _3986_/A vssd1 vssd1 vccd1 vccd1 _5374_/C sky130_fd_sc_hd__and3_1
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6151_ _6399_/CLK _6151_/D vssd1 vssd1 vccd1 vccd1 _6151_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_41_wb_clk_i clkbuf_leaf_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6393_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5102_ _5102_/A _5102_/B vssd1 vssd1 vccd1 vccd1 _5102_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__6078__A1 _4366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3294_ _5315_/A _4273_/B vssd1 vssd1 vccd1 vccd1 _4332_/B sky130_fd_sc_hd__nor2_4
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6082_ _4366_/A _6080_/X _6081_/Y hold520/X _6077_/Y vssd1 vssd1 vccd1 vccd1 _6082_/X
+ sky130_fd_sc_hd__o32a_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5033_ _6372_/Q _5848_/S _5972_/B1 _5032_/X vssd1 vssd1 vccd1 vccd1 _5033_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3836__B1 _3807_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_2_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_5935_ _6421_/Q _6422_/Q _6423_/Q _6424_/Q _5970_/A vssd1 vssd1 vccd1 vccd1 _5935_/Y
+ sky130_fd_sc_hd__o41ai_1
XANTENNA__5684__S0 _5655_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4770__S _4770_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5866_ _5866_/A _6464_/Q _5866_/C vssd1 vssd1 vccd1 vccd1 _5867_/C sky130_fd_sc_hd__or3_1
XFILLER_0_75_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4817_ hold349/X _5098_/S _4815_/X _4816_/X vssd1 vssd1 vccd1 vccd1 _4817_/X sky130_fd_sc_hd__a22o_1
X_5797_ _5796_/X _6362_/Q _5861_/S vssd1 vssd1 vccd1 vccd1 _5797_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_16_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4748_ _6313_/Q _4720_/X wire92/X hold458/X vssd1 vssd1 vccd1 vccd1 _4748_/X sky130_fd_sc_hd__a2bb2o_1
XANTENNA__5761__A0 _6312_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4564__A1 _6313_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4679_ _4713_/A _4678_/X _4714_/S vssd1 vssd1 vccd1 vccd1 _4679_/X sky130_fd_sc_hd__o21a_1
X_6418_ _6422_/CLK _6418_/D fanout173/X vssd1 vssd1 vccd1 vccd1 _6418_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_0_101_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput48 _6301_/Q vssd1 vssd1 vccd1 vccd1 io_out[29] sky130_fd_sc_hd__buf_12
Xoutput37 _6330_/Q vssd1 vssd1 vccd1 vccd1 io_out[19] sky130_fd_sc_hd__buf_12
Xoutput26 _6529_/A vssd1 vssd1 vccd1 vccd1 io_oeb[29] sky130_fd_sc_hd__buf_12
X_6349_ _6377_/CLK _6349_/D fanout176/X vssd1 vssd1 vccd1 vccd1 _6349_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__6069__A1 _6100_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3827__B1 _3852_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5630__A _5644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold548_A _6290_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3150__A _5315_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3763__C1 _6378_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4307__A1 _6312_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4858__A2 _5771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5016__S _5016_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5807__B2 _5977_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3981_ _6285_/Q _6286_/Q vssd1 vssd1 vccd1 vccd1 _3982_/B sky130_fd_sc_hd__xor2_1
XANTENNA__4243__B1 _5322_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5720_ _6224_/Q _5721_/A2 _5721_/B1 _6117_/Q _5730_/C1 vssd1 vssd1 vccd1 vccd1 _5722_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_84_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5991__B1 _3489_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5338__A3 _5387_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5651_ _6421_/Q _5643_/X _5646_/X _5792_/A _5650_/X vssd1 vssd1 vccd1 vccd1 _5651_/X
+ sky130_fd_sc_hd__a221o_1
X_5582_ _6489_/Q _6101_/C _5593_/S vssd1 vssd1 vccd1 vccd1 _5584_/B sky130_fd_sc_hd__mux2_1
X_4602_ _4605_/C _4607_/B vssd1 vssd1 vccd1 vccd1 _4602_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_53_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4533_ hold85/X _4441_/X _4536_/S vssd1 vssd1 vccd1 vccd1 hold86/A sky130_fd_sc_hd__mux2_1
XFILLER_0_25_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold303 _6433_/Q vssd1 vssd1 vccd1 vccd1 _3480_/B sky130_fd_sc_hd__clkbuf_2
Xhold314 _6357_/Q vssd1 vssd1 vccd1 vccd1 _4354_/A sky130_fd_sc_hd__buf_1
Xhold325 _4302_/X vssd1 vssd1 vccd1 vccd1 _6122_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold347 _6160_/Q vssd1 vssd1 vccd1 vccd1 hold347/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold369 _6328_/Q vssd1 vssd1 vccd1 vccd1 hold369/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold336 _6326_/Q vssd1 vssd1 vccd1 vccd1 hold336/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold358 _5859_/X vssd1 vssd1 vccd1 vccd1 _6418_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4464_ hold260/X _4463_/X _4464_/S vssd1 vssd1 vccd1 vccd1 _4464_/X sky130_fd_sc_hd__mux2_1
X_6203_ _6452_/CLK _6203_/D vssd1 vssd1 vccd1 vccd1 _6203_/Q sky130_fd_sc_hd__dfxtp_1
X_3415_ _4784_/D _3412_/Y _3413_/Y _3674_/A vssd1 vssd1 vccd1 vccd1 _3415_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_68_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4395_ hold105/X _4138_/X _4397_/S vssd1 vssd1 vccd1 vccd1 _4395_/X sky130_fd_sc_hd__mux2_1
X_3346_ _4268_/A _3334_/B _3345_/X _3329_/X _3334_/C vssd1 vssd1 vccd1 vccd1 _3346_/X
+ sky130_fd_sc_hd__o2111a_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6134_ _6399_/CLK _6134_/D vssd1 vssd1 vccd1 vccd1 _6134_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4765__S _5232_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6065_ _6101_/B _4920_/B _5496_/Y _6036_/X vssd1 vssd1 vccd1 vccd1 _6065_/X sky130_fd_sc_hd__o22a_1
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3277_ _3699_/A _4324_/B vssd1 vssd1 vccd1 vccd1 _4263_/A sky130_fd_sc_hd__or2_2
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5016_ _6404_/Q _5015_/Y _5016_/S vssd1 vssd1 vccd1 vccd1 _5016_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4234__B1 _5721_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5918_ _5964_/A _5918_/B vssd1 vssd1 vccd1 vccd1 _5918_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_91_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4880__S1 _5100_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5849_ _5817_/A _5848_/X _4901_/Y vssd1 vssd1 vccd1 vccd1 _5849_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_90_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5344__B _5344_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5265__A2 _6339_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3799__B _3818_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4776__A1 _5866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3055__A _3168_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3200_ _4782_/B _3547_/C vssd1 vssd1 vccd1 vccd1 _5360_/B sky130_fd_sc_hd__nand2_1
XANTENNA__4700__A1 _4715_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4180_ hold7/X _4462_/A2 _4463_/S vssd1 vssd1 vccd1 vccd1 _4180_/X sky130_fd_sc_hd__o21a_1
X_3131_ _3205_/B _3332_/A vssd1 vssd1 vccd1 vccd1 _5345_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_38_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3062_ _6159_/Q vssd1 vssd1 vccd1 vccd1 _3062_/Y sky130_fd_sc_hd__inv_2
XANTENNA__6085__B _6107_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4767__B2 _4957_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4767__A1 _6316_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3964_ _4190_/A _3948_/B _3902_/Y vssd1 vssd1 vccd1 vccd1 _3966_/C sky130_fd_sc_hd__o21bai_1
X_5703_ _6338_/Q _5628_/X _5643_/X _6426_/Q vssd1 vssd1 vccd1 vccd1 _5713_/B sky130_fd_sc_hd__a22o_1
XANTENNA__4862__S1 _5078_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3895_ _4430_/B _4425_/A _4425_/B _5300_/C _3858_/Y vssd1 vssd1 vccd1 vccd1 _4437_/B
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_72_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5634_ hold87/A _4406_/B _4420_/S hold65/A _3909_/Y vssd1 vssd1 vccd1 vccd1 _5634_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3727__C1 _4948_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5565_ _5565_/A _5565_/B vssd1 vssd1 vccd1 vccd1 _5565_/Y sky130_fd_sc_hd__xnor2_1
Xhold100 _4498_/X vssd1 vssd1 vccd1 vccd1 _6207_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold144 _6030_/X vssd1 vssd1 vccd1 vccd1 _6471_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold111 _6140_/Q vssd1 vssd1 vccd1 vccd1 hold111/X sky130_fd_sc_hd__dlygate4sd3_1
X_4516_ _4138_/X hold222/X _4518_/S vssd1 vssd1 vccd1 vccd1 _6223_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_13_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold122 _4385_/X vssd1 vssd1 vccd1 vccd1 _6149_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold133 _4534_/X vssd1 vssd1 vccd1 vccd1 _6239_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5496_ _5496_/A _5496_/B vssd1 vssd1 vccd1 vccd1 _5496_/Y sky130_fd_sc_hd__xnor2_1
Xhold166 _4550_/X vssd1 vssd1 vccd1 vccd1 _6262_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold177 _6155_/Q vssd1 vssd1 vccd1 vccd1 hold177/X sky130_fd_sc_hd__dlygate4sd3_1
X_4447_ hold67/X hold176/X hold99/X hold132/X _5721_/C1 _5721_/B1 vssd1 vssd1 vccd1
+ vccd1 _4447_/X sky130_fd_sc_hd__mux4_1
Xhold155 _6452_/Q vssd1 vssd1 vccd1 vccd1 hold155/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold199 _6187_/Q vssd1 vssd1 vccd1 vccd1 hold199/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold188 _4471_/X vssd1 vssd1 vccd1 vccd1 _6183_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6117_ _6239_/CLK _6117_/D vssd1 vssd1 vccd1 vccd1 _6117_/Q sky130_fd_sc_hd__dfxtp_1
X_4378_ hold163/X _3911_/X _4385_/S vssd1 vssd1 vccd1 vccd1 _4378_/X sky130_fd_sc_hd__mux2_1
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4495__S _4500_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3329_ _5774_/C _4325_/C _3557_/B _3329_/D vssd1 vssd1 vccd1 vccd1 _3329_/X sky130_fd_sc_hd__and4b_1
XANTENNA__6150__RESET_B fanout183/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6048_ _5384_/A _6046_/X _6047_/Y hold460/X _6040_/Y vssd1 vssd1 vccd1 vccd1 _6048_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_0_83_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5707__B1 _5721_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4694__B1 _4714_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4446__B1 _4463_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4418__B _6355_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4749__A1 _6313_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4749__B2 _4957_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3680_ _5605_/C _5369_/D vssd1 vssd1 vccd1 vccd1 _3680_/Y sky130_fd_sc_hd__nand2_1
X_5350_ _5350_/A _5350_/B vssd1 vssd1 vccd1 vccd1 _5350_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__4921__A1 _6367_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5281_ _6067_/A _5280_/X _5292_/S vssd1 vssd1 vccd1 vccd1 _5282_/A sky130_fd_sc_hd__mux2_1
X_4301_ _6311_/Q _3091_/Y _4310_/S vssd1 vssd1 vccd1 vccd1 _4301_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_10_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3216__C _5388_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4232_ _6356_/Q _4463_/S vssd1 vssd1 vccd1 vccd1 _5732_/A sky130_fd_sc_hd__nand2_4
X_4163_ _4212_/A _4203_/B _4161_/X vssd1 vssd1 vccd1 vccd1 _4163_/Y sky130_fd_sc_hd__o21ai_1
X_4094_ _4095_/A _4095_/B vssd1 vssd1 vccd1 vccd1 _4094_/Y sky130_fd_sc_hd__nand2_1
X_3114_ _6300_/Q _6299_/Q vssd1 vssd1 vccd1 vccd1 _3326_/B sky130_fd_sc_hd__nand2_8
XFILLER_0_65_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5634__C1 _3909_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout151_A _4675_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4996_ _6459_/Q _4995_/X _5974_/S vssd1 vssd1 vccd1 vccd1 _4996_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_58_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3947_ _3947_/A _3947_/B _3947_/C vssd1 vssd1 vccd1 vccd1 _3948_/B sky130_fd_sc_hd__or3_4
XANTENNA__5874__S _5874_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3878_ _3892_/A _3878_/B _3878_/C vssd1 vssd1 vccd1 vccd1 _3878_/X sky130_fd_sc_hd__and3_1
XFILLER_0_33_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5617_ _5617_/A _5617_/B vssd1 vssd1 vccd1 vccd1 _5617_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_5_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5548_ _6460_/Q _5547_/X _5598_/S vssd1 vssd1 vccd1 vccd1 _5548_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4912__A1 _6366_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5479_ _5492_/A _5479_/B _5479_/C vssd1 vssd1 vccd1 vccd1 _5481_/A sky130_fd_sc_hd__and3_1
XFILLER_0_1_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4140__A2 _3793_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5114__S _5974_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout64_A _5887_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5640__A2 _5732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3651__A1 hold526/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold628_A _6465_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5928__A0 _6461_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5079__S1 _5100_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3796__C _3884_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout61 _3387_/Y vssd1 vssd1 vccd1 vccd1 _5109_/A1 sky130_fd_sc_hd__clkbuf_8
Xfanout83 _4408_/S vssd1 vssd1 vccd1 vccd1 _4235_/S sky130_fd_sc_hd__buf_4
Xfanout72 _5531_/A vssd1 vssd1 vccd1 vccd1 _5594_/A sky130_fd_sc_hd__buf_4
XFILLER_0_36_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout94 _5016_/S vssd1 vssd1 vccd1 vccd1 _4957_/S sky130_fd_sc_hd__clkbuf_8
XANTENNA__4701__B _4714_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4903__A1 _6366_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5024__S _5105_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3333__A _4273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4419__B1 _5731_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4754__A1_N _6314_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4863__S _5101_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5092__A0 _6408_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5631__A2 _5645_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_36_wb_clk_i_A clkbuf_leaf_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__4164__A _6290_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4850_ _4883_/C _4850_/B vssd1 vssd1 vccd1 vccd1 _4852_/B sky130_fd_sc_hd__nor2_1
XANTENNA__5919__B1 _5771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3801_ _3865_/S _3818_/C vssd1 vssd1 vccd1 vccd1 _3801_/X sky130_fd_sc_hd__and2_2
X_4781_ _4557_/C _4784_/B _5774_/B _5372_/B _4335_/C vssd1 vssd1 vccd1 vccd1 _4803_/B
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_43_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3945__A2 _3804_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3732_ _3852_/A _3885_/A _3884_/S vssd1 vssd1 vccd1 vccd1 _4519_/A sky130_fd_sc_hd__or3_1
X_3663_ _3665_/A _5478_/S vssd1 vssd1 vccd1 vccd1 _5295_/B sky130_fd_sc_hd__nand2_1
X_6451_ _6456_/CLK _6451_/D vssd1 vssd1 vccd1 vccd1 _6451_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4611__B _4611_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5402_ _4595_/B _3527_/X _5400_/X hold346/X vssd1 vssd1 vccd1 vccd1 _6359_/D sky130_fd_sc_hd__a22o_1
X_6382_ _6384_/CLK _6382_/D vssd1 vssd1 vccd1 vccd1 _6382_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_42_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5333_ _5757_/B hold230/X _5331_/X _5332_/X vssd1 vssd1 vccd1 vccd1 _5333_/X sky130_fd_sc_hd__a22o_1
X_3594_ _3594_/A _3594_/B vssd1 vssd1 vccd1 vccd1 _3602_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5264_ _5264_/A _5264_/B _5264_/C vssd1 vssd1 vccd1 vccd1 _5264_/X sky130_fd_sc_hd__or3_1
XFILLER_0_76_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5195_ _5195_/A _5195_/B vssd1 vssd1 vccd1 vccd1 _5195_/Y sky130_fd_sc_hd__xnor2_1
X_4215_ _6291_/Q _3770_/A _3773_/Y _5171_/B vssd1 vssd1 vccd1 vccd1 _4216_/A sky130_fd_sc_hd__a22oi_1
X_4146_ _4190_/A _4146_/B vssd1 vssd1 vccd1 vccd1 _4147_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_78_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4077_ _6462_/Q _4076_/X _6347_/Q vssd1 vssd1 vccd1 vccd1 _4077_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_78_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4979_ _6152_/Q hold91/A _6135_/Q _6179_/Q _5100_/S0 _5100_/S1 vssd1 vssd1 vccd1
+ vccd1 _4979_/X sky130_fd_sc_hd__mux4_1
XANTENNA__5617__B _5617_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6279__SET_B fanout183/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3107__A_N _3168_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4948__S _4948_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4683__S _4712_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5613__A2 _5388_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5377__A1 _5364_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5808__A _5866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4337__C1 _5388_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4000_ _5136_/A _6381_/Q vssd1 vssd1 vccd1 vccd1 _4004_/B sky130_fd_sc_hd__nor2_1
XANTENNA__3063__A _4324_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3213__D _4595_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5065__B1 _4963_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5951_ _5951_/A _5970_/A vssd1 vssd1 vccd1 vccd1 _5952_/B sky130_fd_sc_hd__or2_1
XANTENNA__6093__B _6107_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4902_ _6366_/Q _4790_/X _4789_/B vssd1 vssd1 vccd1 vccd1 _4902_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_62_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5882_ _6420_/Q _5970_/A vssd1 vssd1 vccd1 vccd1 _5883_/B sky130_fd_sc_hd__nor2_1
X_4833_ _5892_/S _4832_/X _4818_/X vssd1 vssd1 vccd1 vccd1 _4833_/X sky130_fd_sc_hd__a21o_1
X_4764_ _4177_/Y _4763_/X _4770_/S vssd1 vssd1 vccd1 vccd1 _4764_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_43_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3715_ _5295_/A _3711_/Y _4948_/S vssd1 vssd1 vccd1 vccd1 _3715_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_0_7_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4695_ _4715_/B2 _4691_/Y _4694_/X hold316/X _4672_/Y vssd1 vssd1 vccd1 vccd1 _4695_/X
+ sky130_fd_sc_hd__o32a_1
X_6434_ _6439_/CLK _6434_/D fanout178/X vssd1 vssd1 vccd1 vccd1 _6434_/Q sky130_fd_sc_hd__dfrtp_4
X_3646_ _6468_/Q _3645_/Y _3640_/A vssd1 vssd1 vccd1 vccd1 _3646_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_3_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout114_A _6108_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4343__A2 _5362_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3577_ _5387_/B _4325_/C _4386_/B _4675_/C _5607_/B2 vssd1 vssd1 vccd1 vccd1 _3577_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_60_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6365_ _6475_/CLK _6365_/D fanout181/X vssd1 vssd1 vccd1 vccd1 _6365_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__4768__S _4768_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5540__A1 _5002_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5453__A _5492_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6296_ _6446_/CLK _6296_/D fanout184/X vssd1 vssd1 vccd1 vccd1 _6296_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__3551__B1 _3525_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5316_ _5364_/A _5316_/B vssd1 vssd1 vccd1 vccd1 _5316_/Y sky130_fd_sc_hd__nor2_1
X_5247_ _6383_/Q _5257_/B _5247_/S vssd1 vssd1 vccd1 vccd1 _5247_/X sky130_fd_sc_hd__mux2_1
Xhold37 hold37/A vssd1 vssd1 vccd1 vccd1 hold37/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 hold26/A vssd1 vssd1 vccd1 vccd1 hold26/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold15 hold15/A vssd1 vssd1 vccd1 vccd1 hold15/X sky130_fd_sc_hd__dlygate4sd3_1
X_5178_ _6334_/Q _5178_/B vssd1 vssd1 vccd1 vccd1 _5178_/Y sky130_fd_sc_hd__nand2_1
Xhold59 hold59/A vssd1 vssd1 vccd1 vccd1 hold59/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold48 hold48/A vssd1 vssd1 vccd1 vccd1 hold48/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5599__S _6104_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4129_ _4190_/A _4131_/B vssd1 vssd1 vccd1 vccd1 _4130_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_97_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3701__A _4418_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3909__A2 _4418_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5628__A _5644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4678__S _4712_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4334__A2 _3632_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6087__A2 _5021_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xci2406_z80_205 vssd1 vssd1 vccd1 vccd1 ci2406_z80_205/HI io_oeb[20] sky130_fd_sc_hd__conb_1
Xci2406_z80_216 vssd1 vssd1 vccd1 vccd1 io_oeb[31] ci2406_z80_216/LO sky130_fd_sc_hd__conb_1
XFILLER_0_16_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3500_ _3500_/A _3501_/B vssd1 vssd1 vccd1 vccd1 _5418_/A sky130_fd_sc_hd__and2_4
Xhold507 _4635_/X vssd1 vssd1 vccd1 vccd1 _6289_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4480_ hold176/X _4448_/X _4482_/S vssd1 vssd1 vccd1 vccd1 _6191_/D sky130_fd_sc_hd__mux2_1
Xhold518 _6420_/Q vssd1 vssd1 vccd1 vccd1 hold518/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold529 _6286_/Q vssd1 vssd1 vccd1 vccd1 hold529/X sky130_fd_sc_hd__dlygate4sd3_1
X_3431_ _5980_/A _3431_/B _3431_/C vssd1 vssd1 vccd1 vccd1 _3464_/B sky130_fd_sc_hd__and3_1
X_3362_ _3219_/B _3511_/B _4116_/A _6335_/Q _3361_/Y vssd1 vssd1 vccd1 vccd1 _3370_/A
+ sky130_fd_sc_hd__a221oi_2
X_6150_ _6340_/CLK _6150_/D fanout183/X vssd1 vssd1 vccd1 vccd1 _6150_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3505__B _5769_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5101_ _5100_/X _5099_/X _5101_/S vssd1 vssd1 vccd1 vccd1 _5102_/B sky130_fd_sc_hd__mux2_2
X_3293_ _3288_/X _3291_/X _3292_/X _4263_/A vssd1 vssd1 vccd1 vccd1 _3336_/B sky130_fd_sc_hd__a31o_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6081_ _6081_/A _6107_/S vssd1 vssd1 vccd1 vccd1 _6081_/Y sky130_fd_sc_hd__nor2_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5032_ _6405_/Q _5031_/X _5971_/S vssd1 vssd1 vccd1 vccd1 _5032_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_10_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6472_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_95_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5934_ _5934_/A _5934_/B vssd1 vssd1 vccd1 vccd1 _5937_/A sky130_fd_sc_hd__nand2_1
XANTENNA__5684__S1 _5734_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5865_ hold524/X _6023_/A _5864_/X vssd1 vssd1 vccd1 vccd1 _5865_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_75_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4816_ _4303_/A _6070_/A _5098_/S vssd1 vssd1 vccd1 vccd1 _4816_/X sky130_fd_sc_hd__o21ba_1
XANTENNA__4013__A1 _6285_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5796_ hold474/X _5892_/S _4818_/X vssd1 vssd1 vccd1 vccd1 _5796_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_7_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4747_ hold642/X _4746_/X _5232_/S vssd1 vssd1 vccd1 vccd1 _6312_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4678_ _6382_/Q _4677_/X _4712_/S vssd1 vssd1 vccd1 vccd1 _4678_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_98_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3629_ _4325_/A _3629_/B vssd1 vssd1 vccd1 vccd1 _3629_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__4316__A2 _4310_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4498__S _4500_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6417_ _6417_/CLK _6417_/D fanout173/X vssd1 vssd1 vccd1 vccd1 _6417_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_0_101_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6348_ _6441_/CLK hold44/X fanout185/X vssd1 vssd1 vccd1 vccd1 hold43/A sky130_fd_sc_hd__dfrtp_1
Xoutput49 _3656_/X vssd1 vssd1 vccd1 vccd1 io_out[2] sky130_fd_sc_hd__buf_12
XFILLER_0_3_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput38 _6457_/Q vssd1 vssd1 vccd1 vccd1 io_out[1] sky130_fd_sc_hd__buf_12
Xoutput27 _5581_/S vssd1 vssd1 vccd1 vccd1 io_out[0] sky130_fd_sc_hd__buf_12
XANTENNA__6069__A2 _4949_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6279_ _6312_/CLK _6279_/D fanout183/X vssd1 vssd1 vccd1 vccd1 _6279_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA__3827__A1 _3885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5029__A0 _6461_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5630__B _5645_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4246__B _5757_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4961__S _5101_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold610_A _6337_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5752__A1 _4036_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4307__A2 _4322_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5821__A _5866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5807__A2 _5785_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3980_ _6334_/Q _3079_/Y _4107_/B vssd1 vssd1 vccd1 vccd1 _3982_/A sky130_fd_sc_hd__mux2_1
XANTENNA__4243__A1 _5388_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xmax_cap91 wire92/X vssd1 vssd1 vccd1 vccd1 _5224_/A2 sky130_fd_sc_hd__clkbuf_2
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5268__A _5268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5650_ _6458_/Q _5645_/X _5647_/X _5653_/A _5649_/X vssd1 vssd1 vccd1 vccd1 _5650_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_5_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4601_ _5767_/A _4605_/B vssd1 vssd1 vccd1 vccd1 _4607_/B sky130_fd_sc_hd__nor2_1
X_5581_ hold562/X _5580_/X _5581_/S vssd1 vssd1 vccd1 vccd1 _5581_/X sky130_fd_sc_hd__mux2_1
X_4532_ hold151/X _4435_/X _4536_/S vssd1 vssd1 vccd1 vccd1 _4532_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_4_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold326 _6303_/Q vssd1 vssd1 vccd1 vccd1 hold326/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold304 _3569_/B vssd1 vssd1 vccd1 vccd1 _3488_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold315 _5397_/Y vssd1 vssd1 vccd1 vccd1 hold315/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4463_ _4458_/X _4462_/X _4463_/S vssd1 vssd1 vccd1 vccd1 _4463_/X sky130_fd_sc_hd__mux2_2
X_3414_ _5387_/A _3414_/B vssd1 vssd1 vccd1 vccd1 _5619_/A sky130_fd_sc_hd__or2_2
XFILLER_0_68_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold348 _3528_/X vssd1 vssd1 vccd1 vccd1 _6160_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6202_ _6449_/CLK hold76/X vssd1 vssd1 vccd1 vccd1 hold75/A sky130_fd_sc_hd__dfxtp_1
Xhold359 _6406_/Q vssd1 vssd1 vccd1 vccd1 hold359/X sky130_fd_sc_hd__buf_1
Xhold337 _4998_/X vssd1 vssd1 vccd1 vccd1 _6326_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4394_ hold177/X _4085_/X _4397_/S vssd1 vssd1 vccd1 vccd1 _4394_/X sky130_fd_sc_hd__mux2_1
X_6133_ _6242_/CLK _6133_/D fanout180/X vssd1 vssd1 vccd1 vccd1 _6133_/Q sky130_fd_sc_hd__dfrtp_1
X_3345_ _3304_/B _3344_/X _3342_/X _3317_/X vssd1 vssd1 vccd1 vccd1 _3345_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_68_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3276_ _3699_/A _4324_/B vssd1 vssd1 vccd1 vccd1 _3276_/Y sky130_fd_sc_hd__nor2_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6064_ _4366_/A _6062_/X _6063_/Y hold498/X _6040_/Y vssd1 vssd1 vccd1 vccd1 _6064_/X
+ sky130_fd_sc_hd__o32a_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5015_ _5771_/A _5013_/X _5014_/Y vssd1 vssd1 vccd1 vccd1 _5015_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_84_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout181_A fanout185/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5917_ _6371_/Q _5848_/S _5972_/B1 _5916_/X vssd1 vssd1 vccd1 vccd1 _5918_/B sky130_fd_sc_hd__a22o_1
XANTENNA__5178__A _6334_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5848_ _5847_/X _6366_/Q _5848_/S vssd1 vssd1 vccd1 vccd1 _5848_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_90_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5779_ _5866_/A _5866_/C hold43/A vssd1 vssd1 vccd1 vccd1 _5867_/B sky130_fd_sc_hd__o21bai_4
XFILLER_0_8_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout94_A _5016_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3145__B _3168_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4956__S _5974_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold560_A _6426_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3984__A0 _6285_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4776__A2 _4774_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5725__A1 _6315_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4720__A _5866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4084__S0 _5721_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3130_ _3639_/C _3163_/A vssd1 vssd1 vccd1 vccd1 _3332_/A sky130_fd_sc_hd__or2_1
XANTENNA__3071__A hold1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3061_ _3665_/A vssd1 vssd1 vccd1 vccd1 _4325_/A sky130_fd_sc_hd__inv_6
XFILLER_0_89_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3963_ _3814_/Y _3948_/B _4190_/A vssd1 vssd1 vccd1 vccd1 _3966_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_70_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5702_ _6480_/Q _5629_/X _5646_/X _5852_/A vssd1 vssd1 vccd1 vccd1 _5713_/A sky130_fd_sc_hd__a22o_1
X_3894_ _5300_/C _3894_/B vssd1 vssd1 vccd1 vccd1 _4431_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_45_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5633_ _6226_/Q _4406_/B _4420_/S _6449_/Q _5731_/C1 vssd1 vssd1 vccd1 vccd1 _5633_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5716__A1 _6339_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5564_ _5545_/A _5544_/Y _5553_/A _5563_/Y vssd1 vssd1 vccd1 vccd1 _5565_/B sky130_fd_sc_hd__o31a_1
XFILLER_0_13_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold101 _6138_/Q vssd1 vssd1 vccd1 vccd1 hold101/X sky130_fd_sc_hd__dlygate4sd3_1
X_4515_ _4085_/X hold297/X _4518_/S vssd1 vssd1 vccd1 vccd1 _6222_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_13_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3246__A _5605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold123 _6205_/Q vssd1 vssd1 vccd1 vccd1 hold123/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold112 _4375_/X vssd1 vssd1 vccd1 vccd1 _6140_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold134 _6139_/Q vssd1 vssd1 vccd1 vccd1 hold134/X sky130_fd_sc_hd__dlygate4sd3_1
X_5495_ _5483_/A _5483_/B _5481_/A vssd1 vssd1 vccd1 vccd1 _5496_/B sky130_fd_sc_hd__a21oi_1
X_4446_ hold27/X _4462_/A2 _4463_/S vssd1 vssd1 vccd1 vccd1 _4446_/X sky130_fd_sc_hd__o21a_1
Xhold145 _6185_/Q vssd1 vssd1 vccd1 vccd1 hold145/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold167 _6201_/Q vssd1 vssd1 vccd1 vccd1 hold167/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold156 _6007_/X vssd1 vssd1 vccd1 vccd1 _6452_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold178 _4394_/X vssd1 vssd1 vccd1 vccd1 _6155_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4377_ _4546_/A _4474_/A vssd1 vssd1 vccd1 vccd1 _4385_/S sky130_fd_sc_hd__nor2_4
Xhold189 _6188_/Q vssd1 vssd1 vccd1 vccd1 hold189/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_95_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3328_ _4344_/A _5617_/A vssd1 vssd1 vccd1 vccd1 _5774_/C sky130_fd_sc_hd__nand2_1
X_6116_ _6223_/CLK _6116_/D vssd1 vssd1 vccd1 vccd1 _6116_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3259_ _4557_/C _3376_/B _3232_/C vssd1 vssd1 vccd1 vccd1 _3261_/B sky130_fd_sc_hd__or3b_1
X_6047_ _6081_/A _6071_/S vssd1 vssd1 vccd1 vccd1 _6047_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_95_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5404__A0 _5404_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5955__A1 _5786_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5955__B2 _5976_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3855__S _3883_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4686__S _4711_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4143__B1 _3810_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4694__A1 _4713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4418__C _4418_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_26_wb_clk_i_A _6448_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3957__B1 _3801_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3066__A _5593_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4921__A2 _4790_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5280_ _5279_/X _5277_/X _5291_/S vssd1 vssd1 vccd1 vccd1 _5280_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_50_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4300_ _4300_/A _4300_/B vssd1 vssd1 vccd1 vccd1 _4302_/S sky130_fd_sc_hd__nor2_1
XFILLER_0_49_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4231_ _6356_/Q _4463_/S vssd1 vssd1 vccd1 vccd1 _5655_/B sky130_fd_sc_hd__and2_4
XANTENNA__4685__A1 _4715_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4162_ _4162_/A _4162_/B vssd1 vssd1 vccd1 vccd1 _4203_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_4_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4093_ _4064_/X _4065_/X _4068_/B vssd1 vssd1 vccd1 vccd1 _4095_/B sky130_fd_sc_hd__a21bo_1
X_3113_ _6300_/Q _6299_/Q vssd1 vssd1 vccd1 vccd1 _4248_/B sky130_fd_sc_hd__and2_1
XFILLER_0_4_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5220__S _5489_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4995_ _5964_/A _4994_/X _4982_/Y vssd1 vssd1 vccd1 vccd1 _4995_/X sky130_fd_sc_hd__a21bo_1
XANTENNA_fanout144_A _4273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3946_ _6112_/Q _3731_/X _3810_/X _6179_/Q _3945_/X vssd1 vssd1 vccd1 vccd1 _3947_/C
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3563__A1_N _6431_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3877_ _3878_/B _3878_/C vssd1 vssd1 vccd1 vccd1 _4611_/A sky130_fd_sc_hd__nand2_1
XANTENNA__4360__A _5600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5616_ _3575_/Y _4583_/X _5614_/Y _5615_/Y vssd1 vssd1 vccd1 vccd1 _5616_/X sky130_fd_sc_hd__o31a_1
XFILLER_0_60_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5547_ hold541/X _5546_/X _6070_/A vssd1 vssd1 vccd1 vccd1 _5547_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5478_ _6480_/Q _4901_/B _5478_/S vssd1 vssd1 vccd1 vccd1 _5479_/C sky130_fd_sc_hd__mux2_1
XANTENNA__4125__B1 _3801_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4429_ hold125/X _4428_/X _4464_/S vssd1 vssd1 vccd1 vccd1 _6172_/D sky130_fd_sc_hd__mux2_1
XANTENNA__6371__RESET_B fanout172/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4428__A1 _4441_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3651__A2 hold1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3939__A0 _5427_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout73 _3909_/Y vssd1 vssd1 vccd1 vccd1 _5730_/C1 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_91_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout95 _3496_/X vssd1 vssd1 vccd1 vccd1 _5016_/S sky130_fd_sc_hd__buf_4
Xfanout84 _4408_/S vssd1 vssd1 vccd1 vccd1 _4420_/S sky130_fd_sc_hd__buf_4
XFILLER_0_101_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6105__A1 _6101_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6459__RESET_B fanout181/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6105__B2 _6036_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4736__A2_N _4720_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output38_A _6457_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5040__S _5101_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4780_ _5817_/A _5413_/B _5974_/S vssd1 vssd1 vccd1 vccd1 _4780_/X sky130_fd_sc_hd__o21a_1
XANTENNA__5975__S _5975_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3800_ _3884_/S _3818_/C vssd1 vssd1 vccd1 vccd1 _4528_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_27_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3731_ _3816_/B _3883_/S _3865_/S vssd1 vssd1 vccd1 vccd1 _3731_/X sky130_fd_sc_hd__and3_4
XFILLER_0_55_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_35_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6428_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_27_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3662_ _3098_/Y _3660_/X _3661_/Y _6165_/Q vssd1 vssd1 vccd1 vccd1 _3662_/X sky130_fd_sc_hd__a22o_2
XFILLER_0_42_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6450_ _6452_/CLK _6450_/D vssd1 vssd1 vccd1 vccd1 _6450_/Q sky130_fd_sc_hd__dfxtp_1
X_3593_ _5980_/A _3530_/A _3592_/X _3699_/A vssd1 vssd1 vccd1 vccd1 _3593_/X sky130_fd_sc_hd__o22a_1
X_5401_ _5315_/A _3527_/X _5400_/X _3390_/B vssd1 vssd1 vccd1 vccd1 _5401_/X sky130_fd_sc_hd__a22o_1
X_6381_ _6383_/CLK _6381_/D vssd1 vssd1 vccd1 vccd1 _6381_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_42_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5332_ _5757_/B _5320_/X _6431_/Q _6160_/Q vssd1 vssd1 vccd1 vccd1 _5332_/X sky130_fd_sc_hd__and4bb_1
XFILLER_0_11_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5263_ _5263_/A _5263_/B _5263_/C vssd1 vssd1 vccd1 vccd1 _5264_/C sky130_fd_sc_hd__or3_1
X_5194_ _5194_/A _5194_/B vssd1 vssd1 vccd1 vccd1 _5195_/B sky130_fd_sc_hd__xnor2_1
X_4214_ _4206_/Y _4213_/X _6334_/Q vssd1 vssd1 vccd1 vccd1 _5171_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_76_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3243__B _3304_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4145_ _4190_/A _4146_/B vssd1 vssd1 vccd1 vccd1 _4147_/A sky130_fd_sc_hd__and2_1
XFILLER_0_92_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4076_ _3738_/X _5257_/A _4075_/X _4057_/Y vssd1 vssd1 vccd1 vccd1 _4076_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_92_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3397__A1 _5398_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4978_ _4977_/X hold415/X _5098_/S vssd1 vssd1 vccd1 vccd1 _4978_/X sky130_fd_sc_hd__mux2_1
X_3929_ _3986_/A _4720_/C _4223_/A _6379_/Q vssd1 vssd1 vccd1 vccd1 _3929_/X sky130_fd_sc_hd__o31a_1
XFILLER_0_80_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3434__A _3632_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5846__B1 _5784_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5377__A2 _5607_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3388__A1 _3530_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5808__B _6460_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4888__B2 _4881_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5035__S _5974_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5950_ _6426_/Q _5970_/A vssd1 vssd1 vccd1 vccd1 _5950_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__5065__B2 _6314_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4901_ _5102_/A _4901_/B vssd1 vssd1 vccd1 vccd1 _4901_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__6014__A0 _4658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5881_ _6420_/Q _5970_/A vssd1 vssd1 vccd1 vccd1 _5890_/A sky130_fd_sc_hd__and2_1
X_4832_ _6414_/Q _4793_/Y _4825_/X _4831_/X vssd1 vssd1 vccd1 vccd1 _4832_/X sky130_fd_sc_hd__a211o_1
XANTENNA__4576__B1 _5364_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4763_ _4761_/X _4762_/X _5289_/S vssd1 vssd1 vccd1 vccd1 _4763_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4040__A2 _4462_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4114__S _4716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4694_ _4713_/A _4693_/X _4714_/S vssd1 vssd1 vccd1 vccd1 _4694_/X sky130_fd_sc_hd__o21a_1
X_3714_ _6359_/Q hold5/A _3714_/S vssd1 vssd1 vccd1 vccd1 _3714_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_43_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6433_ _6444_/CLK _6433_/D fanout178/X vssd1 vssd1 vccd1 vccd1 _6433_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3645_ _3373_/B _3640_/C _3644_/C vssd1 vssd1 vccd1 vccd1 _3645_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_3_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3576_ _3587_/B _5777_/B vssd1 vssd1 vccd1 vccd1 _4675_/C sky130_fd_sc_hd__or2_1
X_6364_ _6475_/CLK _6364_/D fanout181/X vssd1 vssd1 vccd1 vccd1 _6364_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_3_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6295_ _6446_/CLK _6295_/D fanout184/X vssd1 vssd1 vccd1 vccd1 _6295_/Q sky130_fd_sc_hd__dfrtp_1
X_5315_ _5315_/A _5315_/B vssd1 vssd1 vccd1 vccd1 _5315_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__5828__A0 _6364_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5246_ _6338_/Q _5131_/Y _5245_/X _4957_/S _5151_/B vssd1 vssd1 vccd1 vccd1 _5246_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_53_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold38 hold38/A vssd1 vssd1 vccd1 vccd1 hold38/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold27 hold27/A vssd1 vssd1 vccd1 vccd1 hold27/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold16 hold16/A vssd1 vssd1 vccd1 vccd1 hold16/X sky130_fd_sc_hd__dlygate4sd3_1
X_5177_ _5177_/A _5177_/B vssd1 vssd1 vccd1 vccd1 _5180_/A sky130_fd_sc_hd__xnor2_1
Xhold49 hold49/A vssd1 vssd1 vccd1 vccd1 hold49/X sky130_fd_sc_hd__dlygate4sd3_1
X_4128_ _4128_/A _4128_/B vssd1 vssd1 vccd1 vccd1 _4131_/B sky130_fd_sc_hd__or2_2
X_4059_ _4199_/A _6382_/Q vssd1 vssd1 vccd1 vccd1 _4063_/B sky130_fd_sc_hd__nor2_1
XANTENNA__3701__B _3701_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3429__A _4324_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4031__A2 _3793_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3790__A1 _4675_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5644__A _5644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold590_A _6367_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3542__A1 _5384_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3845__A2 _3731_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xci2406_z80_206 vssd1 vssd1 vccd1 vccd1 ci2406_z80_206/HI io_oeb[21] sky130_fd_sc_hd__conb_1
Xci2406_z80_217 vssd1 vssd1 vccd1 vccd1 io_oeb[35] ci2406_z80_217/LO sky130_fd_sc_hd__conb_1
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4723__A _5124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6474__RESET_B fanout180/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold508 _6382_/Q vssd1 vssd1 vccd1 vccd1 _4078_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4869__S _4948_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3430_ _3424_/X _3425_/Y _3417_/X vssd1 vssd1 vccd1 vccd1 _3431_/C sky130_fd_sc_hd__a21oi_1
XFILLER_0_52_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold519 _5888_/X vssd1 vssd1 vccd1 vccd1 _6420_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3361_ _4217_/A _3511_/A _6335_/Q _3986_/A vssd1 vssd1 vccd1 vccd1 _3361_/Y sky130_fd_sc_hd__nor4b_1
XANTENNA__3074__A _6436_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3505__C _5418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5100_ _6266_/Q _6201_/Q _6225_/Q _6118_/Q _5100_/S0 _5100_/S1 vssd1 vssd1 vccd1
+ vccd1 _5100_/X sky130_fd_sc_hd__mux4_1
X_6080_ _6101_/A _6079_/X _6107_/S vssd1 vssd1 vccd1 vccd1 _6080_/X sky130_fd_sc_hd__o21a_1
X_3292_ _4338_/A _4386_/A _3668_/A _5146_/B _5405_/A vssd1 vssd1 vccd1 vccd1 _3292_/X
+ sky130_fd_sc_hd__o221a_1
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5031_ _6424_/Q _4793_/Y _5023_/X _5030_/X vssd1 vssd1 vccd1 vccd1 _5031_/X sky130_fd_sc_hd__a211o_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3836__A2 _3804_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5933_ _5933_/A _5970_/A vssd1 vssd1 vccd1 vccd1 _5934_/B sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_50_wb_clk_i clkbuf_leaf_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6454_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_5864_ _6021_/S _5863_/X _5887_/S vssd1 vssd1 vccd1 vccd1 _5864_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_75_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4815_ _6361_/Q _5771_/A _4780_/X _4814_/X _5783_/A vssd1 vssd1 vccd1 vccd1 _4815_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4013__A2 _6286_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5795_ _5977_/S _5794_/X _5784_/X _5792_/A vssd1 vssd1 vccd1 vccd1 _5795_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_28_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4746_ _4029_/Y _4745_/X _4770_/S vssd1 vssd1 vccd1 vccd1 _4746_/X sky130_fd_sc_hd__mux2_1
X_4677_ _6378_/Q _6284_/Q _4711_/S vssd1 vssd1 vccd1 vccd1 _4677_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_71_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4779__S _4919_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5464__A _5757_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3628_ hold59/A _6132_/Q _6133_/Q _6130_/Q vssd1 vssd1 vccd1 vccd1 _3629_/B sky130_fd_sc_hd__or4_1
XFILLER_0_3_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6416_ _6417_/CLK _6416_/D fanout173/X vssd1 vssd1 vccd1 vccd1 _6416_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_0_101_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6347_ _6441_/CLK _6347_/D fanout184/X vssd1 vssd1 vccd1 vccd1 _6347_/Q sky130_fd_sc_hd__dfrtp_4
Xoutput39 _6331_/Q vssd1 vssd1 vccd1 vccd1 io_out[20] sky130_fd_sc_hd__buf_12
XANTENNA__4721__B1 _4720_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput28 _6318_/Q vssd1 vssd1 vccd1 vccd1 io_out[10] sky130_fd_sc_hd__buf_12
XFILLER_0_101_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3559_ _3411_/A _3674_/B _5387_/C vssd1 vssd1 vccd1 vccd1 _3559_/X sky130_fd_sc_hd__a21o_1
X_6278_ _6312_/CLK _6278_/D fanout182/X vssd1 vssd1 vccd1 vccd1 _6278_/Q sky130_fd_sc_hd__dfstp_1
X_5229_ _3774_/A _5226_/X _5228_/X _4023_/X vssd1 vssd1 vccd1 vccd1 _5229_/X sky130_fd_sc_hd__a211o_1
XANTENNA__4808__A _5108_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4019__S _4716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3150__C _3281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4237__C1 _5730_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5639__A _5655_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_hold603_A _6336_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4712__A0 _6287_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3515__A1 _4332_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5060__S0 _5100_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5821__B _6461_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5440__A1 _4844_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3451__B1 _5995_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4600_ _4600_/A _4641_/B vssd1 vssd1 vccd1 vccd1 _4600_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_38_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5580_ _6463_/Q _5579_/X _5598_/S vssd1 vssd1 vccd1 vccd1 _5580_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_13_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4531_ hold69/X _4428_/X _4536_/S vssd1 vssd1 vccd1 vccd1 hold70/A sky130_fd_sc_hd__mux2_1
XFILLER_0_40_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold305 _3489_/C vssd1 vssd1 vccd1 vccd1 hold305/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold316 _6304_/Q vssd1 vssd1 vccd1 vccd1 hold316/X sky130_fd_sc_hd__dlygate4sd3_1
X_4462_ hold13/X _4462_/A2 _4461_/X vssd1 vssd1 vccd1 vccd1 _4462_/X sky130_fd_sc_hd__o21a_1
X_3413_ _5387_/A _3414_/B vssd1 vssd1 vccd1 vccd1 _3413_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__4703__A0 _6285_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold327 _4690_/X vssd1 vssd1 vccd1 vccd1 _6303_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold338 _6120_/Q vssd1 vssd1 vccd1 vccd1 _4303_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6201_ _6489_/CLK _6201_/D vssd1 vssd1 vccd1 vccd1 _6201_/Q sky130_fd_sc_hd__dfxtp_1
Xhold349 _6317_/Q vssd1 vssd1 vccd1 vccd1 hold349/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4393_ hold73/X _4042_/X _4397_/S vssd1 vssd1 vccd1 vccd1 hold74/A sky130_fd_sc_hd__mux2_1
X_3344_ _3180_/B _3338_/X _3343_/X _3627_/C vssd1 vssd1 vccd1 vccd1 _3344_/X sky130_fd_sc_hd__o211a_1
X_6132_ _6444_/CLK _6132_/D fanout177/X vssd1 vssd1 vccd1 vccd1 _6132_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3275_ _5315_/B _3274_/X _3122_/Y vssd1 vssd1 vccd1 vccd1 _3336_/A sky130_fd_sc_hd__o21a_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6063_ _6097_/A _6071_/S vssd1 vssd1 vccd1 vccd1 _6063_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_84_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5014_ _6460_/Q _5771_/A vssd1 vssd1 vccd1 vccd1 _5014_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_84_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3690__B1 _5317_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout174_A fanout175/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4234__A2 _5721_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4363__A _4363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5916_ _6404_/Q _6423_/Q _5971_/S vssd1 vssd1 vccd1 vccd1 _5916_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_75_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5847_ _6418_/Q _5971_/S _4902_/X vssd1 vssd1 vccd1 vccd1 _5847_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_33_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5778_ _5776_/X _5777_/X _5322_/A vssd1 vssd1 vccd1 vccd1 _5778_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_44_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4729_ hold632/X _4728_/X _5232_/S vssd1 vssd1 vccd1 vccd1 _4729_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4810__B _5108_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5498__A1 input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4170__A1 _6290_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5360__C _5360_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3442__A _3489_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_16_wb_clk_i_A _6448_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4273__A _4273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3984__A1 _6287_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6110__3 _6470_/CLK vssd1 vssd1 vccd1 vccd1 _6167_/CLK sky130_fd_sc_hd__inv_2
X_3060_ _4335_/B vssd1 vssd1 vccd1 vccd1 _5145_/A sky130_fd_sc_hd__inv_4
XFILLER_0_89_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5279__A _6459_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5701_ _4300_/A _4078_/A _5611_/Y _5700_/X vssd1 vssd1 vccd1 vccd1 _5701_/X sky130_fd_sc_hd__a22o_1
X_3962_ _4190_/A _3962_/B vssd1 vssd1 vccd1 vccd1 _4045_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_70_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3893_ _4425_/A _4425_/B vssd1 vssd1 vccd1 vccd1 _3894_/B sky130_fd_sc_hd__or2_1
XANTENNA__6477__SET_B fanout176/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5632_ _5632_/A vssd1 vssd1 vccd1 vccd1 _5632_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_72_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5563_ _5542_/B _5551_/B _5594_/A vssd1 vssd1 vccd1 vccd1 _5563_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_26_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4514_ _4042_/X hold194/X _4518_/S vssd1 vssd1 vccd1 vccd1 _6221_/D sky130_fd_sc_hd__mux2_1
XANTENNA__3246__B _4268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold124 _4496_/X vssd1 vssd1 vccd1 vccd1 _6205_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold135 _4374_/X vssd1 vssd1 vccd1 vccd1 _6139_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold102 _4373_/X vssd1 vssd1 vccd1 vccd1 _6138_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold113 _6208_/Q vssd1 vssd1 vccd1 vccd1 hold113/X sky130_fd_sc_hd__dlygate4sd3_1
X_5494_ _5494_/A _5494_/B vssd1 vssd1 vccd1 vccd1 _5496_/A sky130_fd_sc_hd__nor2_1
Xhold157 _6182_/Q vssd1 vssd1 vccd1 vccd1 hold157/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold146 _4473_/X vssd1 vssd1 vccd1 vccd1 _6185_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 _4491_/X vssd1 vssd1 vccd1 vccd1 _6201_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4445_ _4438_/A _5301_/B _4123_/Y vssd1 vssd1 vccd1 vccd1 _4445_/X sky130_fd_sc_hd__a21o_1
Xhold179 _6246_/Q vssd1 vssd1 vccd1 vccd1 _3493_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4376_ hold183/X _4240_/X _4376_/S vssd1 vssd1 vccd1 vccd1 _4376_/X sky130_fd_sc_hd__mux2_1
X_3327_ _5617_/A vssd1 vssd1 vccd1 vccd1 _3405_/A sky130_fd_sc_hd__inv_2
X_6115_ _6399_/CLK _6115_/D vssd1 vssd1 vccd1 vccd1 _6115_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3258_ _3691_/B _3258_/B vssd1 vssd1 vccd1 vccd1 _3278_/A sky130_fd_sc_hd__nand2_2
XANTENNA__5652__A1 _5757_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6046_ _5567_/B _6045_/X _6071_/S vssd1 vssd1 vccd1 vccd1 _6046_/X sky130_fd_sc_hd__o21a_1
XANTENNA__5888__S _5977_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3189_ _6299_/Q _6300_/Q vssd1 vssd1 vccd1 vccd1 _3376_/B sky130_fd_sc_hd__nand2b_2
XFILLER_0_95_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5707__A2 _5721_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3156__B _3168_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3172__A _3172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4268__A _4268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4446__A2 _4462_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6247__RESET_B fanout180/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4230_ hold11/X _4462_/A2 _4463_/S vssd1 vssd1 vccd1 vccd1 _4230_/X sky130_fd_sc_hd__o21a_1
X_4161_ _4203_/A _4162_/A _4162_/B vssd1 vssd1 vccd1 vccd1 _4161_/X sky130_fd_sc_hd__a21o_1
XANTENNA__3082__A _6380_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4092_ _4096_/B _4092_/B vssd1 vssd1 vccd1 vccd1 _4095_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_65_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3112_ _4792_/A vssd1 vssd1 vccd1 vccd1 _4802_/A sky130_fd_sc_hd__inv_2
XANTENNA__3232__D _4248_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3810__A _3852_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5820__A1_N _5977_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4994_ _6370_/Q _5848_/S _5972_/B1 _4993_/X vssd1 vssd1 vccd1 vccd1 _4994_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_58_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3945_ _6219_/Q _3804_/X _3807_/X _6135_/Q vssd1 vssd1 vccd1 vccd1 _3945_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_45_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5615_ _4675_/A _5605_/D _4585_/Y _3590_/A _5364_/A vssd1 vssd1 vccd1 vccd1 _5615_/Y
+ sky130_fd_sc_hd__a221oi_1
X_3876_ _3883_/S _3874_/X _3875_/X _3816_/B vssd1 vssd1 vccd1 vccd1 _3878_/C sky130_fd_sc_hd__a211o_1
XFILLER_0_83_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5546_ hold541/X _5520_/B _5545_/Y _5415_/X vssd1 vssd1 vccd1 vccd1 _5546_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_14_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5477_ _5757_/A _6463_/Q vssd1 vssd1 vccd1 vccd1 _5479_/B sky130_fd_sc_hd__or2_1
X_4428_ _4441_/S _4424_/X _4426_/X _4427_/X vssd1 vssd1 vccd1 vccd1 _4428_/X sky130_fd_sc_hd__a22o_2
XANTENNA__5873__A1 _5976_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4359_ _5522_/A _4359_/B _4359_/C vssd1 vssd1 vccd1 vccd1 _4361_/B sky130_fd_sc_hd__and3_2
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6029_ _3700_/A _6026_/S _6023_/Y _5478_/S vssd1 vssd1 vccd1 vccd1 _6029_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_5_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6412_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_68_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6050__A1 _5567_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold516_A _6469_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout63 _5874_/S vssd1 vssd1 vccd1 vccd1 _5977_/S sky130_fd_sc_hd__clkbuf_8
Xfanout74 _5731_/C1 vssd1 vssd1 vccd1 vccd1 _5721_/C1 sky130_fd_sc_hd__buf_6
XFILLER_0_91_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout96 _3297_/B vssd1 vssd1 vccd1 vccd1 _4595_/B sky130_fd_sc_hd__buf_4
Xfanout85 _3700_/Y vssd1 vssd1 vccd1 vccd1 _4462_/A2 sky130_fd_sc_hd__clkbuf_8
XANTENNA__3167__A _3205_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4697__S _4711_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4667__A2 _4652_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5864__A1 _6021_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6428__RESET_B fanout172/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4419__A2 _4408_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6041__A1 _6101_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6041__B2 _6036_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3730_ _3712_/Y _3715_/Y _3725_/X _3728_/X vssd1 vssd1 vccd1 vccd1 _3861_/S sky130_fd_sc_hd__o31a_4
XFILLER_0_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3661_ _6283_/Q _3098_/Y _6168_/Q vssd1 vssd1 vccd1 vccd1 _3661_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_0_82_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3592_ _5777_/A _3285_/B _5777_/B _3591_/X vssd1 vssd1 vccd1 vccd1 _3592_/X sky130_fd_sc_hd__o31a_1
X_5400_ _5400_/A _5400_/B vssd1 vssd1 vccd1 vccd1 _5400_/X sky130_fd_sc_hd__or2_1
X_6380_ _6465_/CLK _6380_/D vssd1 vssd1 vccd1 vccd1 _6380_/Q sky130_fd_sc_hd__dfxtp_2
X_5331_ _4289_/C _5325_/X _5330_/X hold604/X _5322_/Y vssd1 vssd1 vccd1 vccd1 _5331_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_11_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3805__A _3852_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5262_ _5262_/A _5262_/B _5262_/C _5262_/D vssd1 vssd1 vccd1 vccd1 _5263_/C sky130_fd_sc_hd__or4_1
X_5193_ _6288_/Q _6289_/Q vssd1 vssd1 vccd1 vccd1 _5194_/B sky130_fd_sc_hd__xor2_1
X_4213_ _4203_/A _5178_/B _4212_/X _4211_/A vssd1 vssd1 vccd1 vccd1 _4213_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_76_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3866__B1 _3852_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4144_ _4144_/A _4144_/B vssd1 vssd1 vccd1 vccd1 _4146_/B sky130_fd_sc_hd__or2_2
XANTENNA__5607__B2 _5607_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4075_ _6288_/Q _3770_/A _4074_/X _6382_/Q _4072_/X vssd1 vssd1 vccd1 vccd1 _4075_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5231__S _5292_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4815__C1 _5783_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4977_ hold361/X _4976_/X _5016_/S vssd1 vssd1 vccd1 vccd1 _4977_/X sky130_fd_sc_hd__mux2_1
X_3928_ _3928_/A _3928_/B vssd1 vssd1 vccd1 vccd1 _3928_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_73_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3859_ _3892_/A _3859_/B vssd1 vssd1 vccd1 vccd1 _4430_/B sky130_fd_sc_hd__nor2_1
XANTENNA__4346__B2 _3284_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5529_ _6484_/Q _4982_/B _5593_/S vssd1 vssd1 vccd1 vccd1 _5531_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_41_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4310__S _4310_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4353__A1_N _6435_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3388__A2 _3497_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4034__B1 _3810_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5782__B1 _5418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5808__C _5866_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4337__A1 _5605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4900_ _4899_/X _4898_/X _5101_/S vssd1 vssd1 vccd1 vccd1 _4901_/B sky130_fd_sc_hd__mux2_2
X_5880_ _5866_/A _6465_/Q _5866_/C _5867_/B vssd1 vssd1 vccd1 vccd1 _5901_/B sky130_fd_sc_hd__o31a_2
XFILLER_0_87_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4831_ _5109_/A1 _4827_/X _4830_/Y _4924_/C vssd1 vssd1 vccd1 vccd1 _4831_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4576__A1 _4595_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4762_ hold512/X _4320_/A _4768_/S vssd1 vssd1 vccd1 vccd1 _4762_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_83_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4693_ _6385_/Q _4692_/X _4712_/S vssd1 vssd1 vccd1 vccd1 _4693_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_70_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3713_ _5295_/A _3711_/Y _3687_/X _5296_/A vssd1 vssd1 vccd1 vccd1 _3714_/S sky130_fd_sc_hd__a211o_1
XFILLER_0_15_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6432_ _6439_/CLK _6432_/D fanout178/X vssd1 vssd1 vccd1 vccd1 _6432_/Q sky130_fd_sc_hd__dfrtp_4
X_3644_ _5295_/A _6474_/Q _3644_/C vssd1 vssd1 vccd1 vccd1 _3647_/C sky130_fd_sc_hd__or3_1
XFILLER_0_15_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3575_ _5605_/A _4264_/B vssd1 vssd1 vccd1 vccd1 _3575_/Y sky130_fd_sc_hd__nand2_1
X_6363_ _6475_/CLK _6363_/D fanout175/X vssd1 vssd1 vccd1 vccd1 _6363_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_3_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6294_ _6446_/CLK _6294_/D fanout184/X vssd1 vssd1 vccd1 vccd1 _6294_/Q sky130_fd_sc_hd__dfrtp_1
X_5314_ _5360_/C _4325_/A _5314_/S vssd1 vssd1 vccd1 vccd1 _5314_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_3_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5245_ _6280_/Q wire92/X _5123_/Y _5244_/X vssd1 vssd1 vccd1 vccd1 _5245_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_46_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold28 hold28/A vssd1 vssd1 vccd1 vccd1 hold28/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold17 hold17/A vssd1 vssd1 vccd1 vccd1 hold17/X sky130_fd_sc_hd__dlygate4sd3_1
X_5176_ _5176_/A _5176_/B vssd1 vssd1 vccd1 vccd1 _5177_/B sky130_fd_sc_hd__xnor2_1
Xhold39 hold39/A vssd1 vssd1 vccd1 vccd1 hold39/X sky130_fd_sc_hd__dlygate4sd3_1
X_4127_ _6116_/Q _3731_/X _3810_/X _6183_/Q _4126_/X vssd1 vssd1 vccd1 vccd1 _4128_/B
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4366__A _4366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4058_ _6287_/Q _6289_/Q _4716_/A vssd1 vssd1 vccd1 vccd1 _5262_/C sky130_fd_sc_hd__mux2_1
XFILLER_0_78_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5764__A0 _6315_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4567__A1 _6316_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3148__C _5369_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3790__A2 _5317_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5644__B _5734_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5819__B2 _5786_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5819__A1 _5976_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3180__A _3304_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4276__A _4276_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xci2406_z80_207 vssd1 vssd1 vccd1 vccd1 ci2406_z80_207/HI io_oeb[32] sky130_fd_sc_hd__conb_1
XFILLER_0_69_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4723__B _5757_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold509 _5701_/X vssd1 vssd1 vccd1 vccd1 _6382_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_33_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3360_ _3547_/B _3360_/B vssd1 vssd1 vccd1 vccd1 _4073_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_0_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3291_ _4338_/A _3285_/D _3668_/A _3581_/B _3352_/B vssd1 vssd1 vccd1 vccd1 _3291_/X
+ sky130_fd_sc_hd__o221a_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5030_ _5109_/A1 _5025_/X _5029_/X _4924_/C vssd1 vssd1 vccd1 vccd1 _5030_/X sky130_fd_sc_hd__a22o_1
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5691__C1 _5730_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3090__A _6309_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3802__B _3818_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5932_ _5933_/A _5970_/A vssd1 vssd1 vccd1 vccd1 _5934_/A sky130_fd_sc_hd__nand2_1
X_5863_ _6367_/Q _5862_/X _5863_/S vssd1 vssd1 vccd1 vccd1 _5863_/X sky130_fd_sc_hd__mux2_1
X_5794_ _5786_/Y _5789_/Y _5793_/Y _5976_/S vssd1 vssd1 vccd1 vccd1 _5794_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_28_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4814_ _6361_/Q _5861_/S _5842_/B1 _4813_/X _5102_/A vssd1 vssd1 vccd1 vccd1 _4814_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4013__A3 _6287_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4745_ _4743_/X _4744_/X _5289_/S vssd1 vssd1 vccd1 vccd1 _4745_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_16_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4676_ _4676_/A _4676_/B vssd1 vssd1 vccd1 vccd1 _4711_/S sky130_fd_sc_hd__and2_4
XFILLER_0_98_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3627_ _5322_/A _3627_/B _3627_/C _3674_/A vssd1 vssd1 vccd1 vccd1 _5294_/B sky130_fd_sc_hd__or4_4
X_6415_ _6417_/CLK _6415_/D fanout174/X vssd1 vssd1 vccd1 vccd1 _6415_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__5464__B _6462_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3558_ _5309_/A _5770_/B vssd1 vssd1 vccd1 vccd1 _3674_/B sky130_fd_sc_hd__nand2_1
X_6346_ _6441_/CLK _6346_/D fanout184/X vssd1 vssd1 vccd1 vccd1 _6346_/Q sky130_fd_sc_hd__dfrtp_4
Xoutput29 _6322_/Q vssd1 vssd1 vccd1 vccd1 io_out[11] sky130_fd_sc_hd__buf_12
XFILLER_0_11_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3489_ _5145_/A _3489_/B _3489_/C vssd1 vssd1 vccd1 vccd1 _3489_/Y sky130_fd_sc_hd__nor3_1
X_6277_ _6383_/CLK _6277_/D fanout182/X vssd1 vssd1 vccd1 vccd1 _6277_/Q sky130_fd_sc_hd__dfstp_1
X_5228_ _6336_/Q _5202_/A _5227_/X _5290_/S vssd1 vssd1 vccd1 vccd1 _5228_/X sky130_fd_sc_hd__a211o_1
XANTENNA__4096__A _4150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5159_ _4193_/B _4196_/Y _5158_/X vssd1 vssd1 vccd1 vccd1 _5159_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__5682__C1 _5721_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4824__A _5064_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_hold429_A _6381_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3874__S _3884_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5060__S1 _5100_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_45_wb_clk_i_A clkbuf_leaf_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_27_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5821__C _5866_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4228__B1 _3701_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xmax_cap71 _3723_/Y vssd1 vssd1 vccd1 vccd1 _3885_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_84_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5268__C _6289_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4530_ hold83/X _4416_/X _4536_/S vssd1 vssd1 vccd1 vccd1 hold84/A sky130_fd_sc_hd__mux2_1
XFILLER_0_13_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4951__A1 _5109_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold306 hold658/X vssd1 vssd1 vccd1 vccd1 hold306/X sky130_fd_sc_hd__buf_1
Xhold317 _4695_/X vssd1 vssd1 vccd1 vccd1 _6304_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4461_ _4438_/A _5302_/C _4228_/X vssd1 vssd1 vccd1 vccd1 _4461_/X sky130_fd_sc_hd__a21o_1
X_3412_ _4313_/A _3412_/B vssd1 vssd1 vccd1 vccd1 _3412_/Y sky130_fd_sc_hd__nor2_1
Xhold328 _6132_/Q vssd1 vssd1 vccd1 vccd1 hold328/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3085__A _6459_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold339 _4295_/X vssd1 vssd1 vccd1 vccd1 _6120_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6200_ _6265_/CLK _6200_/D vssd1 vssd1 vccd1 vccd1 _6200_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6131_ _6242_/CLK hold60/X fanout180/X vssd1 vssd1 vccd1 vccd1 hold59/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4392_ hold93/X _3998_/X _4397_/S vssd1 vssd1 vccd1 vccd1 hold94/A sky130_fd_sc_hd__mux2_1
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3343_ _6431_/Q _3320_/Y _3106_/A vssd1 vssd1 vccd1 vccd1 _3343_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5504__S _5593_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3274_ _3187_/X _3274_/B _3274_/C vssd1 vssd1 vccd1 vccd1 _3274_/X sky130_fd_sc_hd__and3b_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6062_ _6101_/A _6061_/X _6071_/S vssd1 vssd1 vccd1 vccd1 _6062_/X sky130_fd_sc_hd__o21a_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5013_ _5102_/A _5012_/Y _5002_/Y vssd1 vssd1 vccd1 vccd1 _5013_/X sky130_fd_sc_hd__o21a_1
XANTENNA__3690__B2 _5777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5967__B1 _5784_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout167_A _5078_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5915_ _5915_/A _5915_/B vssd1 vssd1 vccd1 vccd1 _5915_/X sky130_fd_sc_hd__or2_1
X_5846_ _5977_/S _5845_/X _5784_/X hold379/X vssd1 vssd1 vccd1 vccd1 _5846_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_91_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5777_ _5777_/A _5777_/B _3522_/X vssd1 vssd1 vccd1 vccd1 _5777_/X sky130_fd_sc_hd__or3b_1
XFILLER_0_8_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6365__RESET_B fanout181/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4728_ _3782_/Y _4727_/X _4770_/S vssd1 vssd1 vccd1 vccd1 _4728_/X sky130_fd_sc_hd__mux2_1
X_4659_ _4782_/B _4652_/X _4654_/Y _4658_/X vssd1 vssd1 vccd1 vccd1 _6295_/D sky130_fd_sc_hd__o22a_1
XFILLER_0_71_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5922__B _5970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6329_ _6407_/CLK _6329_/D fanout170/X vssd1 vssd1 vccd1 vccd1 _6329_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__5670__A2 _5655_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3869__S _3884_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5369__B _5369_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_1_wb_clk_i_A clkbuf_leaf_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_10_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4697__A0 _6382_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3352__B _3352_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3672__A1 _3674_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_29_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6316_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__5279__B _6458_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3961_ _3961_/A _3961_/B vssd1 vssd1 vccd1 vccd1 _3962_/B sky130_fd_sc_hd__or2_2
X_5700_ _5700_/A _5700_/B _5700_/C vssd1 vssd1 vccd1 vccd1 _5700_/X sky130_fd_sc_hd__or3_1
XFILLER_0_85_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3892_ _3892_/A _3892_/B vssd1 vssd1 vccd1 vccd1 _4425_/B sky130_fd_sc_hd__xnor2_1
X_5631_ _5644_/A _5645_/A _5610_/B vssd1 vssd1 vccd1 vccd1 _5632_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_5_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5562_ _5562_/A _5562_/B vssd1 vssd1 vccd1 vccd1 _5565_/A sky130_fd_sc_hd__or2_1
XANTENNA__3808__A _3884_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4513_ _3998_/X hold309/X _4518_/S vssd1 vssd1 vccd1 vccd1 _6220_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_41_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold103 _6146_/Q vssd1 vssd1 vccd1 vccd1 hold103/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold114 _6148_/Q vssd1 vssd1 vccd1 vccd1 hold114/X sky130_fd_sc_hd__dlygate4sd3_1
X_5493_ _5492_/A _5492_/B _5492_/C vssd1 vssd1 vccd1 vccd1 _5494_/B sky130_fd_sc_hd__a21oi_1
Xhold125 _6172_/Q vssd1 vssd1 vccd1 vccd1 hold125/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold147 _6197_/Q vssd1 vssd1 vccd1 vccd1 hold147/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold158 _4470_/X vssd1 vssd1 vccd1 vccd1 _6182_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold136 _6179_/Q vssd1 vssd1 vccd1 vccd1 hold136/X sky130_fd_sc_hd__dlygate4sd3_1
X_4444_ _4444_/A _4444_/B vssd1 vssd1 vccd1 vccd1 _5301_/B sky130_fd_sc_hd__xnor2_1
X_4375_ hold111/X _4182_/X _4376_/S vssd1 vssd1 vccd1 vccd1 _4375_/X sky130_fd_sc_hd__mux2_1
Xhold169 _6455_/Q vssd1 vssd1 vccd1 vccd1 hold169/X sky130_fd_sc_hd__dlygate4sd3_1
X_3326_ _3326_/A _3326_/B _3216_/B vssd1 vssd1 vccd1 vccd1 _5617_/A sky130_fd_sc_hd__or3b_4
X_6114_ _6223_/CLK _6114_/D vssd1 vssd1 vccd1 vccd1 _6114_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6045_ _6101_/B _4822_/X _5433_/Y _6036_/X vssd1 vssd1 vccd1 vccd1 _6045_/X sky130_fd_sc_hd__o22a_1
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3257_ _3691_/B _3258_/B vssd1 vssd1 vccd1 vccd1 _3581_/B sky130_fd_sc_hd__and2_2
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3188_ _6299_/Q _6300_/Q vssd1 vssd1 vccd1 vccd1 _3219_/A sky130_fd_sc_hd__and2b_2
XFILLER_0_95_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3415__B2 _3674_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5829_ _6364_/Q _5861_/S _5842_/B1 _5828_/X vssd1 vssd1 vccd1 vccd1 _5829_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_44_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4679__B1 _4714_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5340__A1 _6297_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4143__A2 _3731_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5144__S _5232_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6483__SET_B fanout176/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3654__A1 _4325_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3406__A1 _5317_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3957__A2 _3799_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4906__B2 _4901_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5331__B2 hold604/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4160_ _6290_/Q _4205_/S vssd1 vssd1 vccd1 vccd1 _4162_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__3363__A _4716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3111_ _3699_/A hold347/X _3554_/A _4324_/A vssd1 vssd1 vccd1 vccd1 _4792_/A sky130_fd_sc_hd__o31a_2
XANTENNA__4178__B _6067_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4091_ _6289_/Q _4091_/B _4091_/C vssd1 vssd1 vccd1 vccd1 _4092_/B sky130_fd_sc_hd__nor3_1
XANTENNA__5634__A2 _4406_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3810__B _3883_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4993_ _6403_/Q _4992_/X _5971_/S vssd1 vssd1 vccd1 vccd1 _4993_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_81_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3944_ _6260_/Q _3793_/X _3795_/X _6195_/Q vssd1 vssd1 vccd1 vccd1 _3947_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_18_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4922__A _6366_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3875_ hold83/X _3861_/S _3873_/X _3723_/Y vssd1 vssd1 vccd1 vccd1 _3875_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_18_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6103__A1_N _6067_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4641__B _4641_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5614_ _6432_/Q _4595_/B _3489_/B vssd1 vssd1 vccd1 vccd1 _5614_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_5_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5545_ _5545_/A _5545_/B vssd1 vssd1 vccd1 vccd1 _5545_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_30_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5476_ hold595/X _5475_/X _5513_/S vssd1 vssd1 vccd1 vccd1 _5476_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4125__A2 _3799_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4427_ hold29/X _3700_/Y _3698_/Y vssd1 vssd1 vccd1 vccd1 _4427_/X sky130_fd_sc_hd__o21a_1
XANTENNA__4088__B _6383_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4358_ _5522_/A _4358_/B vssd1 vssd1 vccd1 vccd1 _6101_/B sky130_fd_sc_hd__nand2_8
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3309_ _5600_/B _3609_/A vssd1 vssd1 vccd1 vccd1 _3394_/A sky130_fd_sc_hd__or2_1
X_4289_ _4716_/A _4289_/B _4289_/C vssd1 vssd1 vccd1 vccd1 _4768_/S sky130_fd_sc_hd__and3_4
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6028_ _5478_/S _6026_/S _6023_/Y _3501_/A vssd1 vssd1 vccd1 vccd1 _6469_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_96_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout64 _5887_/S vssd1 vssd1 vccd1 vccd1 _5976_/S sky130_fd_sc_hd__clkbuf_8
XANTENNA_hold411_A _6329_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout97 _5360_/B vssd1 vssd1 vccd1 vccd1 _5314_/S sky130_fd_sc_hd__buf_4
XFILLER_0_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout86 _3698_/Y vssd1 vssd1 vccd1 vccd1 _4463_/S sky130_fd_sc_hd__buf_6
Xfanout75 _3908_/X vssd1 vssd1 vccd1 vccd1 _5731_/C1 sky130_fd_sc_hd__clkbuf_8
XANTENNA__4043__S _4241_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3882__S _3884_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6041__A2 _5413_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3660_ _6168_/Q _6165_/Q input4/X vssd1 vssd1 vccd1 vccd1 _3660_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_70_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3591_ _4338_/A _4386_/A _3673_/B _3588_/Y _3590_/Y vssd1 vssd1 vccd1 vccd1 _3591_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_23_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5330_ _4217_/A _5314_/X _5328_/X _5329_/X vssd1 vssd1 vccd1 vccd1 _5330_/X sky130_fd_sc_hd__a211o_1
X_5261_ _6284_/Q _5261_/B _5261_/C _5170_/B vssd1 vssd1 vccd1 vccd1 _5261_/X sky130_fd_sc_hd__or4b_1
XFILLER_0_11_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3805__B _3885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4212_ _4212_/A _4212_/B vssd1 vssd1 vccd1 vccd1 _4212_/X sky130_fd_sc_hd__or2_1
XANTENNA__3093__A _6314_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5192_ _5192_/A _5192_/B vssd1 vssd1 vccd1 vccd1 _5195_/A sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_44_wb_clk_i clkbuf_leaf_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6263_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__3866__A1 _3885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4143_ _6117_/Q _3731_/X _3810_/X _6184_/Q _4142_/X vssd1 vssd1 vccd1 vccd1 _4144_/B
+ sky130_fd_sc_hd__a221o_1
X_4074_ _4073_/A _4223_/A _4073_/Y _3759_/Y vssd1 vssd1 vccd1 vccd1 _4074_/X sky130_fd_sc_hd__a211o_1
XANTENNA__4636__B _4641_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4652__A _5769_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4976_ _6458_/Q _4975_/X _5974_/S vssd1 vssd1 vccd1 vccd1 _4976_/X sky130_fd_sc_hd__mux2_1
X_3927_ _3986_/A _4720_/C vssd1 vssd1 vccd1 vccd1 _3927_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_73_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3858_ _3892_/A _3859_/B vssd1 vssd1 vccd1 vccd1 _3858_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__4346__A2 _3668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3789_ _3278_/A _3674_/A _3693_/C _3278_/B vssd1 vssd1 vccd1 vccd1 _3789_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_6_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5528_ _5526_/X _5527_/X _4300_/A _5521_/A vssd1 vssd1 vccd1 vccd1 _5528_/X sky130_fd_sc_hd__a2bb2o_1
X_5459_ _5457_/X _5458_/X _5485_/S vssd1 vssd1 vccd1 vccd1 _5459_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_1_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3490__C1 _4800_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold626_A _6460_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3178__A _4268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3906__A _6355_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4830_ _4847_/B _4830_/B vssd1 vssd1 vccd1 vccd1 _4830_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__5222__A0 _6336_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4761_ _6315_/Q _4719_/A _4760_/X _4957_/S vssd1 vssd1 vccd1 vccd1 _4761_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_28_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4692_ _6381_/Q _6287_/Q _4711_/S vssd1 vssd1 vccd1 vccd1 _4692_/X sky130_fd_sc_hd__mux2_1
X_3712_ _5295_/A _3711_/Y _3687_/X _5296_/A vssd1 vssd1 vccd1 vccd1 _3712_/Y sky130_fd_sc_hd__a211oi_4
XFILLER_0_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3643_ _5405_/B _3643_/B vssd1 vssd1 vccd1 vccd1 _3644_/C sky130_fd_sc_hd__or2_2
X_6431_ _6444_/CLK _6431_/D fanout178/X vssd1 vssd1 vccd1 vccd1 _6431_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_43_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4959__S0 _5100_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6362_ _6462_/CLK _6362_/D fanout181/X vssd1 vssd1 vccd1 vccd1 _6362_/Q sky130_fd_sc_hd__dfrtp_4
X_5313_ _3986_/A _5336_/B _5336_/A _4247_/B vssd1 vssd1 vccd1 vccd1 _5313_/X sky130_fd_sc_hd__a211o_1
X_3574_ _6435_/Q _3574_/B _5146_/D vssd1 vssd1 vccd1 vccd1 _3574_/X sky130_fd_sc_hd__or3_1
XFILLER_0_3_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6293_ _6446_/CLK _6293_/D fanout184/X vssd1 vssd1 vccd1 vccd1 _6293_/Q sky130_fd_sc_hd__dfrtp_1
X_5244_ _6314_/Q _5243_/X _5244_/S vssd1 vssd1 vccd1 vccd1 _5244_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_11_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5175_ _5260_/B _5175_/B vssd1 vssd1 vccd1 vccd1 _5176_/B sky130_fd_sc_hd__xnor2_1
Xhold29 hold29/A vssd1 vssd1 vccd1 vccd1 hold29/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold18 hold18/A vssd1 vssd1 vccd1 vccd1 hold18/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5242__S _5489_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4126_ _6223_/Q _3804_/X _3807_/X _6139_/Q vssd1 vssd1 vccd1 vccd1 _4126_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_39_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4057_ _5260_/A _5174_/A vssd1 vssd1 vccd1 vccd1 _4057_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_78_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4959_ _6151_/Q _6134_/Q _6142_/Q _6178_/Q _5100_/S1 _5100_/S0 vssd1 vssd1 vccd1
+ vccd1 _4959_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_19_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_35_wb_clk_i_A clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_100_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4557__A _5322_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3120__A_N _3284_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4276__B _5314_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xci2406_z80_208 vssd1 vssd1 vccd1 vccd1 ci2406_z80_208/HI io_oeb[33] sky130_fd_sc_hd__conb_1
XFILLER_0_96_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5388__A _5388_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4292__A _4313_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5835__B _5867_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3636__A _4800_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3290_ _4335_/B _3786_/A vssd1 vssd1 vccd1 vccd1 _3668_/A sky130_fd_sc_hd__or2_4
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5851__A _5866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5691__B1 _5721_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5931_ _5922_/A _5930_/X _5977_/S vssd1 vssd1 vccd1 vccd1 _5931_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_48_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5862_ _5817_/A _5861_/X _4920_/X vssd1 vssd1 vccd1 vccd1 _5862_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_75_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5793_ _5804_/A _5793_/B vssd1 vssd1 vccd1 vccd1 _5793_/Y sky130_fd_sc_hd__nand2_1
X_4813_ _6361_/Q _4812_/X _5892_/S vssd1 vssd1 vccd1 vccd1 _4813_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4744_ hold407/X _4312_/A _4768_/S vssd1 vssd1 vccd1 vccd1 _4744_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_83_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4675_ _4675_/A _5146_/C _4675_/C vssd1 vssd1 vccd1 vccd1 _4712_/S sky130_fd_sc_hd__or3_4
X_3626_ _3665_/A _5757_/A _3600_/X _3625_/Y vssd1 vssd1 vccd1 vccd1 _6168_/D sky130_fd_sc_hd__a31o_1
X_6414_ _6417_/CLK _6414_/D fanout174/X vssd1 vssd1 vccd1 vccd1 _6414_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA_fanout112_A _6108_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6345_ _6446_/CLK _6345_/D fanout184/X vssd1 vssd1 vccd1 vccd1 _6345_/Q sky130_fd_sc_hd__dfrtp_4
X_3557_ _4335_/B _3557_/B _3668_/B vssd1 vssd1 vccd1 vccd1 _3557_/X sky130_fd_sc_hd__or3_1
Xoutput19 _6523_/X vssd1 vssd1 vccd1 vccd1 io_oeb[22] sky130_fd_sc_hd__buf_12
X_6276_ _6312_/CLK _6276_/D fanout183/X vssd1 vssd1 vccd1 vccd1 _6276_/Q sky130_fd_sc_hd__dfstp_1
X_3488_ _3488_/A _3488_/B vssd1 vssd1 vccd1 vccd1 _3489_/C sky130_fd_sc_hd__nand2_1
X_5227_ _6381_/Q _5314_/S _4223_/A _4020_/X vssd1 vssd1 vccd1 vccd1 _5227_/X sky130_fd_sc_hd__a31o_1
XANTENNA__3281__A _3281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3288__A2 _5317_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5682__B1 _5721_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5158_ _5268_/A _5158_/B _4193_/B vssd1 vssd1 vccd1 vccd1 _5158_/X sky130_fd_sc_hd__or3b_1
X_4109_ _6289_/Q _4109_/B vssd1 vssd1 vccd1 vccd1 _4210_/A sky130_fd_sc_hd__xor2_1
X_5089_ _6464_/Q _5108_/S _5088_/X vssd1 vssd1 vccd1 vccd1 _5089_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_94_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4824__B _4835_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3748__A0 _4150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5655__B _5655_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3763__A3 _4557_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5374__C _5374_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5268__D _6290_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5728__A1 _6340_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3366__A _4716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4460_ _4460_/A _4460_/B vssd1 vssd1 vccd1 vccd1 _5302_/C sky130_fd_sc_hd__xnor2_1
Xhold307 _6123_/Q vssd1 vssd1 vccd1 vccd1 _4312_/A sky130_fd_sc_hd__clkbuf_2
X_3411_ _3411_/A _5406_/B vssd1 vssd1 vccd1 vccd1 _3411_/Y sky130_fd_sc_hd__nand2_1
Xhold329 _3526_/X vssd1 vssd1 vccd1 vccd1 _6132_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold318 _6306_/Q vssd1 vssd1 vccd1 vccd1 hold318/X sky130_fd_sc_hd__dlygate4sd3_1
X_4391_ hold161/X _3954_/X _4397_/S vssd1 vssd1 vccd1 vccd1 _4391_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_7_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3342_ _6430_/Q _3332_/A _3310_/Y vssd1 vssd1 vccd1 vccd1 _3342_/X sky130_fd_sc_hd__o21a_1
X_6130_ _6242_/CLK _6130_/D fanout180/X vssd1 vssd1 vccd1 vccd1 _6130_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4197__A _5268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3273_ _3273_/A _3273_/B _3273_/C vssd1 vssd1 vccd1 vccd1 _3274_/C sky130_fd_sc_hd__and3_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6061_ _6101_/B _4901_/B _5483_/X _6036_/X vssd1 vssd1 vccd1 vccd1 _6061_/X sky130_fd_sc_hd__o22a_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3532__C _5777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5012_ _6371_/Q _5848_/S _5972_/B1 _5011_/X vssd1 vssd1 vccd1 vccd1 _5012_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_0_84_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4219__B2 _5268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4219__A1 _6333_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5914_ _5914_/A _5914_/B _5914_/C vssd1 vssd1 vccd1 vccd1 _5915_/B sky130_fd_sc_hd__and3_1
XFILLER_0_91_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5845_ _5887_/S _5840_/Y _5844_/Y _5786_/Y vssd1 vssd1 vccd1 vccd1 _5845_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_36_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4660__A input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5776_ _3627_/B _3627_/C _4386_/B _5775_/Y _5387_/C vssd1 vssd1 vccd1 vccd1 _5776_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_0_44_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4727_ _4722_/X _4726_/X _5289_/S vssd1 vssd1 vccd1 vccd1 _4727_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_44_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4658_ _4658_/A _4668_/B vssd1 vssd1 vccd1 vccd1 _4658_/X sky130_fd_sc_hd__and2_1
XFILLER_0_31_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3609_ _3609_/A _5370_/B _3609_/C vssd1 vssd1 vccd1 vccd1 _5523_/A sky130_fd_sc_hd__or3_2
XFILLER_0_31_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4589_ _3185_/A _5777_/B _4253_/A vssd1 vssd1 vccd1 vccd1 _4589_/Y sky130_fd_sc_hd__o21ai_1
X_6328_ _6407_/CLK _6328_/D fanout170/X vssd1 vssd1 vccd1 vccd1 _6328_/Q sky130_fd_sc_hd__dfrtp_2
X_6259_ _6399_/CLK _6259_/D vssd1 vssd1 vccd1 vccd1 _6259_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__6080__B1 _6107_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4630__B2 _4629_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4720__D _6021_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4697__A1 _6378_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3633__B _4788_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6071__A0 _4227_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3960_ _6113_/Q _3731_/X _3810_/X _6180_/Q _3959_/X vssd1 vssd1 vccd1 vccd1 _3961_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_85_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4621__A1 _4036_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3891_ _3892_/A _3892_/B vssd1 vssd1 vccd1 vccd1 _3891_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_38_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5630_ _5644_/A _5645_/A _5645_/B _5630_/D vssd1 vssd1 vccd1 vccd1 _5630_/X sky130_fd_sc_hd__and4_2
XFILLER_0_5_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5561_ _5594_/A _5561_/B vssd1 vssd1 vccd1 vccd1 _5562_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_5_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4512_ _3954_/X hold218/X _4518_/S vssd1 vssd1 vccd1 vccd1 _4512_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_26_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5492_ _5492_/A _5492_/B _5492_/C vssd1 vssd1 vccd1 vccd1 _5494_/A sky130_fd_sc_hd__and3_1
XFILLER_0_80_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold126 _6210_/Q vssd1 vssd1 vccd1 vccd1 hold126/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold104 _4382_/X vssd1 vssd1 vccd1 vccd1 _6146_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold115 _4384_/X vssd1 vssd1 vccd1 vccd1 _6148_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold148 _4487_/X vssd1 vssd1 vccd1 vccd1 _6197_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold137 _4467_/X vssd1 vssd1 vccd1 vccd1 _6179_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5515__S _5593_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4443_ _4190_/A _3847_/B _3898_/C vssd1 vssd1 vccd1 vccd1 _4444_/B sky130_fd_sc_hd__a21oi_1
Xhold159 _6211_/Q vssd1 vssd1 vccd1 vccd1 hold159/X sky130_fd_sc_hd__dlygate4sd3_1
X_4374_ hold134/X _4138_/X _4376_/S vssd1 vssd1 vccd1 vccd1 _4374_/X sky130_fd_sc_hd__mux2_1
X_3325_ _3379_/A _3412_/B _4253_/A _3324_/Y _3617_/A vssd1 vssd1 vccd1 vccd1 _3329_/D
+ sky130_fd_sc_hd__o221a_1
X_6113_ _6263_/CLK _6113_/D vssd1 vssd1 vccd1 vccd1 _6113_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3256_ _3304_/B _3268_/B vssd1 vssd1 vccd1 vccd1 _3258_/B sky130_fd_sc_hd__or2_4
X_6044_ _5384_/A _6042_/X _6043_/Y hold417/X _6040_/Y vssd1 vssd1 vccd1 vccd1 _6044_/X
+ sky130_fd_sc_hd__o32a_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3187_ _3300_/A _3187_/B _5369_/C _3187_/D vssd1 vssd1 vccd1 vccd1 _3187_/X sky130_fd_sc_hd__or4_1
XFILLER_0_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5828_ _6364_/Q _6416_/Q _5892_/S vssd1 vssd1 vccd1 vccd1 _5828_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5759_ _6310_/Q hold456/X _5765_/S vssd1 vssd1 vccd1 vccd1 _5759_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_44_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5933__B _5970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3156__D _3205_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4679__A1 _4713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5340__A2 _5317_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold660 _6467_/Q vssd1 vssd1 vccd1 vccd1 hold660/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_hold489_A _6378_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5723__S0 _5655_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4851__A1 _6460_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4851__B2 _5109_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4504__S _4509_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3342__A1 _6430_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3110_ _3110_/A _3652_/B vssd1 vssd1 vccd1 vccd1 _3530_/A sky130_fd_sc_hd__and2_4
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4766__A1_N _6316_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4090_ _4091_/B _4091_/C _6289_/Q vssd1 vssd1 vccd1 vccd1 _4096_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_65_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4194__B _6385_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4992_ _6422_/Q _4793_/Y _4984_/X _4991_/X vssd1 vssd1 vccd1 vccd1 _4992_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_58_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3943_ _6152_/Q _3799_/X _3801_/X hold91/A vssd1 vssd1 vccd1 vccd1 _3947_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_18_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4922__B _6367_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3874_ hold79/X hold63/X _3884_/S vssd1 vssd1 vccd1 vccd1 _3874_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5613_ _5600_/A _5388_/A _4338_/X _4324_/X vssd1 vssd1 vccd1 vccd1 _5613_/X sky130_fd_sc_hd__a31o_1
X_5544_ _5545_/B vssd1 vssd1 vccd1 vccd1 _5544_/Y sky130_fd_sc_hd__inv_2
X_5475_ _6462_/Q _5474_/X _5512_/S vssd1 vssd1 vccd1 vccd1 _5475_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4426_ _4438_/A _3894_/B _4425_/Y _3995_/Y vssd1 vssd1 vccd1 vccd1 _4426_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_1_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4357_ _5522_/A _4359_/B _4357_/C vssd1 vssd1 vccd1 vccd1 _6100_/A sky130_fd_sc_hd__and3_2
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3308_ _5774_/B _3308_/B vssd1 vssd1 vccd1 vccd1 _4785_/A sky130_fd_sc_hd__or2_1
X_4288_ _4289_/B _4289_/C vssd1 vssd1 vccd1 vccd1 _4724_/C sky130_fd_sc_hd__and2_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3239_ _3314_/B _3632_/D vssd1 vssd1 vccd1 vccd1 _4784_/C sky130_fd_sc_hd__or2_1
X_6027_ _6468_/Q _6026_/S _6023_/Y _3594_/A vssd1 vssd1 vccd1 vccd1 _6027_/X sky130_fd_sc_hd__a22o_1
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4597__B1 _5607_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout65 _5842_/B1 vssd1 vssd1 vccd1 vccd1 _5972_/B1 sky130_fd_sc_hd__buf_4
XFILLER_0_36_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout98 _5892_/S vssd1 vssd1 vccd1 vccd1 _5971_/S sky130_fd_sc_hd__clkbuf_8
Xfanout87 _5817_/A vssd1 vssd1 vccd1 vccd1 _5964_/A sky130_fd_sc_hd__buf_4
Xfanout76 _3734_/X vssd1 vssd1 vccd1 vccd1 _4438_/A sky130_fd_sc_hd__buf_4
XANTENNA__5010__A1 _6423_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5155__S _5232_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3572__A1 _5314_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold490 _5652_/X vssd1 vssd1 vccd1 vccd1 _6378_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3639__A _5605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3358__B _4716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3590_ _3590_/A _5317_/B vssd1 vssd1 vccd1 vccd1 _3590_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_23_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3563__B2 _5146_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5260_ _5260_/A _5260_/B _5175_/B vssd1 vssd1 vccd1 vccd1 _5261_/C sky130_fd_sc_hd__or3b_1
XFILLER_0_23_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4211_ _4211_/A _4212_/B vssd1 vssd1 vccd1 vccd1 _5178_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_11_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5191_ _5267_/A _5267_/B vssd1 vssd1 vccd1 vccd1 _5192_/B sky130_fd_sc_hd__xor2_1
X_4142_ _6224_/Q _3804_/X _3807_/X _6140_/Q vssd1 vssd1 vccd1 vccd1 _4142_/X sky130_fd_sc_hd__a22o_1
X_4073_ _4073_/A _4168_/B vssd1 vssd1 vccd1 vccd1 _4073_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_78_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_13_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6242_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_78_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6017__A0 input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4652__B _5418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4975_ _5964_/A _4974_/X _4962_/Y vssd1 vssd1 vccd1 vccd1 _4975_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_25_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3926_ _6284_/Q _6286_/Q _4217_/A vssd1 vssd1 vccd1 vccd1 _5264_/B sky130_fd_sc_hd__mux2_1
XANTENNA__3549__A _5124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3857_ _3892_/A _3859_/B vssd1 vssd1 vccd1 vccd1 _4430_/A sky130_fd_sc_hd__and2_1
X_3788_ _3672_/X _3675_/X _3784_/Y _3787_/Y vssd1 vssd1 vccd1 vccd1 _3788_/Y sky130_fd_sc_hd__a31oi_4
XFILLER_0_26_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_25_wb_clk_i_A _6448_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5527_ _5593_/S _5411_/B _5525_/B _4300_/A vssd1 vssd1 vccd1 vccd1 _5527_/X sky130_fd_sc_hd__a31o_1
XANTENNA__3284__A _4782_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5458_ _4716_/A _6364_/Q _5484_/S vssd1 vssd1 vccd1 vccd1 _5458_/X sky130_fd_sc_hd__mux2_1
X_5389_ _5362_/C _4272_/X _5362_/D _5388_/X _4244_/Y vssd1 vssd1 vccd1 vccd1 _5391_/B
+ sky130_fd_sc_hd__o41a_1
X_4409_ hold63/X _4406_/B _4420_/S hold79/X _5731_/C1 vssd1 vssd1 vccd1 vccd1 _4409_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA__3731__B _3883_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4034__A2 _3731_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5782__A2 _5867_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3906__B _4441_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4258__C1 _5607_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output36_A _6329_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3136__C_N _3205_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5773__A2 _4248_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4760_ _6315_/Q _4720_/X _5224_/A2 _6273_/Q vssd1 vssd1 vccd1 vccd1 _4760_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_83_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4691_ _6089_/A _4714_/S vssd1 vssd1 vccd1 vccd1 _4691_/Y sky130_fd_sc_hd__nor2_1
X_3711_ _5607_/B2 _3689_/Y _3693_/X _5478_/S _3665_/A vssd1 vssd1 vccd1 vccd1 _3711_/Y
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_0_15_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3642_ _5522_/A _5478_/S _3642_/C _4357_/C vssd1 vssd1 vccd1 vccd1 _3650_/A sky130_fd_sc_hd__and4_1
XFILLER_0_70_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6430_ _6444_/CLK _6430_/D fanout178/X vssd1 vssd1 vccd1 vccd1 _6430_/Q sky130_fd_sc_hd__dfrtp_4
X_6361_ _6384_/CLK _6361_/D fanout175/X vssd1 vssd1 vccd1 vccd1 _6361_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_3_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4959__S1 _5100_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5312_ _5387_/C _3413_/Y _5311_/X vssd1 vssd1 vccd1 vccd1 _5336_/B sky130_fd_sc_hd__a21o_1
X_3573_ _3560_/X _3567_/X _3571_/X _3572_/Y _5322_/A vssd1 vssd1 vccd1 vccd1 _3573_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_0_87_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6292_ _6441_/CLK _6292_/D fanout185/X vssd1 vssd1 vccd1 vccd1 _6292_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__5289__A1 hold572/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5243_ _6338_/Q _3093_/Y _5243_/S vssd1 vssd1 vccd1 vccd1 _5243_/X sky130_fd_sc_hd__mux2_1
X_5174_ _5174_/A _5174_/B vssd1 vssd1 vccd1 vccd1 _5176_/A sky130_fd_sc_hd__xnor2_1
Xhold19 hold19/A vssd1 vssd1 vccd1 vccd1 hold19/X sky130_fd_sc_hd__dlygate4sd3_1
X_4125_ _6156_/Q _3799_/X _3801_/X _6147_/Q _4124_/X vssd1 vssd1 vccd1 vccd1 _4128_/A
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4139__S _4241_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4056_ _6288_/Q _4056_/B vssd1 vssd1 vccd1 vccd1 _5174_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_66_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4421__C1 _5731_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4958_ _4957_/X hold383/X _5098_/S vssd1 vssd1 vccd1 vccd1 _4958_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3775__B2 _6284_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3909_ _6127_/Q _4418_/C _3907_/X vssd1 vssd1 vccd1 vccd1 _3909_/Y sky130_fd_sc_hd__o21ai_4
X_4889_ _6462_/Q _4963_/B _4887_/X _5109_/A1 vssd1 vssd1 vccd1 vccd1 _4889_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3742__A _6284_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_2_1__f_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xci2406_z80_209 vssd1 vssd1 vccd1 vccd1 ci2406_z80_209/HI io_oeb[34] sky130_fd_sc_hd__conb_1
XFILLER_0_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5452__A1 _4863_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5669__A _5732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5204__B2 _6335_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3766__A1 _5268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3917__A _6285_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4512__S _4518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5851__B _6463_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5930_ _5929_/X _5924_/Y _5976_/S vssd1 vssd1 vccd1 vccd1 _5930_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_18_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5861_ _5860_/X _6367_/Q _5861_/S vssd1 vssd1 vccd1 vccd1 _5861_/X sky130_fd_sc_hd__mux2_1
X_5792_ _5792_/A _5792_/B vssd1 vssd1 vccd1 vccd1 _5793_/B sky130_fd_sc_hd__or2_1
X_4812_ _6413_/Q _4793_/Y _4799_/X _4811_/X vssd1 vssd1 vccd1 vccd1 _4812_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_28_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4743_ _6312_/Q _4719_/A _4742_/X _4957_/S vssd1 vssd1 vccd1 vccd1 _4743_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4930__B _4930_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4674_ _5146_/C _5777_/B vssd1 vssd1 vccd1 vccd1 _4676_/B sky130_fd_sc_hd__nor2_1
XANTENNA__3509__A1 _4324_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6413_ _6417_/CLK _6413_/D fanout174/X vssd1 vssd1 vccd1 vccd1 _6413_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3625_ _3603_/Y _3620_/X _3665_/A vssd1 vssd1 vccd1 vccd1 _3625_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_3_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6344_ _6446_/CLK _6344_/D fanout184/X vssd1 vssd1 vccd1 vccd1 _6344_/Q sky130_fd_sc_hd__dfrtp_4
X_3556_ _5400_/A _3527_/C _3555_/X vssd1 vssd1 vccd1 vccd1 _6161_/D sky130_fd_sc_hd__a21o_1
XANTENNA__4182__B2 _4441_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4658__A _4658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6275_ _6307_/CLK _6275_/D fanout183/X vssd1 vssd1 vccd1 vccd1 _6275_/Q sky130_fd_sc_hd__dfstp_1
X_5226_ _6381_/Q _5256_/B _5247_/S vssd1 vssd1 vccd1 vccd1 _5226_/X sky130_fd_sc_hd__mux2_1
X_3487_ _3488_/A _3487_/B vssd1 vssd1 vccd1 vccd1 _3492_/B sky130_fd_sc_hd__and2b_1
XANTENNA__3281__B _5398_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5157_ _5156_/X _6474_/Q _5289_/S vssd1 vssd1 vccd1 vccd1 _5157_/X sky130_fd_sc_hd__mux2_1
X_4108_ _6289_/Q _4109_/B vssd1 vssd1 vccd1 vccd1 _4207_/C sky130_fd_sc_hd__or2_1
X_5088_ _5107_/B _5087_/Y _5108_/S vssd1 vssd1 vccd1 vccd1 _5088_/X sky130_fd_sc_hd__o21a_1
XANTENNA__5434__B2 _5415_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4237__A2 _4406_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4039_ _4438_/A _5303_/B _4030_/Y vssd1 vssd1 vccd1 vccd1 _4039_/X sky130_fd_sc_hd__a21o_1
XANTENNA__3445__B1 _3673_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5428__S _5478_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5833__A1_N _5977_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3472__A _3530_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5425__A1 _5489_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4507__S _4509_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4228__A2 _4227_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3436__B1 _3489_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xmax_cap62 _4794_/Y vssd1 vssd1 vccd1 vccd1 _5104_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_85_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3366__B _5605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6023__A _6023_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold308 _4308_/X vssd1 vssd1 vccd1 vccd1 _6123_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5361__B1 hold604/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3410_ _3557_/B _4344_/A vssd1 vssd1 vccd1 vccd1 _3410_/Y sky130_fd_sc_hd__nand2_1
Xhold319 _4705_/X vssd1 vssd1 vccd1 vccd1 _6306_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4390_ hold109/X _3911_/X _4397_/S vssd1 vssd1 vccd1 vccd1 _4390_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_40_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3341_ _3288_/X _3291_/X _3340_/Y _4263_/A vssd1 vssd1 vccd1 vccd1 _3341_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_0_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3911__B2 _4441_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4197__B _6385_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3272_ _5327_/B _3272_/B _5327_/C _3272_/D vssd1 vssd1 vccd1 vccd1 _3273_/C sky130_fd_sc_hd__and4_1
XANTENNA__5664__A1 _5757_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6060_ _4366_/A _6058_/X _6059_/Y hold442/X _6040_/Y vssd1 vssd1 vccd1 vccd1 _6060_/X
+ sky130_fd_sc_hd__o32a_1
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5011_ _6404_/Q _5010_/X _5971_/S vssd1 vssd1 vccd1 vccd1 _5011_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4417__S _4464_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5102__A _5102_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5913_ _5914_/B _5914_/C _5914_/A vssd1 vssd1 vccd1 vccd1 _5915_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__4941__A _4949_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5844_ _6365_/Q _5863_/S _5843_/X vssd1 vssd1 vccd1 vccd1 _5844_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_29_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4660__B _4668_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5775_ _6430_/Q _5773_/X _5774_/X vssd1 vssd1 vccd1 vccd1 _5775_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_44_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4726_ hold361/X _4303_/A _4768_/S vssd1 vssd1 vccd1 vccd1 _4726_/X sky130_fd_sc_hd__mux2_1
X_4657_ _4782_/A _4652_/X _4654_/Y _4656_/X vssd1 vssd1 vccd1 vccd1 _6294_/D sky130_fd_sc_hd__o22a_1
XFILLER_0_71_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3276__B _4324_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3608_ _3608_/A _3608_/B vssd1 vssd1 vccd1 vccd1 _4804_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_31_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4588_ _4588_/A _4588_/B vssd1 vssd1 vccd1 vccd1 _4588_/X sky130_fd_sc_hd__or2_1
X_6327_ _6426_/CLK _6327_/D fanout171/X vssd1 vssd1 vccd1 vccd1 _6327_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_0_101_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3539_ _5522_/A _3536_/X _3538_/Y vssd1 vssd1 vccd1 vccd1 _3539_/Y sky130_fd_sc_hd__a21oi_1
X_6258_ _6441_/CLK hold50/X fanout181/X vssd1 vssd1 vccd1 vccd1 hold49/A sky130_fd_sc_hd__dfrtp_1
X_5209_ _5279_/C _5209_/B vssd1 vssd1 vccd1 vccd1 _5215_/A sky130_fd_sc_hd__nand2_1
X_6189_ _6472_/CLK hold82/X vssd1 vssd1 vccd1 vccd1 hold81/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__6374__RESET_B fanout172/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6303__RESET_B fanout185/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4835__B _4835_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold601_A _6366_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5018__S0 _5100_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4997__S _5016_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3914__B _6379_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3890_ _3880_/B _4401_/B _3878_/X vssd1 vssd1 vccd1 vccd1 _4425_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__3377__A _5777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5560_ _5594_/A _5561_/B vssd1 vssd1 vccd1 vccd1 _5562_/A sky130_fd_sc_hd__and2_1
X_4511_ _3911_/X hold291/X _4518_/S vssd1 vssd1 vccd1 vccd1 _6218_/D sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_38_wb_clk_i clkbuf_leaf_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6480_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_5491_ _6481_/Q _4920_/B _5593_/S vssd1 vssd1 vccd1 vccd1 _5492_/C sky130_fd_sc_hd__mux2_1
XFILLER_0_80_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold105 _6156_/Q vssd1 vssd1 vccd1 vccd1 hold105/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold116 _6157_/Q vssd1 vssd1 vccd1 vccd1 hold116/X sky130_fd_sc_hd__dlygate4sd3_1
X_4442_ hold271/X _4441_/X _4464_/S vssd1 vssd1 vccd1 vccd1 _6174_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_79_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold127 _4502_/X vssd1 vssd1 vccd1 vccd1 _6210_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 _6200_/Q vssd1 vssd1 vccd1 vccd1 hold138/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold149 _6226_/Q vssd1 vssd1 vccd1 vccd1 hold149/X sky130_fd_sc_hd__dlygate4sd3_1
X_4373_ hold101/X _4085_/X _4376_/S vssd1 vssd1 vccd1 vccd1 _4373_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3324_ _3674_/A _4338_/B vssd1 vssd1 vccd1 vccd1 _3324_/Y sky130_fd_sc_hd__nor2_1
X_6112_ _6263_/CLK _6112_/D vssd1 vssd1 vccd1 vccd1 _6112_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3255_ _3639_/C _3268_/B vssd1 vssd1 vccd1 vccd1 _3691_/B sky130_fd_sc_hd__or2_4
X_6043_ _6076_/A _6071_/S vssd1 vssd1 vccd1 vccd1 _6043_/Y sky130_fd_sc_hd__nor2_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3186_ _5345_/C _3186_/B _3186_/C _3610_/A vssd1 vssd1 vccd1 vccd1 _3187_/D sky130_fd_sc_hd__or4_1
XFILLER_0_14_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout172_A fanout175/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5767__A _5767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4612__A2 _4611_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3820__B1 _3807_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3287__A _4276_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5827_ _5839_/B _5827_/B vssd1 vssd1 vccd1 vccd1 _5827_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5758_ _6309_/Q hold361/X _5765_/S vssd1 vssd1 vccd1 vccd1 _5758_/X sky130_fd_sc_hd__mux2_1
X_4709_ _4713_/A _4708_/X _4714_/S vssd1 vssd1 vccd1 vccd1 _4709_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_32_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5689_ hold442/X _5629_/X _5646_/X hold379/X vssd1 vssd1 vccd1 vccd1 _5700_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_8_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5876__A1 _6368_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold661 _6248_/Q vssd1 vssd1 vccd1 vccd1 hold661/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold650 _6291_/Q vssd1 vssd1 vccd1 vccd1 hold650/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3887__B1 _3852_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4836__C1 _5771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5723__S1 _5734_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4284__C _4605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4851__A2 _4963_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6053__B2 _6036_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6053__A1 _6101_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4603__A2 _4641_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4367__A1 _5769_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4520__S _4527_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4748__A2_N _4720_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6044__A1 _5384_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4991_ _5109_/A1 _4986_/X _4990_/Y _4924_/C vssd1 vssd1 vccd1 vccd1 _4991_/X sky130_fd_sc_hd__a22o_1
X_3942_ _3734_/X _6081_/A _3700_/Y vssd1 vssd1 vccd1 vccd1 _3942_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_73_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3873_ _3714_/S _3717_/B _3726_/Y _3727_/Y _6187_/Q vssd1 vssd1 vccd1 vccd1 _3873_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_0_45_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5612_ _5645_/A _5645_/B vssd1 vssd1 vccd1 vccd1 _5653_/A sky130_fd_sc_hd__nor2_1
X_5543_ _5543_/A _5543_/B vssd1 vssd1 vccd1 vccd1 _5545_/B sky130_fd_sc_hd__and2_1
XFILLER_0_26_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_15_wb_clk_i_A _6448_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5474_ _5472_/X _5473_/X _5567_/B vssd1 vssd1 vccd1 vccd1 _5474_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5858__A1 _5786_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5858__B2 _5887_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4425_ _4425_/A _4425_/B vssd1 vssd1 vccd1 vccd1 _4425_/Y sky130_fd_sc_hd__nand2_1
X_4356_ hold332/X _4355_/X _5769_/S vssd1 vssd1 vccd1 vccd1 _4356_/X sky130_fd_sc_hd__mux2_1
X_3307_ _3307_/A _3307_/B vssd1 vssd1 vccd1 vccd1 _3308_/B sky130_fd_sc_hd__nand2_2
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4666__A input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3570__A _5605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4287_ hold5/X _4286_/X _5769_/S vssd1 vssd1 vccd1 vccd1 hold6/A sky130_fd_sc_hd__mux2_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3238_ _3627_/B _3627_/C vssd1 vssd1 vccd1 vccd1 _3632_/D sky130_fd_sc_hd__nor2_4
X_6026_ _6025_/X _3594_/A _6026_/S vssd1 vssd1 vccd1 vccd1 _6467_/D sky130_fd_sc_hd__mux2_1
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4294__B1 _6309_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3169_ _5387_/A _4557_/C _4557_/D vssd1 vssd1 vccd1 vccd1 _4556_/C sky130_fd_sc_hd__nor3_4
XFILLER_0_49_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout88 _4360_/Y vssd1 vssd1 vccd1 vccd1 _5817_/A sky130_fd_sc_hd__buf_4
Xfanout99 _4791_/Y vssd1 vssd1 vccd1 vccd1 _5892_/S sky130_fd_sc_hd__clkbuf_8
Xfanout77 _5901_/B vssd1 vssd1 vccd1 vccd1 _5970_/A sky130_fd_sc_hd__buf_4
Xfanout66 _4789_/Y vssd1 vssd1 vccd1 vccd1 _5842_/B1 sky130_fd_sc_hd__buf_2
XFILLER_0_51_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5436__S _5499_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold480 _5999_/X vssd1 vssd1 vccd1 vccd1 _6435_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold491 _6436_/Q vssd1 vssd1 vccd1 vccd1 hold491/X sky130_fd_sc_hd__buf_1
XFILLER_0_87_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5785__B1 _5977_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4515__S _4518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3260__A1 _3172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3639__B _5322_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3655__A _6023_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4210_ _4210_/A _4210_/B vssd1 vssd1 vccd1 vccd1 _4212_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_50_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5190_ _5267_/C _5267_/D vssd1 vssd1 vccd1 vccd1 _5192_/A sky130_fd_sc_hd__xor2_1
X_4141_ _6157_/Q _3799_/X _3801_/X _6148_/Q _4140_/X vssd1 vssd1 vccd1 vccd1 _4144_/A
+ sky130_fd_sc_hd__a221o_1
X_4072_ _4073_/A _3759_/Y _4115_/A _5262_/C _3979_/A vssd1 vssd1 vccd1 vccd1 _4072_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4815__A2 _5771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4579__B2 _6159_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4974_ _5521_/A _5861_/S _5842_/B1 _4973_/X vssd1 vssd1 vccd1 vccd1 _4974_/X sky130_fd_sc_hd__a22o_1
X_3925_ _6379_/Q _6383_/Q _6343_/Q vssd1 vssd1 vccd1 vccd1 _5267_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_86_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3549__B _5388_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5528__B1 _4300_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout135_A _4313_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3856_ _3816_/B _3855_/X _3852_/X vssd1 vssd1 vccd1 vccd1 _3859_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_81_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3787_ _3557_/B _3786_/Y _5522_/A vssd1 vssd1 vccd1 vccd1 _3787_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_61_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5526_ _6101_/A _5485_/S _5519_/Y _5521_/Y _5598_/S vssd1 vssd1 vccd1 vccd1 _5526_/X
+ sky130_fd_sc_hd__o311a_1
XANTENNA__3284__B _3284_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5457_ _5457_/A _5457_/B vssd1 vssd1 vccd1 vccd1 _5457_/X sky130_fd_sc_hd__xor2_1
X_4408_ _6211_/Q _6203_/Q _4408_/S vssd1 vssd1 vccd1 vccd1 _4408_/X sky130_fd_sc_hd__mux2_1
X_5388_ _5388_/A _5388_/B _5388_/C _5387_/X vssd1 vssd1 vccd1 vccd1 _5388_/X sky130_fd_sc_hd__or4b_1
X_4339_ _4782_/A _5314_/S _4338_/X _4325_/C vssd1 vssd1 vccd1 vccd1 _4339_/X sky130_fd_sc_hd__a31o_1
XANTENNA__3711__C1 _5478_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6009_ _4448_/X hold246/X _6011_/S vssd1 vssd1 vccd1 vccd1 _6454_/D sky130_fd_sc_hd__mux2_1
XANTENNA__4019__A0 _6286_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3490__A1 _3530_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4990__A1 _5427_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3475__A _5995_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3194__B _3205_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5298__A2 _5299_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5758__A0 _6309_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3710_ _3695_/Y _3717_/A _3709_/X _5384_/A vssd1 vssd1 vccd1 vccd1 _4546_/A sky130_fd_sc_hd__a31o_4
XFILLER_0_7_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4690_ _4715_/B2 _4688_/Y _4689_/X hold326/X _4672_/Y vssd1 vssd1 vccd1 vccd1 _4690_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_0_43_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3641_ hold298/X _3648_/C _3648_/B vssd1 vssd1 vccd1 vccd1 _3641_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_43_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5076__S _6070_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3536__A2 _5617_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3572_ _5314_/S _3412_/B _4325_/C vssd1 vssd1 vccd1 vccd1 _3572_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__3385__A _4324_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6360_ _6377_/CLK _6360_/D vssd1 vssd1 vccd1 vccd1 _6360_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3816__C _3885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5311_ _5311_/A _5311_/B _5311_/C _5311_/D vssd1 vssd1 vccd1 vccd1 _5311_/X sky130_fd_sc_hd__or4_1
XFILLER_0_3_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6291_ _6441_/CLK _6291_/D vssd1 vssd1 vccd1 vccd1 _6291_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5242_ hold610/X _5241_/X _5489_/S vssd1 vssd1 vccd1 vccd1 _6337_/D sky130_fd_sc_hd__mux2_1
X_5173_ _5174_/A _5173_/B vssd1 vssd1 vccd1 vccd1 _5261_/B sky130_fd_sc_hd__nand2_1
XANTENNA__5694__C1 _5730_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4124_ _6264_/Q _3793_/X _3795_/X _6199_/Q vssd1 vssd1 vccd1 vccd1 _4124_/X sky130_fd_sc_hd__a22o_1
Xinput1 custom_settings[0] vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__clkbuf_2
X_4055_ _6334_/Q _3933_/Y _4107_/C _4054_/Y vssd1 vssd1 vccd1 vccd1 _4056_/B sky130_fd_sc_hd__o22a_1
XANTENNA__5997__B1 _4363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4421__B1 _4408_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4957_ hold274/X _4956_/X _4957_/S vssd1 vssd1 vccd1 vccd1 _4957_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_74_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3908_ _6127_/Q _4418_/C _3907_/X vssd1 vssd1 vccd1 vccd1 _3908_/X sky130_fd_sc_hd__o21a_1
XANTENNA__4972__A1 _6421_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4888_ _6479_/Q _5104_/A2 _4796_/Y _4881_/X _4793_/Y vssd1 vssd1 vccd1 vccd1 _4888_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_61_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3839_ _4052_/A _3839_/B vssd1 vssd1 vccd1 vccd1 _4444_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__5921__B1 _5784_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5509_ hold592/X _5520_/B _5508_/Y _5485_/S vssd1 vssd1 vccd1 vccd1 _5509_/Y sky130_fd_sc_hd__o2bb2ai_1
X_6489_ _6489_/CLK _6489_/D fanout176/X vssd1 vssd1 vccd1 vccd1 _6489_/Q sky130_fd_sc_hd__dfstp_2
XANTENNA__4838__B _5783_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4557__C _4557_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold631_A _6313_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4292__C _5418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3518__A2 _5314_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4715__B2 _4715_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6489__SET_B fanout176/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5851__C _5866_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5140__A1 _5605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5691__A2 _5721_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4651__B1 _5567_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5860_ _6419_/Q _4791_/Y _4921_/X vssd1 vssd1 vccd1 vccd1 _5860_/X sky130_fd_sc_hd__a21o_1
X_4811_ _4924_/C _4809_/Y _4810_/X _4801_/X _5109_/A1 vssd1 vssd1 vccd1 vccd1 _4811_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_68_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5791_ _5792_/A _5792_/B vssd1 vssd1 vccd1 vccd1 _5804_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_7_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4703__S _4712_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4742_ _6312_/Q _4720_/X _5224_/A2 hold476/X vssd1 vssd1 vccd1 vccd1 _4742_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_56_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4954__A1 _6368_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4673_ _6076_/A _4714_/S vssd1 vssd1 vccd1 vccd1 _4673_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_71_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3624_ _3665_/A _5757_/A vssd1 vssd1 vccd1 vccd1 _3624_/Y sky130_fd_sc_hd__nand2_1
X_6412_ _6412_/CLK hold20/X vssd1 vssd1 vccd1 vccd1 hold19/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4004__A _6287_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6343_ _6446_/CLK _6343_/D fanout184/X vssd1 vssd1 vccd1 vccd1 _6343_/Q sky130_fd_sc_hd__dfrtp_4
X_3555_ _4363_/A _5400_/A _5600_/C _5400_/B _4324_/B vssd1 vssd1 vccd1 vccd1 _3555_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_3_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3486_ _3480_/B _3481_/B _3492_/A hold432/X vssd1 vssd1 vccd1 vccd1 _3486_/X sky130_fd_sc_hd__a211o_1
X_6274_ _6336_/CLK _6274_/D fanout182/X vssd1 vssd1 vccd1 vccd1 _6274_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA__4658__B _4668_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3562__B _3619_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5225_ _6336_/Q _5131_/Y _5224_/X _5016_/S _5151_/B vssd1 vssd1 vccd1 vccd1 _5225_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5667__C1 _5730_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5682__A2 _5721_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5156_ _6335_/Q _6277_/Q _5288_/S vssd1 vssd1 vccd1 vccd1 _5156_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_98_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4107_ _6288_/Q _4107_/B _4107_/C vssd1 vssd1 vccd1 vccd1 _4109_/B sky130_fd_sc_hd__or3_1
X_5087_ _6374_/Q _5086_/C _6375_/Q vssd1 vssd1 vccd1 vccd1 _5087_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_79_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5434__A2 _5520_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4038_ _4038_/A _4038_/B vssd1 vssd1 vccd1 vccd1 _5303_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_2_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5198__B2 _6381_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5198__A1 _6384_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5989_ _4335_/B _5978_/Y _5980_/Y _5988_/X vssd1 vssd1 vccd1 vccd1 _5989_/X sky130_fd_sc_hd__a22o_1
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3381__B1 _3673_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3532__A_N _5617_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5189__A1 _5866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4523__S _4527_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold309 _6220_/Q vssd1 vssd1 vccd1 vccd1 hold309/X sky130_fd_sc_hd__dlygate4sd3_1
X_3340_ _4264_/B _3673_/B _3424_/B vssd1 vssd1 vccd1 vccd1 _3340_/Y sky130_fd_sc_hd__a21oi_1
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3271_ _3163_/A _3161_/B _3222_/X vssd1 vssd1 vccd1 vccd1 _3272_/D sky130_fd_sc_hd__a21o_1
X_5010_ _6423_/Q _4793_/Y _5004_/X _5009_/X vssd1 vssd1 vccd1 vccd1 _5010_/X sky130_fd_sc_hd__a211o_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3675__B2 _3674_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5912_ _5912_/A _5912_/B vssd1 vssd1 vccd1 vccd1 _5914_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_75_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5843_ _5817_/A _5842_/X _4882_/X vssd1 vssd1 vccd1 vccd1 _5843_/X sky130_fd_sc_hd__a21o_1
XANTENNA__5529__S _5593_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4927__B2 _4920_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5774_ _5774_/A _5774_/B _5774_/C _3379_/B vssd1 vssd1 vccd1 vccd1 _5774_/X sky130_fd_sc_hd__or4b_1
XFILLER_0_44_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4725_ _6033_/A _4725_/B vssd1 vssd1 vccd1 vccd1 _4770_/S sky130_fd_sc_hd__nand2_4
XFILLER_0_44_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4656_ _4656_/A _4668_/B vssd1 vssd1 vccd1 vccd1 _4656_/X sky130_fd_sc_hd__and2_1
X_3607_ _3110_/A _3281_/A _3300_/B _5371_/C _5369_/A vssd1 vssd1 vccd1 vccd1 _3608_/B
+ sky130_fd_sc_hd__a2111o_1
X_4587_ _4359_/B _3547_/X _3322_/C vssd1 vssd1 vccd1 vccd1 _4588_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_101_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3538_ _5317_/A _3352_/B _5146_/C vssd1 vssd1 vccd1 vccd1 _3538_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_12_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6326_ _6419_/CLK _6326_/D fanout173/X vssd1 vssd1 vccd1 vccd1 _6326_/Q sky130_fd_sc_hd__dfrtp_1
X_6257_ _6441_/CLK _6257_/D fanout181/X vssd1 vssd1 vccd1 vccd1 _6257_/Q sky130_fd_sc_hd__dfrtp_1
X_3469_ _3469_/A _3469_/B vssd1 vssd1 vccd1 vccd1 _3636_/B sky130_fd_sc_hd__nand2_4
X_5208_ _6463_/Q _6462_/Q vssd1 vssd1 vccd1 vccd1 _5209_/B sky130_fd_sc_hd__nand2_1
X_6188_ _6449_/CLK _6188_/D vssd1 vssd1 vccd1 vccd1 _6188_/Q sky130_fd_sc_hd__dfxtp_1
X_5139_ _6343_/Q _4150_/A _6333_/Q _6346_/Q vssd1 vssd1 vccd1 vccd1 _5139_/X sky130_fd_sc_hd__o211a_1
XANTENNA__3418__A1 _3284_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_8_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6444_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_39_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_hold427_A _6330_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3467__B _3501_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5018__S1 _5100_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5343__A1 _5364_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4777__S0 _5078_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4518__S _4518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5582__A1 _6101_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4510_ _4546_/A _6003_/A vssd1 vssd1 vccd1 vccd1 _4518_/S sky130_fd_sc_hd__or2_4
X_5490_ _5757_/A _6464_/Q vssd1 vssd1 vccd1 vccd1 _5492_/B sky130_fd_sc_hd__or2_1
XFILLER_0_79_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold106 _4395_/X vssd1 vssd1 vccd1 vccd1 _6156_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold117 _4396_/X vssd1 vssd1 vccd1 vccd1 _6157_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4441_ _4439_/X _4440_/X _4441_/S vssd1 vssd1 vccd1 vccd1 _4441_/X sky130_fd_sc_hd__mux2_2
Xhold128 _6265_/Q vssd1 vssd1 vccd1 vccd1 hold128/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5084__S _5105_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold139 _6158_/Q vssd1 vssd1 vccd1 vccd1 hold139/X sky130_fd_sc_hd__dlygate4sd3_1
X_4372_ hold174/X _4042_/X _4376_/S vssd1 vssd1 vccd1 vccd1 _4372_/X sky130_fd_sc_hd__mux2_1
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6111_ _6393_/CLK _6111_/D vssd1 vssd1 vccd1 vccd1 _6111_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4001__B _6381_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3323_ _3323_/A _3326_/A _5387_/A vssd1 vssd1 vccd1 vccd1 _4253_/A sky130_fd_sc_hd__or3_4
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3254_ _3273_/A _3273_/B vssd1 vssd1 vccd1 vccd1 _3254_/Y sky130_fd_sc_hd__nand2_1
X_6042_ _5567_/B _6041_/X _6071_/S vssd1 vssd1 vccd1 vccd1 _6042_/X sky130_fd_sc_hd__o21a_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3185_ _3185_/A _4804_/D vssd1 vssd1 vccd1 vccd1 _3610_/A sky130_fd_sc_hd__nand2_1
XANTENNA_fanout165_A _5600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5217__A1_N _5291_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_44_wb_clk_i_A clkbuf_leaf_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__3568__A _5317_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3287__B _3489_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5826_ _5826_/A _5826_/B _5824_/X vssd1 vssd1 vccd1 vccd1 _5827_/B sky130_fd_sc_hd__or3b_1
XANTENNA__5022__B1 _5021_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5757_ _5757_/A _5757_/B _5757_/C _4724_/C vssd1 vssd1 vccd1 vccd1 _5765_/S sky130_fd_sc_hd__or4b_4
XFILLER_0_44_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4708_ _6286_/Q _4707_/X _4712_/S vssd1 vssd1 vccd1 vccd1 _4708_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5783__A _5783_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5325__A1 _4675_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5688_ _5757_/B _4027_/A _5611_/Y _5687_/X vssd1 vssd1 vccd1 vccd1 _5688_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_44_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4639_ hold440/X _4604_/X _4605_/X _6489_/Q _4638_/X vssd1 vssd1 vccd1 vccd1 _4639_/X
+ sky130_fd_sc_hd__a221o_1
Xhold651 _4645_/X vssd1 vssd1 vccd1 vccd1 _6291_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold640 _6468_/Q vssd1 vssd1 vccd1 vccd1 _3500_/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3887__A1 _3883_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6309_ _6336_/CLK _6309_/D fanout182/X vssd1 vssd1 vccd1 vccd1 _6309_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__6053__A2 _4863_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4367__A2 _5078_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4801__S _4948_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3941__A _6081_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4055__A1 _6334_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5252__A0 _6097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4990_ _5427_/B _4808_/Y _4989_/X vssd1 vssd1 vccd1 vccd1 _4990_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_58_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3941_ _6081_/A vssd1 vssd1 vccd1 vccd1 _3941_/Y sky130_fd_sc_hd__inv_2
X_3872_ _3723_/Y _3869_/X _3871_/X _3852_/A vssd1 vssd1 vccd1 vccd1 _3878_/B sky130_fd_sc_hd__a211o_1
X_5611_ _5644_/A _5646_/B _4300_/A vssd1 vssd1 vccd1 vccd1 _5611_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__5555__B2 _5415_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4711__S _4711_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5542_ _5594_/A _5542_/B vssd1 vssd1 vccd1 vccd1 _5543_/B sky130_fd_sc_hd__or2_1
XFILLER_0_14_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5473_ hold595/X input6/X _5510_/S vssd1 vssd1 vccd1 vccd1 _5473_/X sky130_fd_sc_hd__mux2_1
X_4424_ _5732_/A _4421_/X _4422_/X _4423_/X vssd1 vssd1 vccd1 vccd1 _4424_/X sky130_fd_sc_hd__o31a_1
X_4355_ _6359_/Q _5601_/A _4355_/S vssd1 vssd1 vccd1 vccd1 _4355_/X sky130_fd_sc_hd__mux2_1
X_3306_ _3307_/A _3307_/B vssd1 vssd1 vccd1 vccd1 _3433_/B sky130_fd_sc_hd__and2_1
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4666__B _4668_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4286_ _6359_/Q _6377_/Q _4286_/S vssd1 vssd1 vccd1 vccd1 _4286_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4818__B1 _4789_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3237_ _4273_/A _6300_/Q _6299_/Q _4268_/A vssd1 vssd1 vccd1 vccd1 _3627_/C sky130_fd_sc_hd__or4b_4
X_6025_ _6025_/A _6025_/B vssd1 vssd1 vccd1 vccd1 _6025_/X sky130_fd_sc_hd__or2_1
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4294__B2 _4322_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3168_ _4782_/A _3168_/B _4782_/B _3547_/B vssd1 vssd1 vccd1 vccd1 _4557_/D sky130_fd_sc_hd__or4b_4
XANTENNA_clkbuf_leaf_0_wb_clk_i_A clkbuf_leaf_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_55_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3099_ _3099_/A vssd1 vssd1 vccd1 vccd1 _6446_/D sky130_fd_sc_hd__inv_2
XFILLER_0_89_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5243__A0 _6338_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xci2406_z80_190 vssd1 vssd1 vccd1 vccd1 ci2406_z80_190/HI io_oeb[5] sky130_fd_sc_hd__conb_1
XANTENNA__5794__B2 _5976_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5794__A1 _5786_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout78 _4776_/Y vssd1 vssd1 vccd1 vccd1 _5771_/A sky130_fd_sc_hd__buf_4
Xfanout89 _4418_/C vssd1 vssd1 vccd1 vccd1 _4441_/S sky130_fd_sc_hd__buf_6
X_5809_ _6415_/Q _5867_/B _5809_/C vssd1 vssd1 vccd1 vccd1 _5826_/A sky130_fd_sc_hd__and3_1
XANTENNA__5546__B2 _5415_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout67 _5861_/S vssd1 vssd1 vccd1 vccd1 _5848_/S sky130_fd_sc_hd__buf_4
XFILLER_0_17_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4621__S _4641_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3745__B _6333_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold470 _6287_/Q vssd1 vssd1 vccd1 vccd1 hold470/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold481 _6281_/Q vssd1 vssd1 vccd1 vccd1 hold481/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold492 _3653_/X vssd1 vssd1 vccd1 vccd1 _6436_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5452__S _5593_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5785__A1 _6023_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4531__S _4536_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6446__RESET_B fanout185/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4140_ _6265_/Q _3793_/X _3795_/X _6200_/Q vssd1 vssd1 vccd1 vccd1 _4140_/X sky130_fd_sc_hd__a22o_1
X_4071_ _5161_/A vssd1 vssd1 vccd1 vccd1 _5257_/A sky130_fd_sc_hd__inv_2
XANTENNA__5776__B2 _5387_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4973_ _6402_/Q _4972_/X _5892_/S vssd1 vssd1 vccd1 vccd1 _4973_/X sky130_fd_sc_hd__mux2_1
X_3924_ _5136_/A _6285_/Q _6379_/Q _4060_/B _3923_/X vssd1 vssd1 vccd1 vccd1 _5162_/B
+ sky130_fd_sc_hd__o41a_2
XANTENNA__3549__C _4248_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5537__S _5581_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4441__S _4441_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3855_ _3853_/X _3854_/X _3883_/S vssd1 vssd1 vccd1 vccd1 _3855_/X sky130_fd_sc_hd__mux2_1
X_3786_ _3786_/A _4786_/C vssd1 vssd1 vccd1 vccd1 _3786_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_73_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout128_A hold526/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_22_wb_clk_i _6448_/CLK vssd1 vssd1 vccd1 vccd1 _6336_/CLK sky130_fd_sc_hd__clkbuf_16
X_5525_ _5593_/S _5525_/B vssd1 vssd1 vccd1 vccd1 _5598_/S sky130_fd_sc_hd__nand2_4
XFILLER_0_74_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5456_ _5445_/A _5445_/B _5443_/A vssd1 vssd1 vccd1 vccd1 _5457_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_41_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4407_ _6187_/Q _4408_/S _5731_/C1 _4406_/X vssd1 vssd1 vccd1 vccd1 _4407_/X sky130_fd_sc_hd__o211a_1
X_5387_ _5387_/A _5387_/B _5387_/C vssd1 vssd1 vccd1 vccd1 _5387_/X sky130_fd_sc_hd__or3_1
X_4338_ _4338_/A _4338_/B vssd1 vssd1 vccd1 vccd1 _4338_/X sky130_fd_sc_hd__or2_1
XFILLER_0_5_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4269_ _5522_/D _4268_/Y _4267_/Y vssd1 vssd1 vccd1 vccd1 _4269_/X sky130_fd_sc_hd__o21a_1
X_6008_ _4441_/X hold296/X _6011_/S vssd1 vssd1 vccd1 vccd1 _6453_/D sky130_fd_sc_hd__mux2_1
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5216__B1 _5291_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4616__S _4641_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3475__B _4363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4258__A1 _4782_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5211__A _6465_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4526__S _4527_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3640_ _3640_/A _6446_/Q _3640_/C vssd1 vssd1 vccd1 vccd1 _3648_/C sky130_fd_sc_hd__and3_1
X_3571_ _4344_/A _5617_/A _4344_/B _3569_/X vssd1 vssd1 vccd1 vccd1 _3571_/X sky130_fd_sc_hd__a31o_1
X_5310_ _5369_/A _5369_/D _5346_/B _5310_/D vssd1 vssd1 vccd1 vccd1 _5311_/D sky130_fd_sc_hd__or4_1
X_6290_ _6441_/CLK _6290_/D vssd1 vssd1 vccd1 vccd1 _6290_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_51_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5241_ _6093_/A _5292_/S _5147_/X _5240_/X vssd1 vssd1 vccd1 vccd1 _5241_/X sky130_fd_sc_hd__a2bb2o_1
XANTENNA__4041__S0 _5721_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5172_ _5172_/A _5172_/B vssd1 vssd1 vccd1 vccd1 _5177_/A sky130_fd_sc_hd__xnor2_1
X_4123_ _4438_/A _6097_/A _4462_/A2 vssd1 vssd1 vccd1 vccd1 _4123_/Y sky130_fd_sc_hd__o21ai_1
X_4054_ _6334_/Q _6337_/Q vssd1 vssd1 vccd1 vccd1 _4054_/Y sky130_fd_sc_hd__nand2_1
Xinput2 custom_settings[1] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__buf_1
XFILLER_0_78_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4436__S _4464_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4956_ _6368_/Q _4955_/X _5974_/S vssd1 vssd1 vccd1 vccd1 _4956_/X sky130_fd_sc_hd__mux2_1
X_3907_ _6377_/Q _4463_/S vssd1 vssd1 vccd1 vccd1 _3907_/X sky130_fd_sc_hd__or2_1
X_4887_ _4881_/X _4886_/X _4948_/S vssd1 vssd1 vccd1 vccd1 _4887_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_34_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3838_ _3838_/A _3838_/B _3838_/C vssd1 vssd1 vccd1 vccd1 _3839_/B sky130_fd_sc_hd__or3_2
XFILLER_0_61_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4185__B1 _3801_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3932__B1 _6287_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3769_ _3772_/B _4156_/A _6346_/Q vssd1 vssd1 vccd1 vccd1 _3770_/A sky130_fd_sc_hd__and3b_4
XANTENNA__6368__RESET_B fanout181/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5508_ _5508_/A _5508_/B vssd1 vssd1 vccd1 vccd1 _5508_/Y sky130_fd_sc_hd__xnor2_2
X_6488_ _6488_/CLK _6488_/D fanout172/X vssd1 vssd1 vccd1 vccd1 _6488_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_0_100_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5439_ _5757_/A _6460_/Q vssd1 vssd1 vccd1 vccd1 _5441_/B sky130_fd_sc_hd__or2_1
XANTENNA__5685__B1 _5684_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5437__A0 _6459_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout60_A _5975_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold624_A _6461_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4412__A1 _5732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5140__A2 _5268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3652__C _5388_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6037__A _6070_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4651__A1 _5995_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4810_ _6361_/Q _5108_/S vssd1 vssd1 vccd1 vccd1 _4810_/X sky130_fd_sc_hd__or2_1
XFILLER_0_68_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5790_ _5866_/A _5411_/B _5866_/C _5867_/B vssd1 vssd1 vccd1 vccd1 _5792_/B sky130_fd_sc_hd__o31ai_1
XFILLER_0_90_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3396__A _5388_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4741_ hold635/X _4740_/X _5232_/S vssd1 vssd1 vccd1 vccd1 _6311_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_83_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4672_ _4713_/A _4714_/S _4715_/B2 vssd1 vssd1 vccd1 vccd1 _4672_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_0_28_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3623_ _3621_/X _3622_/Y _3665_/A vssd1 vssd1 vccd1 vccd1 _6169_/D sky130_fd_sc_hd__mux2_1
X_6411_ _6472_/CLK hold42/X vssd1 vssd1 vccd1 vccd1 hold41/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__6461__RESET_B fanout181/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6342_ _6441_/CLK _6342_/D fanout184/X vssd1 vssd1 vccd1 vccd1 _6342_/Q sky130_fd_sc_hd__dfrtp_1
X_3554_ _3554_/A _5400_/B vssd1 vssd1 vccd1 vccd1 _3554_/X sky130_fd_sc_hd__and2_1
XFILLER_0_3_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3485_ _5995_/C _3487_/B _3484_/X _3472_/B _3477_/X vssd1 vssd1 vccd1 vccd1 _3485_/X
+ sky130_fd_sc_hd__a221o_1
X_6273_ _6312_/CLK _6273_/D fanout182/X vssd1 vssd1 vccd1 vccd1 _6273_/Q sky130_fd_sc_hd__dfstp_1
X_5224_ _6278_/Q _5224_/A2 _5123_/Y _5223_/X vssd1 vssd1 vccd1 vccd1 _5224_/X sky130_fd_sc_hd__a22o_1
X_5155_ hold645/X _5154_/X _5232_/S vssd1 vssd1 vccd1 vccd1 _6334_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_47_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5550__S _5593_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4106_ _4106_/A _4205_/S vssd1 vssd1 vccd1 vccd1 _4162_/A sky130_fd_sc_hd__or2_1
XANTENNA__4674__B _5777_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5086_ _6374_/Q _6375_/Q _5086_/C vssd1 vssd1 vccd1 vccd1 _5107_/B sky130_fd_sc_hd__and3_1
XANTENNA__6092__B1 _6107_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4037_ _4190_/A _3962_/B _3967_/A vssd1 vssd1 vccd1 vccd1 _4038_/B sky130_fd_sc_hd__a21o_1
XANTENNA__3445__A2 _3685_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5198__A2 _4332_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5988_ _6437_/Q _5988_/B vssd1 vssd1 vccd1 vccd1 _5988_/X sky130_fd_sc_hd__and2b_1
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4939_ _6209_/Q _6217_/Q _6456_/Q _6233_/Q _5404_/A0 _5078_/S1 vssd1 vssd1 vccd1
+ vccd1 _4939_/X sky130_fd_sc_hd__mux4_2
XFILLER_0_74_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3905__B1 _4463_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6131__RESET_B fanout180/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3381__A1 _6431_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4330__B1 _5362_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4865__A _6364_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5189__A2 _6335_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3663__B _5478_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3270_ _3229_/A _3057_/Y _3219_/Y _3264_/X _3685_/A vssd1 vssd1 vccd1 vccd1 _5327_/C
+ sky130_fd_sc_hd__o311a_1
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4321__B1 _4322_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3675__A2 _3673_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6074__B1 _6101_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_34_wb_clk_i_A clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_5911_ _6421_/Q _6422_/Q _5901_/B vssd1 vssd1 vccd1 vccd1 _5914_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_48_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4714__S _4714_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5842_ _6365_/Q _5861_/S _5842_/B1 _5841_/X vssd1 vssd1 vccd1 vccd1 _5842_/X sky130_fd_sc_hd__a22o_1
X_5773_ _4248_/B _4248_/C _3308_/B _3396_/B _4335_/C vssd1 vssd1 vccd1 vccd1 _5773_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_90_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4724_ _5605_/B _6469_/Q _4724_/C vssd1 vssd1 vccd1 vccd1 _5289_/S sky130_fd_sc_hd__and3_4
XFILLER_0_8_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4655_ _3168_/B _4652_/X _4654_/Y _4650_/X vssd1 vssd1 vccd1 vccd1 _6293_/D sky130_fd_sc_hd__o22a_1
XANTENNA__5337__C1 _3632_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3606_ _3282_/A _3180_/B _3253_/A _5522_/B vssd1 vssd1 vccd1 vccd1 _4806_/A sky130_fd_sc_hd__o211a_1
X_4586_ _4267_/Y _4583_/X _4585_/Y _5774_/A _5388_/A vssd1 vssd1 vccd1 vccd1 _4586_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_71_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3537_ _5315_/B _5388_/A _5314_/S vssd1 vssd1 vccd1 vccd1 _3574_/B sky130_fd_sc_hd__or3_1
X_6325_ _6407_/CLK _6325_/D fanout170/X vssd1 vssd1 vccd1 vccd1 _6325_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3468_ _6021_/S _3594_/B vssd1 vssd1 vccd1 vccd1 _3469_/B sky130_fd_sc_hd__nor2_1
X_6256_ _6456_/CLK _6256_/D vssd1 vssd1 vccd1 vccd1 _6256_/Q sky130_fd_sc_hd__dfxtp_1
X_3399_ _5369_/C _3399_/B _5372_/A _5311_/A vssd1 vssd1 vccd1 vccd1 _3399_/X sky130_fd_sc_hd__or4_2
XANTENNA__5280__S _5291_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5207_ _6463_/Q _6462_/Q vssd1 vssd1 vccd1 vccd1 _5279_/C sky130_fd_sc_hd__or2_1
X_6187_ _6412_/CLK _6187_/D vssd1 vssd1 vccd1 vccd1 _6187_/Q sky130_fd_sc_hd__dfxtp_1
X_5138_ _5233_/B _5137_/Y _5138_/S vssd1 vssd1 vccd1 vccd1 _5138_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_79_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5069_ _6463_/Q _5068_/X _5108_/S vssd1 vssd1 vccd1 vccd1 _5069_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_47_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4777__S1 _5404_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4534__S _4536_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5031__A1 _6424_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3674__A _3674_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold107 _6184_/Q vssd1 vssd1 vccd1 vccd1 hold107/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4440_ hold249/X hold211/X hold197/X hold85/X _5721_/C1 _5721_/B1 vssd1 vssd1 vccd1
+ vccd1 _4440_/X sky130_fd_sc_hd__mux4_2
XANTENNA__3345__A1 _3304_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold118 _6173_/Q vssd1 vssd1 vccd1 vccd1 hold118/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold129 _4553_/X vssd1 vssd1 vccd1 vccd1 _6265_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4371_ hold257/X _3998_/X _4376_/S vssd1 vssd1 vccd1 vccd1 _6136_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_95_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3322_ _3323_/A _4782_/B _3322_/C vssd1 vssd1 vccd1 vccd1 _4784_/D sky130_fd_sc_hd__and3b_2
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3253_ _3253_/A _3253_/B _3253_/C vssd1 vssd1 vccd1 vccd1 _3273_/B sky130_fd_sc_hd__and3_1
X_6041_ _6101_/B _5413_/B _5414_/Y _6036_/X vssd1 vssd1 vccd1 vccd1 _6041_/X sky130_fd_sc_hd__o22a_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3184_ _5315_/A _5774_/A vssd1 vssd1 vccd1 vccd1 _4804_/D sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_47_wb_clk_i clkbuf_leaf_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6239_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout158_A _4782_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5825_ _5826_/A _5826_/B _5824_/X vssd1 vssd1 vccd1 vccd1 _5839_/B sky130_fd_sc_hd__o21ba_1
XANTENNA__3820__A2 _3804_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5022__A1 _6312_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5756_ hold11/X _4190_/B _6104_/S vssd1 vssd1 vccd1 vccd1 hold12/A sky130_fd_sc_hd__mux2_1
X_4707_ _6384_/Q _6380_/Q _4711_/S vssd1 vssd1 vccd1 vccd1 _4707_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3584__A1 _3581_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5687_ _5687_/A _5687_/B _5687_/C vssd1 vssd1 vccd1 vccd1 _5687_/X sky130_fd_sc_hd__or3_1
XFILLER_0_71_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4638_ _6464_/Q _4606_/X _4607_/X _6315_/Q _4637_/X vssd1 vssd1 vccd1 vccd1 _4638_/X
+ sky130_fd_sc_hd__a221o_1
Xhold630 _6310_/Q vssd1 vssd1 vccd1 vccd1 hold630/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4569_ hold527/X _6334_/Q _4575_/S vssd1 vssd1 vccd1 vccd1 _4569_/X sky130_fd_sc_hd__mux2_1
Xhold641 _6129_/Q vssd1 vssd1 vccd1 vccd1 hold641/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold652 _6355_/Q vssd1 vssd1 vccd1 vccd1 hold652/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5730__C1 _5730_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6308_ _6308_/CLK _6308_/D fanout185/X vssd1 vssd1 vccd1 vccd1 _6308_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__5089__A1 _6464_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6239_ _6239_/CLK _6239_/D vssd1 vssd1 vccd1 vccd1 _6239_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5958__B _5970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5013__A1 _5102_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4447__S0 _5721_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4772__B1 _3503_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5721__C1 _5721_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4529__S _4536_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5788__C1 _5102_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3940_ _3928_/A _3939_/X _4227_/S vssd1 vssd1 vccd1 vccd1 _6081_/A sky130_fd_sc_hd__mux2_4
XFILLER_0_85_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3871_ hold266/X _3861_/S _3870_/X _3883_/S vssd1 vssd1 vccd1 vccd1 _3871_/X sky130_fd_sc_hd__o211a_1
X_5610_ _5645_/A _5610_/B vssd1 vssd1 vccd1 vccd1 _5646_/B sky130_fd_sc_hd__and2_1
XANTENNA__5555__A2 _5520_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5541_ _5594_/A _5542_/B vssd1 vssd1 vccd1 vccd1 _5543_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_81_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6336__SET_B fanout183/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5472_ _5470_/X _5471_/X _5485_/S vssd1 vssd1 vccd1 vccd1 _5472_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4423_ _5730_/C1 _4420_/X _4419_/X _5655_/B vssd1 vssd1 vccd1 vccd1 _4423_/X sky130_fd_sc_hd__a211o_1
X_4354_ _4354_/A _4354_/B _5644_/A _5645_/A vssd1 vssd1 vccd1 vccd1 _4355_/S sky130_fd_sc_hd__or4b_1
XFILLER_0_1_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3305_ _3305_/A _3305_/B vssd1 vssd1 vccd1 vccd1 _5774_/B sky130_fd_sc_hd__or2_2
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5124__A _5124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6024_ _6466_/Q _6026_/S _6023_/Y hold45/X vssd1 vssd1 vccd1 vccd1 hold46/A sky130_fd_sc_hd__a22o_1
X_4285_ _5767_/B _5767_/A vssd1 vssd1 vccd1 vccd1 _4286_/S sky130_fd_sc_hd__nand2b_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3236_ _3614_/A _3414_/B vssd1 vssd1 vccd1 vccd1 _3314_/B sky130_fd_sc_hd__nor2_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5491__A1 _4920_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3167_ _3205_/B _3167_/B _4359_/C vssd1 vssd1 vccd1 vccd1 _5344_/B sky130_fd_sc_hd__and3_2
XANTENNA__4963__A _6309_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3098_ input5/X vssd1 vssd1 vccd1 vccd1 _3098_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_55_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xci2406_z80_191 vssd1 vssd1 vccd1 vccd1 ci2406_z80_191/HI io_oeb[6] sky130_fd_sc_hd__conb_1
XFILLER_0_64_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout68 _5816_/S vssd1 vssd1 vccd1 vccd1 _5861_/S sky130_fd_sc_hd__buf_4
Xfanout79 _5863_/S vssd1 vssd1 vccd1 vccd1 _5974_/S sky130_fd_sc_hd__clkbuf_8
X_5808_ _5866_/A _6460_/Q _5866_/C vssd1 vssd1 vccd1 vccd1 _5809_/C sky130_fd_sc_hd__or3_1
XANTENNA__5546__A2 _5520_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5739_ _3096_/Y _5299_/B _5769_/S vssd1 vssd1 vccd1 vccd1 _5740_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_72_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold471 _4625_/X vssd1 vssd1 vccd1 vccd1 _6287_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold460 _6476_/Q vssd1 vssd1 vccd1 vccd1 hold460/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout90_A _4361_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3190__C1 _4557_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold482 _4574_/X vssd1 vssd1 vccd1 vccd1 _6281_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold493 _6477_/Q vssd1 vssd1 vccd1 vccd1 hold493/X sky130_fd_sc_hd__buf_1
XFILLER_0_99_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_18 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5785__A2 _5976_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5846__A1_N _5977_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4070_ _4070_/A _4070_/B vssd1 vssd1 vccd1 vccd1 _5161_/A sky130_fd_sc_hd__nand2_1
XANTENNA__5473__A1 input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4783__A _5322_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5225__A1 _6336_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5225__B2 _5016_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4972_ _6421_/Q _4793_/Y _4964_/X _4971_/X vssd1 vssd1 vccd1 vccd1 _4972_/X sky130_fd_sc_hd__a211o_1
X_3923_ _4060_/B _3920_/X _3974_/B _3922_/X vssd1 vssd1 vccd1 vccd1 _3923_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_86_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3854_ _6452_/Q _6229_/Q _3861_/S vssd1 vssd1 vccd1 vccd1 _3854_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4736__B1 wire92/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5119__A _6076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3785_ _6432_/Q _3785_/B _5317_/B vssd1 vssd1 vccd1 vccd1 _4786_/C sky130_fd_sc_hd__or3_1
XFILLER_0_54_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5524_ _5405_/A _3643_/B _5523_/X vssd1 vssd1 vccd1 vccd1 _5525_/B sky130_fd_sc_hd__o21ai_4
XFILLER_0_6_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5455_ _5455_/A _5455_/B vssd1 vssd1 vccd1 vccd1 _5457_/A sky130_fd_sc_hd__and2_1
X_4406_ hold83/A _4406_/B _4418_/C vssd1 vssd1 vccd1 vccd1 _4406_/X sky130_fd_sc_hd__or3_1
XANTENNA__3581__B _3581_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3711__A1 _5607_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5386_ _5513_/S _6033_/B vssd1 vssd1 vccd1 vccd1 _5386_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_10_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4169__S _4716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4337_ _5605_/B _4330_/X _4336_/X _5388_/A vssd1 vssd1 vccd1 vccd1 _4337_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4268_ _4268_/A _5145_/A vssd1 vssd1 vccd1 vccd1 _4268_/Y sky130_fd_sc_hd__nor2_1
X_3219_ _3219_/A _3219_/B vssd1 vssd1 vccd1 vccd1 _3219_/Y sky130_fd_sc_hd__nand2_2
XANTENNA__4898__S0 _5100_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6007_ _4435_/X hold155/X _6011_/S vssd1 vssd1 vccd1 vccd1 _6007_/X sky130_fd_sc_hd__mux2_1
X_4199_ _4199_/A _4199_/B vssd1 vssd1 vccd1 vccd1 _4199_/Y sky130_fd_sc_hd__nand2_1
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold290 _6233_/Q vssd1 vssd1 vccd1 vccd1 hold290/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4258__A2 _4324_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5211__B _6464_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4108__A _6289_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4966__A0 _4962_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4542__S _4545_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3666__B _6021_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4718__B1 _5783_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3570_ _5605_/A _3570_/B vssd1 vssd1 vccd1 vccd1 _4344_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_70_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5881__B _5970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5240_ _5151_/Y _5237_/X _5239_/X _5236_/X _5151_/B vssd1 vssd1 vccd1 vccd1 _5240_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_87_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4041__S1 _5721_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5171_ _5171_/A _5171_/B vssd1 vssd1 vccd1 vccd1 _5172_/B sky130_fd_sc_hd__xor2_1
X_4122_ _6097_/A vssd1 vssd1 vccd1 vccd1 _4122_/Y sky130_fd_sc_hd__inv_2
X_4053_ _4053_/A _4053_/B vssd1 vssd1 vccd1 vccd1 _4053_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__5446__B2 _5415_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput3 custom_settings[2] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4955_ _5964_/A _4954_/X _4942_/Y vssd1 vssd1 vccd1 vccd1 _4955_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_86_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3906_ _6355_/Q _4441_/S vssd1 vssd1 vccd1 vccd1 _4408_/S sky130_fd_sc_hd__nor2_4
XFILLER_0_19_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4421__A2 _6355_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3576__B _5777_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4886_ _6417_/Q _6365_/Q _5105_/S vssd1 vssd1 vccd1 vccd1 _4886_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4709__B1 _4714_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3837_ _6231_/Q _3731_/X _3810_/X _6254_/Q _3836_/X vssd1 vssd1 vccd1 vccd1 _3838_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_34_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3768_ _5182_/A vssd1 vssd1 vccd1 vccd1 _5264_/A sky130_fd_sc_hd__inv_2
XANTENNA__5382__B1 _6021_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3932__A1 _6285_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4688__A _6085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5507_ _5505_/Y _5507_/B vssd1 vssd1 vccd1 vccd1 _5508_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__5283__S _5489_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3699_ _3699_/A _3699_/B _5344_/B vssd1 vssd1 vccd1 vccd1 _3701_/B sky130_fd_sc_hd__and3_2
XFILLER_0_42_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6487_ _6488_/CLK _6487_/D fanout176/X vssd1 vssd1 vccd1 vccd1 _6487_/Q sky130_fd_sc_hd__dfstp_2
X_5438_ hold570/X _5437_/X _5489_/S vssd1 vssd1 vccd1 vccd1 _5438_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_2_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5685__A1 _6461_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5369_ _5369_/A _5369_/B _5369_/C _5369_/D vssd1 vssd1 vccd1 vccd1 _5523_/C sky130_fd_sc_hd__or4_1
XFILLER_0_10_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3448__B1 _4289_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3652__D _4595_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_24_wb_clk_i_A _6448_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4651__A2 _4324_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output34_A _6327_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4740_ _3994_/Y _4739_/X _4770_/S vssd1 vssd1 vccd1 vccd1 _4740_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5039__S0 _5100_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4671_ _5117_/A _4725_/B vssd1 vssd1 vccd1 vccd1 _4714_/S sky130_fd_sc_hd__nand2_8
X_3622_ _3594_/A _3594_/B _4653_/A vssd1 vssd1 vccd1 vccd1 _3622_/Y sky130_fd_sc_hd__o21ai_1
X_6410_ _6419_/CLK _6410_/D fanout173/X vssd1 vssd1 vccd1 vccd1 _6410_/Q sky130_fd_sc_hd__dfrtp_1
X_6341_ _6465_/CLK _6341_/D vssd1 vssd1 vccd1 vccd1 _6341_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3553_ _3525_/Y _3550_/X _3551_/Y hold49/X vssd1 vssd1 vccd1 vccd1 hold50/A sky130_fd_sc_hd__a22o_1
XFILLER_0_51_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3484_ hold37/X _3493_/B hold47/X _3493_/C vssd1 vssd1 vccd1 vccd1 _3484_/X sky130_fd_sc_hd__or4_1
X_6272_ _6312_/CLK _6272_/D fanout182/X vssd1 vssd1 vccd1 vccd1 _6272_/Q sky130_fd_sc_hd__dfstp_1
X_5223_ _6312_/Q _5222_/X _5244_/S vssd1 vssd1 vccd1 vccd1 _5223_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_51_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5154_ _6081_/A _5292_/S _5147_/X _5153_/X vssd1 vssd1 vccd1 vccd1 _5154_/X sky130_fd_sc_hd__a2bb2o_1
X_4105_ _6288_/Q _6289_/Q _4105_/C vssd1 vssd1 vccd1 vccd1 _4205_/S sky130_fd_sc_hd__and3_1
XANTENNA__5419__A1 _4650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5085_ _6101_/C _5084_/X _5106_/S vssd1 vssd1 vccd1 vccd1 _5085_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_2_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4036_ _4052_/A _4036_/B vssd1 vssd1 vccd1 vccd1 _4038_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4642__A2 _4611_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3587__A _5605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5987_ _3636_/C _3635_/Y _5986_/Y _3636_/B _4335_/B vssd1 vssd1 vccd1 vccd1 _5987_/X
+ sky130_fd_sc_hd__a32o_1
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4938_ _4937_/X _5101_/S vssd1 vssd1 vccd1 vccd1 _4938_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_62_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4869_ _4863_/X _4868_/X _4948_/S vssd1 vssd1 vccd1 vccd1 _4869_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_30_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5658__A1 _5732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4330__A1 _3668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5741__S _5769_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4330__B2 _5315_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6083__A1 _6101_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6083__B2 _6036_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4105__B _6289_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4872__A2 _4930_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6074__B2 _4962_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4791__A _6431_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5910_ _6423_/Q _5970_/A vssd1 vssd1 vccd1 vccd1 _5914_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_88_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5841_ _6365_/Q _6417_/Q _5892_/S vssd1 vssd1 vccd1 vccd1 _5841_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_29_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5772_ _4957_/S _5771_/Y _3503_/B vssd1 vssd1 vccd1 vccd1 _5874_/S sky130_fd_sc_hd__o21a_2
XFILLER_0_8_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4723_ _5124_/A _5757_/A _4724_/C vssd1 vssd1 vccd1 vccd1 _4723_/X sky130_fd_sc_hd__or3b_1
X_4654_ _4957_/S _5418_/C _4652_/X vssd1 vssd1 vccd1 vccd1 _4654_/Y sky130_fd_sc_hd__o21ai_4
X_4585_ _5619_/B vssd1 vssd1 vccd1 vccd1 _4585_/Y sky130_fd_sc_hd__inv_2
X_3605_ _3691_/B _5146_/D _3604_/X vssd1 vssd1 vccd1 vccd1 _3605_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_12_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3536_ _3405_/A _5617_/B _5522_/D _3535_/X vssd1 vssd1 vccd1 vccd1 _3536_/X sky130_fd_sc_hd__a31o_1
XANTENNA__4560__A1 _6309_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout103_A _3390_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6324_ _6419_/CLK _6324_/D fanout173/X vssd1 vssd1 vccd1 vccd1 _6324_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6255_ _6455_/CLK hold72/X vssd1 vssd1 vccd1 vccd1 hold71/A sky130_fd_sc_hd__dfxtp_1
X_5206_ _5206_/A _5206_/B _5200_/X vssd1 vssd1 vccd1 vccd1 _5206_/X sky130_fd_sc_hd__or3b_1
X_3467_ _5295_/A _3501_/B vssd1 vssd1 vccd1 vccd1 _3594_/B sky130_fd_sc_hd__nor2_1
X_3398_ _3617_/B _5522_/C vssd1 vssd1 vccd1 vccd1 _5311_/A sky130_fd_sc_hd__nand2_1
X_6186_ _6449_/CLK hold56/X vssd1 vssd1 vccd1 vccd1 hold55/A sky130_fd_sc_hd__dfxtp_1
X_5137_ _6345_/Q _6344_/Q vssd1 vssd1 vccd1 vccd1 _5137_/Y sky130_fd_sc_hd__nor2_1
X_5068_ _6374_/Q _5086_/C vssd1 vssd1 vccd1 vccd1 _5068_/X sky130_fd_sc_hd__xor2_1
XANTENNA__6065__B2 _6036_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6065__A1 _6101_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4019_ _6286_/Q _6288_/Q _4716_/A vssd1 vssd1 vccd1 vccd1 _5262_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_94_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5500__A0 _6464_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4595__B _4595_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6056__A1 _4366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5319__B1 _5607_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3593__A2 _3530_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4550__S _4554_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold108 _4472_/X vssd1 vssd1 vccd1 vccd1 _6184_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold119 _4436_/X vssd1 vssd1 vccd1 vccd1 _6173_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4370_ hold195/X _3954_/X _4376_/S vssd1 vssd1 vccd1 vccd1 _4370_/X sky130_fd_sc_hd__mux2_1
X_3321_ _5605_/A _4276_/A _4595_/B vssd1 vssd1 vccd1 vccd1 _3412_/B sky130_fd_sc_hd__and3_1
XANTENNA__4786__A _5322_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5381__S _5769_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3252_ _4784_/C _3307_/B _4344_/A _3252_/D vssd1 vssd1 vccd1 vccd1 _3253_/C sky130_fd_sc_hd__and4b_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6040_ _6071_/S _6039_/Y _4366_/A vssd1 vssd1 vccd1 vccd1 _6040_/Y sky130_fd_sc_hd__a21oi_4
X_3183_ _3183_/A _3316_/B vssd1 vssd1 vccd1 vccd1 _3183_/X sky130_fd_sc_hd__or2_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4058__A0 _6287_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_16_wb_clk_i _6448_/CLK vssd1 vssd1 vccd1 vccd1 _6446_/CLK sky130_fd_sc_hd__clkbuf_16
X_5824_ _5839_/A _5824_/B vssd1 vssd1 vccd1 vccd1 _5824_/X sky130_fd_sc_hd__or2_1
XFILLER_0_8_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5022__A2 _4963_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5755_ hold7/X _4146_/B _6104_/S vssd1 vssd1 vccd1 vccd1 hold8/A sky130_fd_sc_hd__mux2_1
XANTENNA__5556__S _6070_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4230__B1 _4463_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4781__A1 _4557_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4706_ _6067_/A _4714_/S vssd1 vssd1 vccd1 vccd1 _4706_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_44_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5686_ _6312_/Q _5630_/X _5653_/X _6486_/Q _5685_/X vssd1 vssd1 vccd1 vccd1 _5687_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_44_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4637_ _4146_/B _4611_/B _4602_/Y _4636_/X vssd1 vssd1 vccd1 vccd1 _4637_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_32_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold620 _6463_/Q vssd1 vssd1 vccd1 vccd1 hold620/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4568_ hold514/X _6333_/Q _4575_/S vssd1 vssd1 vccd1 vccd1 _4568_/X sky130_fd_sc_hd__mux2_1
Xhold642 _6312_/Q vssd1 vssd1 vccd1 vccd1 hold642/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold631 _6313_/Q vssd1 vssd1 vccd1 vccd1 hold631/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold653 _6349_/Q vssd1 vssd1 vccd1 vccd1 _3709_/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4696__A _6093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3519_ _3516_/X _3518_/X _5384_/A vssd1 vssd1 vccd1 vccd1 _3519_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__5291__S _5291_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6307_ _6307_/CLK _6307_/D fanout183/X vssd1 vssd1 vccd1 vccd1 _6307_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__5089__A2 _5108_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4499_ _4456_/X hold113/X _4500_/S vssd1 vssd1 vccd1 vccd1 _6208_/D sky130_fd_sc_hd__mux2_1
XANTENNA__4297__B1 _4322_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6238_ _6456_/CLK hold86/X vssd1 vssd1 vccd1 vccd1 hold85/A sky130_fd_sc_hd__dfxtp_1
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6169_ _6467_/CLK _6169_/D fanout177/X vssd1 vssd1 vccd1 vccd1 _6169_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_0_99_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3105__A _5124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6038__A1 _6101_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4049__B1 _3807_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4447__S1 _5721_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4772__A1 _6023_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4370__S _4376_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5721__B1 _5721_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6029__B2 _5478_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4545__S _4545_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3870_ _3714_/S _3717_/B _3726_/Y _3727_/Y _6227_/Q vssd1 vssd1 vccd1 vccd1 _3870_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_0_85_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3685__A _3685_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4354__D_N _5645_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5540_ _6485_/Q _5002_/B _5593_/S vssd1 vssd1 vccd1 vccd1 _5542_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_26_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5471_ _5605_/B _6365_/Q _5484_/S vssd1 vssd1 vccd1 vccd1 _5471_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4422_ _6451_/Q _6355_/Q _4420_/S hold272/X _5730_/C1 vssd1 vssd1 vccd1 vccd1 _4422_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_41_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4353_ _6435_/Q _4352_/Y _4324_/X _3284_/B vssd1 vssd1 vccd1 vccd1 _5645_/A sky130_fd_sc_hd__a2bb2o_2
X_3304_ _3326_/B _3304_/B vssd1 vssd1 vccd1 vccd1 _3305_/B sky130_fd_sc_hd__nor2_2
X_4284_ _6357_/Q _4354_/B _4605_/B vssd1 vssd1 vccd1 vccd1 _5767_/B sky130_fd_sc_hd__or3_1
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3235_ _3235_/A _3235_/B _5327_/A vssd1 vssd1 vccd1 vccd1 _3274_/B sky130_fd_sc_hd__and3_1
XANTENNA__5124__B _5322_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4279__B1 _5607_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6023_ _6023_/A _6026_/S vssd1 vssd1 vccd1 vccd1 _6023_/Y sky130_fd_sc_hd__nor2_2
XANTENNA__4818__A2 _4790_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3166_ _3326_/B _4260_/B vssd1 vssd1 vccd1 vccd1 _4784_/B sky130_fd_sc_hd__nor2_2
XANTENNA__4963__B _4963_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3097_ _3097_/A vssd1 vssd1 vccd1 vccd1 _3097_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_89_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xci2406_z80_192 vssd1 vssd1 vccd1 vccd1 ci2406_z80_192/HI io_oeb[7] sky130_fd_sc_hd__conb_1
XFILLER_0_36_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5807_ hold474/X _5785_/Y _5806_/X _5977_/S vssd1 vssd1 vccd1 vccd1 _5807_/X sky130_fd_sc_hd__a22o_1
X_3999_ _3998_/X hold287/X _4241_/S vssd1 vssd1 vccd1 vccd1 _6113_/D sky130_fd_sc_hd__mux2_1
Xfanout69 _3861_/S vssd1 vssd1 vccd1 vccd1 _3865_/S sky130_fd_sc_hd__buf_4
XFILLER_0_91_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3595__A _5387_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5738_ _5757_/B hold419/X _5611_/Y _5737_/X vssd1 vssd1 vccd1 vccd1 _5738_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_17_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5669_ _5732_/A _5669_/B vssd1 vssd1 vccd1 vccd1 _5669_/X sky130_fd_sc_hd__or2_1
Xhold472 _6432_/Q vssd1 vssd1 vccd1 vccd1 hold472/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold450 _6279_/Q vssd1 vssd1 vccd1 vccd1 hold450/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold461 _6048_/X vssd1 vssd1 vccd1 vccd1 _6476_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5315__A _5315_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold483 _6478_/Q vssd1 vssd1 vccd1 vccd1 hold483/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold494 _6052_/X vssd1 vssd1 vccd1 vccd1 _6477_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout83_A _4408_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4365__S _5769_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3489__B _3489_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3245__B2 _5398_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3245__A1 _5315_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4783__B _5146_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4971_ _5109_/A1 _4966_/X _4970_/X _4924_/C vssd1 vssd1 vccd1 vccd1 _4971_/X sky130_fd_sc_hd__a22o_1
X_3922_ _5136_/B _3916_/Y _3921_/A _3753_/X vssd1 vssd1 vccd1 vccd1 _3922_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_86_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3853_ _6205_/Q _6213_/Q _3861_/S vssd1 vssd1 vccd1 vccd1 _3853_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_73_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5119__B _5292_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3784_ _4675_/A _5369_/D vssd1 vssd1 vccd1 vccd1 _3784_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_26_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5523_ _5523_/A _5523_/B _5523_/C _5522_/X vssd1 vssd1 vccd1 vccd1 _5523_/X sky130_fd_sc_hd__or4b_4
XFILLER_0_26_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5454_ _5492_/A _5453_/B _5453_/C vssd1 vssd1 vccd1 vccd1 _5455_/B sky130_fd_sc_hd__a21o_1
X_5385_ _6023_/A _5377_/Y _5384_/Y _3088_/A _6444_/Q vssd1 vssd1 vccd1 vccd1 _5385_/X
+ sky130_fd_sc_hd__a32o_1
X_4405_ hold65/X _4404_/X _4464_/S vssd1 vssd1 vccd1 vccd1 hold66/A sky130_fd_sc_hd__mux2_1
XFILLER_0_41_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4336_ _4782_/A _5388_/B _4333_/X _5624_/A vssd1 vssd1 vccd1 vccd1 _4336_/X sky130_fd_sc_hd__a211o_1
X_4267_ _4313_/A _4267_/B vssd1 vssd1 vccd1 vccd1 _4267_/Y sky130_fd_sc_hd__nor2_1
X_4198_ _5268_/A _6385_/Q vssd1 vssd1 vccd1 vccd1 _4199_/B sky130_fd_sc_hd__nand2_1
X_3218_ _4273_/A _4268_/A vssd1 vssd1 vccd1 vccd1 _3219_/B sky130_fd_sc_hd__and2b_2
XANTENNA__4898__S1 _5100_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_31_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6422_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_6006_ _4428_/X hold294/X _6011_/S vssd1 vssd1 vccd1 vccd1 _6006_/X sky130_fd_sc_hd__mux2_1
X_3149_ _5309_/A _4335_/C _3305_/A vssd1 vssd1 vccd1 vccd1 _3187_/B sky130_fd_sc_hd__or3_1
XANTENNA__4672__B1 _4715_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3227__A1 _3168_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6478__SET_B fanout176/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5744__S _5769_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5152__B2 _5783_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5152__A1 _6334_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold280 _3474_/X vssd1 vssd1 vccd1 vccd1 _6244_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold291 _6218_/Q vssd1 vssd1 vccd1 vccd1 hold291/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_14_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_62_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4179__C1 _3701_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5143__A1 _5292_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5679__C1 _5731_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5694__A2 _5721_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5170_ _6284_/Q _5170_/B vssd1 vssd1 vccd1 vccd1 _5172_/A sky130_fd_sc_hd__xor2_1
X_4121_ _4227_/S _4120_/X _4087_/X vssd1 vssd1 vccd1 vccd1 _6097_/A sky130_fd_sc_hd__a21oi_4
XANTENNA__5446__A2 _5520_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4052_ _4052_/A _4052_/B vssd1 vssd1 vccd1 vccd1 _4053_/B sky130_fd_sc_hd__xnor2_1
Xinput4 custom_settings[3] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__buf_1
XANTENNA__4654__B1 _4652_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4944__D _6364_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4733__S _5289_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4954_ _6368_/Q _5861_/S _5842_/B1 _4953_/X vssd1 vssd1 vccd1 vccd1 _4954_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_19_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3905_ hold9/X _4462_/A2 _4463_/S vssd1 vssd1 vccd1 vccd1 _3905_/X sky130_fd_sc_hd__o21a_1
XANTENNA__4709__A1 _4713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4885_ _4922_/C _4885_/B _4924_/C vssd1 vssd1 vccd1 vccd1 _4885_/X sky130_fd_sc_hd__and3b_1
XANTENNA_fanout133_A _5777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3836_ _6454_/Q _3804_/X _3807_/X _6175_/Q vssd1 vssd1 vccd1 vccd1 _3836_/X sky130_fd_sc_hd__a22o_1
X_3767_ _4716_/A _3079_/Y _3766_/Y vssd1 vssd1 vccd1 vccd1 _5182_/A sky130_fd_sc_hd__a21o_1
XANTENNA__5382__A1 _4605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4185__A2 _3799_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3932__A2 _6286_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5506_ _5594_/A _5506_/B vssd1 vssd1 vccd1 vccd1 _5507_/B sky130_fd_sc_hd__nand2_1
XANTENNA__4688__B _4714_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3698_ _5478_/S _3700_/B vssd1 vssd1 vccd1 vccd1 _3698_/Y sky130_fd_sc_hd__nand2_2
X_6486_ _6488_/CLK _6486_/D fanout172/X vssd1 vssd1 vccd1 vccd1 _6486_/Q sky130_fd_sc_hd__dfstp_1
X_5437_ _6459_/Q _5436_/X _5512_/S vssd1 vssd1 vccd1 vccd1 _5437_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_2_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5368_ hold43/X _5367_/Y _5368_/S vssd1 vssd1 vccd1 vccd1 hold44/A sky130_fd_sc_hd__mux2_1
X_5299_ _5299_/A _5299_/B _5299_/C vssd1 vssd1 vccd1 vccd1 _5299_/X sky130_fd_sc_hd__or3_1
XFILLER_0_10_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4319_ _5232_/S _4319_/B _5783_/A _4319_/D vssd1 vssd1 vccd1 vccd1 _4320_/B sky130_fd_sc_hd__and4_1
XANTENNA__3448__A1 _4276_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6377__RESET_B fanout176/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6306__RESET_B fanout183/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5739__S _5769_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold512_A _6408_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5474__S _5567_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4884__B1 _6365_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4553__S _4554_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output27_A _5581_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4670_ _6032_/C _4670_/B _4670_/C _4670_/D vssd1 vssd1 vccd1 vccd1 _4725_/B sky130_fd_sc_hd__and4_2
XFILLER_0_43_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5039__S1 _5078_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3621_ _3603_/A _3665_/B _3620_/X vssd1 vssd1 vccd1 vccd1 _3621_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_3_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3552_ _3525_/Y _3548_/X _3551_/Y hold365/X vssd1 vssd1 vccd1 vccd1 _3552_/X sky130_fd_sc_hd__a22o_1
X_6340_ _6340_/CLK _6340_/D fanout183/X vssd1 vssd1 vccd1 vccd1 _6340_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_0_71_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3483_ _3493_/C _3472_/B _3487_/B _5995_/C vssd1 vssd1 vccd1 vccd1 _3483_/X sky130_fd_sc_hd__a22o_1
X_6271_ _6316_/CLK _6271_/D fanout174/X vssd1 vssd1 vccd1 vccd1 _6271_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_0_11_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5222_ _6336_/Q _3092_/Y _5243_/S vssd1 vssd1 vccd1 vccd1 _5222_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5667__A2 _5721_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5153_ _5151_/Y _5152_/X _5148_/X vssd1 vssd1 vccd1 vccd1 _5153_/X sky130_fd_sc_hd__a21o_1
XANTENNA__4728__S _4770_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4104_ _6333_/Q _4104_/B vssd1 vssd1 vccd1 vccd1 _4203_/A sky130_fd_sc_hd__or2_4
XFILLER_0_47_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5413__A _6458_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5084_ _6427_/Q _6375_/Q _5105_/S vssd1 vssd1 vccd1 vccd1 _5084_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4029__A _6089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4035_ _4035_/A _4035_/B vssd1 vssd1 vccd1 vccd1 _4036_/B sky130_fd_sc_hd__or2_2
XFILLER_0_2_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5559__S _5593_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4463__S _4463_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5986_ _5995_/C _5985_/X _3426_/B vssd1 vssd1 vccd1 vccd1 _5986_/Y sky130_fd_sc_hd__a21oi_1
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4937_ hold61/A _6193_/Q _6177_/Q _6256_/Q _5404_/A0 _5078_/S1 vssd1 vssd1 vccd1
+ vccd1 _4937_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_34_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4868_ _6416_/Q _6364_/Q _5105_/S vssd1 vssd1 vccd1 vccd1 _4868_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_62_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3819_ _6209_/Q _3793_/X _3816_/X _3817_/X _3818_/X vssd1 vssd1 vccd1 vccd1 _3822_/A
+ sky130_fd_sc_hd__a2111o_1
X_4799_ _6475_/Q _4794_/Y _4798_/X vssd1 vssd1 vccd1 vccd1 _4799_/X sky130_fd_sc_hd__a21o_1
XANTENNA__3905__A2 _4462_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6469_ _6470_/CLK _6469_/D fanout177/X vssd1 vssd1 vccd1 vccd1 _6469_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_30_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5291__A0 _6465_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6083__A2 _5002_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5154__A1_N _6081_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4373__S _4376_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3497__B _3497_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5897__A2 _6023_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4548__S _4554_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4085__B2 _4441_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4791__B _6442_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5379__S _5769_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5840_ _5855_/B _5840_/B vssd1 vssd1 vccd1 vccd1 _5840_/Y sky130_fd_sc_hd__nand2b_1
X_5771_ _5771_/A _5771_/B vssd1 vssd1 vccd1 vccd1 _5771_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_33_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3596__B1 _3619_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4722_ _6309_/Q _4719_/Y _4721_/X _5783_/A vssd1 vssd1 vccd1 vccd1 _4722_/X sky130_fd_sc_hd__o22a_1
XANTENNA__5337__A1 _3172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4653_ _4653_/A hold49/X vssd1 vssd1 vccd1 vccd1 _5418_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_71_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4584_ _4276_/A _4595_/B _4583_/X vssd1 vssd1 vccd1 vccd1 _5619_/B sky130_fd_sc_hd__a21bo_1
X_3604_ _3258_/B _3285_/D _4386_/B vssd1 vssd1 vccd1 vccd1 _3604_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_71_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3535_ _3205_/B _4335_/C _3305_/A _3531_/X _3534_/X vssd1 vssd1 vccd1 vccd1 _3535_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_12_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6323_ _6419_/CLK _6323_/D fanout173/X vssd1 vssd1 vccd1 vccd1 _6323_/Q sky130_fd_sc_hd__dfrtp_1
X_3466_ _6021_/S vssd1 vssd1 vccd1 vccd1 _6023_/A sky130_fd_sc_hd__inv_6
X_6254_ _6454_/CLK _6254_/D vssd1 vssd1 vccd1 vccd1 _6254_/Q sky130_fd_sc_hd__dfxtp_1
X_5205_ _3774_/A _5169_/X _5204_/X vssd1 vssd1 vccd1 vccd1 _5206_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_58_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3397_ _5398_/A _3333_/C _3379_/A _3183_/X _3514_/B vssd1 vssd1 vccd1 vccd1 _5522_/C
+ sky130_fd_sc_hd__o2111a_1
XFILLER_0_42_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6185_ _6489_/CLK _6185_/D vssd1 vssd1 vccd1 vccd1 _6185_/Q sky130_fd_sc_hd__dfxtp_1
X_5136_ _5136_/A _5136_/B vssd1 vssd1 vccd1 vccd1 _5233_/B sky130_fd_sc_hd__nor2_1
XANTENNA__4982__A _5102_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5067_ _5063_/B _5066_/X _5106_/S vssd1 vssd1 vccd1 vccd1 _5067_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6065__A2 _4920_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4018_ _6381_/Q _6385_/Q _6343_/Q vssd1 vssd1 vccd1 vccd1 _5267_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_79_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5289__S _5289_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5025__A0 _5021_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5969_ _5969_/A _5969_/B vssd1 vssd1 vccd1 vccd1 _5970_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_81_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5328__B2 _4313_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4222__A _6385_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5752__S _6104_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4730__A2_N _4720_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold109 _6151_/Q vssd1 vssd1 vccd1 vccd1 hold109/X sky130_fd_sc_hd__dlygate4sd3_1
X_3320_ _5605_/A _6430_/Q vssd1 vssd1 vccd1 vccd1 _3320_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3251_ _3174_/X _3180_/B _4273_/B _3307_/A vssd1 vssd1 vccd1 vccd1 _3253_/B sky130_fd_sc_hd__o22a_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6059__A _6093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3182_ _5387_/A _3316_/B vssd1 vssd1 vccd1 vccd1 _5774_/A sky130_fd_sc_hd__nor2_4
XANTENNA__3502__B1 hold526/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5898__A _5976_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4058__A1 _6289_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5823_ _5867_/B _5822_/C _6416_/Q vssd1 vssd1 vccd1 vccd1 _5824_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__4741__S _5232_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5754_ hold21/X _4131_/B _6104_/S vssd1 vssd1 vccd1 vccd1 hold22/A sky130_fd_sc_hd__mux2_1
X_4705_ _4715_/B2 _4701_/Y _4704_/X hold318/X _4672_/Y vssd1 vssd1 vccd1 vccd1 _4705_/X
+ sky130_fd_sc_hd__o32a_1
X_5685_ _6461_/Q _5645_/X _5684_/X _5632_/Y vssd1 vssd1 vccd1 vccd1 _5685_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_8_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4636_ _4636_/A _4641_/B vssd1 vssd1 vccd1 vccd1 _4636_/X sky130_fd_sc_hd__or2_1
Xhold610 _6337_/Q vssd1 vssd1 vccd1 vccd1 hold610/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold621 _6462_/Q vssd1 vssd1 vccd1 vccd1 hold621/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold643 _6333_/Q vssd1 vssd1 vccd1 vccd1 hold643/X sky130_fd_sc_hd__dlygate4sd3_1
X_6306_ _6307_/CLK _6306_/D fanout183/X vssd1 vssd1 vccd1 vccd1 _6306_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold654 _6470_/Q vssd1 vssd1 vccd1 vccd1 _3699_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold632 _6309_/Q vssd1 vssd1 vccd1 vccd1 hold632/X sky130_fd_sc_hd__dlygate4sd3_1
X_4567_ hold434/X _6316_/Q _4575_/S vssd1 vssd1 vccd1 vccd1 _4567_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4696__B _4714_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3518_ _4325_/C _5314_/S _3517_/Y _3285_/D _5146_/C vssd1 vssd1 vccd1 vccd1 _3518_/X
+ sky130_fd_sc_hd__o32a_1
X_4498_ _4448_/X hold99/X _4500_/S vssd1 vssd1 vccd1 vccd1 _4498_/X sky130_fd_sc_hd__mux2_1
X_3449_ _3449_/A _4328_/A _3449_/C vssd1 vssd1 vccd1 vccd1 _3450_/B sky130_fd_sc_hd__or3_1
X_6237_ _6237_/CLK _6237_/D vssd1 vssd1 vccd1 vccd1 _6237_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6168_ _6467_/CLK _6168_/D fanout177/X vssd1 vssd1 vccd1 vccd1 _6168_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_0_85_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5119_ _6076_/A _5292_/S vssd1 vssd1 vccd1 vccd1 _5119_/Y sky130_fd_sc_hd__nor2_1
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6038__A2 _6036_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6099_ hold597/X _6037_/B _6037_/Y _5587_/X vssd1 vssd1 vccd1 vccd1 _6100_/B sky130_fd_sc_hd__o22a_1
XFILLER_0_79_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3121__A _3205_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold425_A _6379_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5747__S _6104_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4772__A2 _5499_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3980__A0 _6334_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4826__S _5105_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5237__B1 _6337_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5470_ _5470_/A _5470_/B vssd1 vssd1 vccd1 vccd1 _5470_/X sky130_fd_sc_hd__xor2_2
XFILLER_0_100_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4421_ hold125/X _6355_/Q _4408_/S hold264/X _5731_/C1 vssd1 vssd1 vccd1 vccd1 _4421_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA__5712__A1 _6314_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4352_ _5607_/B2 _4351_/X _4349_/X vssd1 vssd1 vccd1 vccd1 _4352_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3303_ _4359_/C _3249_/B _5369_/D _4360_/B _4247_/A vssd1 vssd1 vccd1 vccd1 _3608_/A
+ sky130_fd_sc_hd__a2111o_1
XANTENNA__4279__A1 _3284_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4283_ _4605_/B vssd1 vssd1 vccd1 vccd1 _4283_/Y sky130_fd_sc_hd__inv_2
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3234_ _5124_/A _3268_/B _3230_/Y _3231_/X _3233_/X vssd1 vssd1 vccd1 vccd1 _5327_/A
+ sky130_fd_sc_hd__o311a_1
X_6022_ _6022_/A _6022_/B vssd1 vssd1 vccd1 vccd1 _6026_/S sky130_fd_sc_hd__nand2_4
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3165_ _3326_/B _3282_/A vssd1 vssd1 vccd1 vccd1 _5346_/A sky130_fd_sc_hd__nor2_4
XFILLER_0_55_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5779__A1 _5866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3096_ _3096_/A vssd1 vssd1 vccd1 vccd1 _3096_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_89_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout163_A hold604/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4471__S _4473_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xci2406_z80_193 vssd1 vssd1 vccd1 vccd1 ci2406_z80_193/HI io_oeb[8] sky130_fd_sc_hd__conb_1
XFILLER_0_9_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5806_ _4837_/X _5786_/Y _5798_/X _5805_/Y _5976_/S vssd1 vssd1 vccd1 vccd1 _5806_/X
+ sky130_fd_sc_hd__a32o_1
X_3998_ _3956_/X _3997_/X _4463_/S vssd1 vssd1 vccd1 vccd1 _3998_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_29_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout59 _5116_/S vssd1 vssd1 vccd1 vccd1 _5098_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_0_36_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5737_ _5737_/A _5737_/B _5737_/C vssd1 vssd1 vccd1 vccd1 _5737_/X sky130_fd_sc_hd__or3_1
XFILLER_0_72_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5668_ _6136_/Q _5721_/A2 _4235_/S _6180_/Q _5731_/C1 vssd1 vssd1 vccd1 vccd1 _5669_/B
+ sky130_fd_sc_hd__o221a_1
X_5599_ hold539/X _5598_/X _6104_/S vssd1 vssd1 vccd1 vccd1 _5599_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5703__B2 _6426_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5703__A1 _6338_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4619_ _4602_/Y _4616_/X _4618_/X vssd1 vssd1 vccd1 vccd1 _4619_/X sky130_fd_sc_hd__a21o_1
Xhold451 _4572_/X vssd1 vssd1 vccd1 vccd1 _6279_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold462 _6269_/Q vssd1 vssd1 vccd1 vccd1 hold462/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold440 _6481_/Q vssd1 vssd1 vccd1 vccd1 hold440/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold495 _6441_/Q vssd1 vssd1 vccd1 vccd1 _3633_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold473 _5992_/X vssd1 vssd1 vccd1 vccd1 _6432_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold484 _6056_/X vssd1 vssd1 vccd1 vccd1 _6478_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3116__A _4268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4690__A1 _4715_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4381__S _4385_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_1_wb_clk_i clkbuf_leaf_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6456_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_clkbuf_leaf_43_wb_clk_i_A clkbuf_leaf_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__5458__A0 _4716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4970_ _6458_/Q _4969_/Y _5108_/S vssd1 vssd1 vccd1 vccd1 _4970_/X sky130_fd_sc_hd__mux2_1
X_3921_ _3921_/A _3921_/B vssd1 vssd1 vccd1 vccd1 _3974_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_86_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3852_ _3852_/A _3852_/B _3852_/C vssd1 vssd1 vccd1 vccd1 _3852_/X sky130_fd_sc_hd__and3_1
X_5522_ _5522_/A _5522_/B _5522_/C _5522_/D vssd1 vssd1 vccd1 vccd1 _5522_/X sky130_fd_sc_hd__and4_1
XANTENNA__3944__B1 _3795_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3783_ _3734_/X _6076_/A _3700_/Y vssd1 vssd1 vccd1 vccd1 _3783_/Y sky130_fd_sc_hd__o21ai_1
X_5453_ _5492_/A _5453_/B _5453_/C vssd1 vssd1 vccd1 vccd1 _5455_/A sky130_fd_sc_hd__nand3_1
X_5384_ _5384_/A _5384_/B vssd1 vssd1 vccd1 vccd1 _5384_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__5416__A _6434_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4404_ _4418_/C _5637_/B _4402_/X vssd1 vssd1 vccd1 vccd1 _4404_/X sky130_fd_sc_hd__a21o_2
XFILLER_0_1_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6011__S _6011_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4335_ _5605_/A _4335_/B _4335_/C vssd1 vssd1 vccd1 vccd1 _5624_/A sky130_fd_sc_hd__and3_1
XANTENNA__5449__A0 _6460_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5850__S _5974_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4266_ _4328_/B _4265_/X _4258_/X vssd1 vssd1 vccd1 vccd1 _5767_/A sky130_fd_sc_hd__o21ai_4
X_4197_ _5268_/A _6385_/Q vssd1 vssd1 vccd1 vccd1 _4197_/X sky130_fd_sc_hd__or2_1
X_3217_ _5388_/A _5314_/S vssd1 vssd1 vccd1 vccd1 _3221_/C sky130_fd_sc_hd__nand2_1
XANTENNA__4672__A1 _4713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4466__S _4473_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6005_ _4416_/X hold266/X _6011_/S vssd1 vssd1 vccd1 vccd1 _6005_/X sky130_fd_sc_hd__mux2_1
X_3148_ _5371_/A _5369_/A _5369_/B vssd1 vssd1 vccd1 vccd1 _3300_/A sky130_fd_sc_hd__or3_1
XANTENNA__5151__A _5289_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3079_ _6285_/Q vssd1 vssd1 vccd1 vccd1 _3079_/Y sky130_fd_sc_hd__inv_2
XANTENNA__5621__B1 _3668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4424__A1 _5732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4188__B1 _3810_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold270 _6231_/Q vssd1 vssd1 vccd1 vccd1 hold270/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold281 _6351_/Q vssd1 vssd1 vccd1 vccd1 _6032_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold292 _6227_/Q vssd1 vssd1 vccd1 vccd1 hold292/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5760__S _5765_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4376__S _4376_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4262__A_N _5364_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3871__C1 _3883_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3926__A0 _6284_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4120_ _6463_/Q _4119_/X _6347_/Q vssd1 vssd1 vccd1 vccd1 _4120_/X sky130_fd_sc_hd__mux2_1
X_4051_ _4051_/A _4051_/B vssd1 vssd1 vccd1 vccd1 _4052_/B sky130_fd_sc_hd__or2_2
XANTENNA__6484__SET_B fanout172/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6067__A _6067_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput5 custom_settings[4] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__buf_1
XANTENNA__4654__A1 _4957_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4953_ _6368_/Q _4952_/X _5892_/S vssd1 vssd1 vccd1 vccd1 _4953_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_86_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4315__A _4322_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3904_ _4438_/A _5302_/A _3783_/Y vssd1 vssd1 vccd1 vccd1 _3904_/X sky130_fd_sc_hd__a21o_1
XANTENNA__6006__S _6011_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4884_ _6363_/Q _6364_/Q _4847_/B _6365_/Q vssd1 vssd1 vccd1 vccd1 _4885_/B sky130_fd_sc_hd__a31o_1
XFILLER_0_74_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3835_ hold99/A _3793_/X _3795_/X hold67/A vssd1 vssd1 vccd1 vccd1 _3838_/B sky130_fd_sc_hd__a22o_1
X_3766_ _5268_/A _3115_/Y _3765_/X vssd1 vssd1 vccd1 vccd1 _3766_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout126_A _4715_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6485_ _6488_/CLK _6485_/D fanout172/X vssd1 vssd1 vccd1 vccd1 _6485_/Q sky130_fd_sc_hd__dfstp_1
X_5505_ _5594_/A _5506_/B vssd1 vssd1 vccd1 vccd1 _5505_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__3365__S _6340_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3697_ _3699_/A _5478_/S _5344_/B vssd1 vssd1 vccd1 vccd1 _4418_/C sky130_fd_sc_hd__and3_4
X_5436_ _5434_/X _5435_/X _5499_/S vssd1 vssd1 vccd1 vccd1 _5436_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_2_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5367_ _6441_/Q _5367_/B vssd1 vssd1 vccd1 vccd1 _5367_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__4893__A1 _6365_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5298_ _5271_/X _5299_/C _5297_/X vssd1 vssd1 vccd1 vccd1 _5298_/Y sky130_fd_sc_hd__a21oi_1
X_4318_ _4313_/A _4319_/B _4319_/D _4320_/A vssd1 vssd1 vccd1 vccd1 _4318_/X sky130_fd_sc_hd__a31o_1
X_4249_ _4249_/A _4249_/B vssd1 vssd1 vccd1 vccd1 _5362_/C sky130_fd_sc_hd__or2_1
XFILLER_0_93_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5070__A1 _5109_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5070__B2 _4924_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5755__S _6104_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5833__B1 _5784_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5061__A1 _5101_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3620_ _4786_/B _5373_/A _3619_/X _3605_/X _5146_/C vssd1 vssd1 vccd1 vccd1 _3620_/X
+ sky130_fd_sc_hd__o32a_2
XANTENNA__5967__A1_N _5977_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4789__B _4789_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3375__A1 _3668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3551_ _3548_/X _3549_/X _3550_/X _3525_/Y vssd1 vssd1 vccd1 vccd1 _3551_/Y sky130_fd_sc_hd__o31ai_1
XFILLER_0_24_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3482_ hold47/X _3472_/B _3492_/A vssd1 vssd1 vccd1 vccd1 hold48/A sky130_fd_sc_hd__a21o_1
X_6270_ _6312_/CLK _6270_/D fanout182/X vssd1 vssd1 vccd1 vccd1 _6270_/Q sky130_fd_sc_hd__dfstp_1
X_5221_ _5147_/C _5221_/B vssd1 vssd1 vccd1 vccd1 _5221_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5152_ _6334_/Q _5132_/X _5150_/X _5783_/A vssd1 vssd1 vccd1 vccd1 _5152_/X sky130_fd_sc_hd__o22a_1
X_4103_ _6333_/Q _4104_/B vssd1 vssd1 vccd1 vccd1 _4212_/A sky130_fd_sc_hd__nor2_1
XANTENNA__5413__B _5413_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6077__B1 _4366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5083_ _6489_/Q _5104_/A2 _5082_/X vssd1 vssd1 vccd1 vccd1 _5083_/X sky130_fd_sc_hd__a21o_1
XANTENNA__4627__B2 _6313_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4627__A1 _6462_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4034_ _6114_/Q _3731_/X _3810_/X _6181_/Q _4033_/X vssd1 vssd1 vccd1 vccd1 _4035_/B
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4744__S _4768_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6525__A _6529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5985_ _6438_/Q _5995_/B _6437_/Q vssd1 vssd1 vccd1 vccd1 _5985_/X sky130_fd_sc_hd__or3b_1
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4936_ _4935_/X hold381/X _5098_/S vssd1 vssd1 vccd1 vccd1 _4936_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_74_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6001__B1 hold1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_10 _4313_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4867_ _4924_/C _4867_/B _4867_/C vssd1 vssd1 vccd1 vccd1 _4867_/X sky130_fd_sc_hd__and3_1
XFILLER_0_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3818_ _6193_/Q _3865_/S _3818_/C vssd1 vssd1 vccd1 vccd1 _3818_/X sky130_fd_sc_hd__and3_1
XFILLER_0_34_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4798_ _5413_/B _4796_/Y _4963_/B _6458_/Q vssd1 vssd1 vccd1 vccd1 _4798_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_15_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3749_ _3750_/A _3750_/B vssd1 vssd1 vccd1 vccd1 _3749_/X sky130_fd_sc_hd__or2_1
X_6468_ _6470_/CLK _6468_/D fanout177/X vssd1 vssd1 vccd1 vccd1 _6468_/Q sky130_fd_sc_hd__dfrtp_4
X_5419_ hold581/X _4650_/A _5510_/S vssd1 vssd1 vccd1 vccd1 _5419_/X sky130_fd_sc_hd__mux2_1
X_6399_ _6399_/CLK hold22/X vssd1 vssd1 vccd1 vccd1 hold21/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__4919__S _4919_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5485__S _5485_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3794__A _3852_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4306__B1 _4300_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4857__A1 _4361_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3969__A _4150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5770_ _6436_/Q _5770_/B _5770_/C _4787_/B vssd1 vssd1 vccd1 vccd1 _5771_/B sky130_fd_sc_hd__or4b_2
XFILLER_0_29_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4721_ hold466/X _4559_/B _4720_/X _3090_/Y vssd1 vssd1 vccd1 vccd1 _4721_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_44_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4652_ _5769_/S _5418_/A _4652_/C vssd1 vssd1 vccd1 vccd1 _4652_/X sky130_fd_sc_hd__and3_4
XFILLER_0_44_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5395__S _5769_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3603_ _3603_/A _3665_/B vssd1 vssd1 vccd1 vccd1 _3603_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_44_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3209__A _3304_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4583_ _5605_/B _5605_/C _3489_/B _4335_/B vssd1 vssd1 vccd1 vccd1 _4583_/X sky130_fd_sc_hd__a31o_1
X_3534_ _5345_/A _4784_/C _3534_/C _3534_/D vssd1 vssd1 vccd1 vccd1 _3534_/X sky130_fd_sc_hd__or4_1
X_6322_ _6419_/CLK _6322_/D fanout173/X vssd1 vssd1 vccd1 vccd1 _6322_/Q sky130_fd_sc_hd__dfrtp_1
X_3465_ _6025_/B _3465_/B vssd1 vssd1 vccd1 vccd1 _5975_/S sky130_fd_sc_hd__and2b_4
XANTENNA__4739__S _5289_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6253_ _6454_/CLK _6253_/D vssd1 vssd1 vccd1 vccd1 _6253_/Q sky130_fd_sc_hd__dfxtp_1
X_5204_ _3773_/Y _5180_/Y _5202_/A _6335_/Q _5290_/S vssd1 vssd1 vccd1 vccd1 _5204_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4848__B2 _4844_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3396_ _5388_/A _3396_/B vssd1 vssd1 vccd1 vccd1 _5371_/C sky130_fd_sc_hd__or2_1
XANTENNA__3520__A1 _5384_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6184_ _6239_/CLK _6184_/D vssd1 vssd1 vccd1 vccd1 _6184_/Q sky130_fd_sc_hd__dfxtp_1
X_5135_ _5268_/A _4193_/B _4196_/Y vssd1 vssd1 vccd1 vccd1 _5138_/S sky130_fd_sc_hd__a21bo_1
XFILLER_0_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4982__B _4982_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5066_ _6426_/Q _6374_/Q _5105_/S vssd1 vssd1 vccd1 vccd1 _5066_/X sky130_fd_sc_hd__mux2_1
X_4017_ _6334_/Q _4107_/C _4013_/Y _4016_/Y vssd1 vssd1 vccd1 vccd1 _5175_/B sky130_fd_sc_hd__a31o_1
XFILLER_0_74_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5273__A1 _6339_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5968_ _5959_/B _5961_/B _5959_/A vssd1 vssd1 vccd1 vccd1 _5969_/B sky130_fd_sc_hd__o21ba_1
XFILLER_0_47_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4919_ _4918_/X _4917_/X _4919_/S vssd1 vssd1 vccd1 vccd1 _4920_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_35_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5899_ _5912_/A _5898_/Y _5896_/X _5897_/X vssd1 vssd1 vccd1 vccd1 _5899_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_35_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3339__A1 _3489_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4222__B _5374_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5334__A _5757_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4839__A1 _4957_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold572_A _6409_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4384__S _4385_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6361__RESET_B fanout175/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6104__S _6104_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5943__S _5976_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3250_ _5315_/A _4784_/B vssd1 vssd1 vccd1 vccd1 _3252_/D sky130_fd_sc_hd__nand2_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3181_ _3323_/A _3229_/A _3205_/B _3168_/B vssd1 vssd1 vccd1 vccd1 _3316_/B sky130_fd_sc_hd__or4b_4
XANTENNA__3502__A1 _5567_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5822_ _6416_/Q _5867_/B _5822_/C vssd1 vssd1 vccd1 vccd1 _5839_/A sky130_fd_sc_hd__and3_1
X_5753_ hold25/X _4052_/B _6104_/S vssd1 vssd1 vccd1 vccd1 hold26/A sky130_fd_sc_hd__mux2_1
XFILLER_0_29_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4704_ _4713_/A _4703_/X _4714_/S vssd1 vssd1 vccd1 vccd1 _4704_/X sky130_fd_sc_hd__o21a_1
XANTENNA__6014__S _6019_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4861__S0 _5404_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4230__A2 _4462_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5684_ _4434_/X _5680_/X _4041_/X _5683_/X _5655_/B _5734_/S vssd1 vssd1 vccd1 vccd1
+ _5684_/X sky130_fd_sc_hd__mux4_2
XFILLER_0_71_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4635_ _5393_/A1 hold506/X _4582_/Y _4634_/X vssd1 vssd1 vccd1 vccd1 _4635_/X sky130_fd_sc_hd__a22o_1
Xhold611 _6294_/Q vssd1 vssd1 vccd1 vccd1 hold611/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold600 _3544_/X vssd1 vssd1 vccd1 vccd1 _6130_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_25_wb_clk_i _6448_/CLK vssd1 vssd1 vccd1 vccd1 _6462_/CLK sky130_fd_sc_hd__clkbuf_16
X_4566_ hold438/X _6315_/Q _4575_/S vssd1 vssd1 vccd1 vccd1 _4566_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_8_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3517_ _5522_/A _4338_/B _4324_/B vssd1 vssd1 vccd1 vccd1 _3517_/Y sky130_fd_sc_hd__a21oi_1
X_6305_ _6307_/CLK _6305_/D fanout183/X vssd1 vssd1 vccd1 vccd1 _6305_/Q sky130_fd_sc_hd__dfrtp_1
Xhold622 _6474_/Q vssd1 vssd1 vccd1 vccd1 hold622/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold633 _4729_/X vssd1 vssd1 vccd1 vccd1 _6309_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold644 _6360_/Q vssd1 vssd1 vccd1 vccd1 hold644/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4469__S _4473_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5730__A2 _4406_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold655 _6429_/Q vssd1 vssd1 vccd1 vccd1 hold655/X sky130_fd_sc_hd__dlygate4sd3_1
X_4497_ _4441_/X hold197/X _4500_/S vssd1 vssd1 vccd1 vccd1 _4497_/X sky130_fd_sc_hd__mux2_1
X_3448_ _4276_/A _3590_/A _4289_/B _3446_/Y _3786_/A vssd1 vssd1 vccd1 vccd1 _3449_/C
+ sky130_fd_sc_hd__a2111o_1
X_6236_ _6456_/CLK hold70/X vssd1 vssd1 vccd1 vccd1 hold69/A sky130_fd_sc_hd__dfxtp_1
X_3379_ _3379_/A _3379_/B _3379_/C _3379_/D vssd1 vssd1 vccd1 vccd1 _3379_/X sky130_fd_sc_hd__and4_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6167_ _6167_/CLK _6167_/D fanout179/X vssd1 vssd1 vccd1 vccd1 _6167_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_0_85_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5118_ _6032_/B _6032_/C _6073_/A _6032_/A vssd1 vssd1 vccd1 vccd1 _5292_/S sky130_fd_sc_hd__or4b_4
XANTENNA__5246__A1 _6338_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5246__B2 _4957_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4049__A2 _3804_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6098_ _4366_/A _6096_/X _6097_/Y hold468/X _6077_/Y vssd1 vssd1 vccd1 vccd1 _6098_/X
+ sky130_fd_sc_hd__o32a_1
X_5049_ _6462_/Q _5108_/S _5048_/Y vssd1 vssd1 vccd1 vccd1 _5049_/X sky130_fd_sc_hd__o21a_1
XANTENNA__4217__B _6284_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_2_3__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6448_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_79_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5763__S _5765_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4379__S _4385_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5721__A2 _5721_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_33_wb_clk_i_A clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__5064__A _5064_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3496__B1 _4325_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5237__A1 _4716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4996__A0 _6459_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4748__B1 wire92/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5239__A _5783_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4843__S0 _5404_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4420_ _6212_/Q _6204_/Q _4420_/S vssd1 vssd1 vccd1 vccd1 _4420_/X sky130_fd_sc_hd__mux2_1
X_4351_ _5398_/A _4326_/Y _4328_/X _4350_/X vssd1 vssd1 vccd1 vccd1 _4351_/X sky130_fd_sc_hd__a211o_1
X_3302_ _5387_/A _3639_/C vssd1 vssd1 vccd1 vccd1 _3302_/X sky130_fd_sc_hd__or2_1
X_4282_ _4282_/A _4282_/B vssd1 vssd1 vccd1 vccd1 _4605_/B sky130_fd_sc_hd__nand2_4
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3233_ _3226_/X _3227_/Y _3228_/X _3219_/Y _3232_/X vssd1 vssd1 vccd1 vccd1 _3233_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA__4279__A2 _4324_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6021_ _3469_/A _6020_/X _6021_/S vssd1 vssd1 vccd1 vccd1 _6022_/B sky130_fd_sc_hd__mux2_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3164_ _5371_/B _5600_/B vssd1 vssd1 vccd1 vccd1 _5345_/C sky130_fd_sc_hd__or2_2
XANTENNA__5228__A1 _6336_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5779__A2 _5866_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6009__S _6011_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3095_ _6369_/Q vssd1 vssd1 vccd1 vccd1 _4968_/A sky130_fd_sc_hd__inv_2
XFILLER_0_89_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4752__S _4770_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout156_A _3284_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xci2406_z80_194 vssd1 vssd1 vccd1 vccd1 ci2406_z80_194/HI io_oeb[9] sky130_fd_sc_hd__conb_1
XFILLER_0_9_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5805_ _5805_/A _5813_/B vssd1 vssd1 vccd1 vccd1 _5805_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_9_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3997_ hold17/X _4462_/A2 _3996_/X vssd1 vssd1 vccd1 vccd1 _3997_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_91_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5736_ _6428_/Q _5643_/X _5645_/X _6465_/Q _5735_/X vssd1 vssd1 vccd1 vccd1 _5737_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_60_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5667_ _6220_/Q _5721_/A2 _4235_/S _6113_/Q _5730_/C1 vssd1 vssd1 vccd1 vccd1 _5667_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4618_ hold493/X _4604_/X _4605_/X hold363/X _4617_/X vssd1 vssd1 vccd1 vccd1 _4618_/X
+ sky130_fd_sc_hd__a221o_1
X_5598_ _6465_/Q _5597_/X _5598_/S vssd1 vssd1 vccd1 vccd1 _5598_/X sky130_fd_sc_hd__mux2_1
Xhold452 _6284_/Q vssd1 vssd1 vccd1 vccd1 hold452/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold430 _5688_/X vssd1 vssd1 vccd1 vccd1 _6381_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold463 _4562_/X vssd1 vssd1 vccd1 vccd1 _6269_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4549_ _3998_/X hold207/X _4554_/S vssd1 vssd1 vccd1 vccd1 _6261_/D sky130_fd_sc_hd__mux2_1
Xhold441 _6068_/X vssd1 vssd1 vccd1 vccd1 _6481_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold496 _3634_/B vssd1 vssd1 vccd1 vccd1 _5978_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold485 _6280_/Q vssd1 vssd1 vccd1 vccd1 hold485/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold474 _6414_/Q vssd1 vssd1 vccd1 vccd1 hold474/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3116__B _4273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6219_ _6263_/CLK _6219_/D vssd1 vssd1 vccd1 vccd1 _6219_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5467__A1 _5492_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5612__A _5645_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3132__A _4675_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5758__S _5765_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5078__S0 _5404_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4902__B1 _4789_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5458__A1 _6364_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3920_ _3921_/A _3921_/B vssd1 vssd1 vccd1 vccd1 _3920_/X sky130_fd_sc_hd__or2_1
XFILLER_0_46_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3696__B _5344_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3851_ _6173_/Q _3884_/S _3850_/X _3885_/A vssd1 vssd1 vccd1 vccd1 _3852_/C sky130_fd_sc_hd__a211o_1
X_3782_ _6076_/A vssd1 vssd1 vccd1 vccd1 _3782_/Y sky130_fd_sc_hd__inv_2
XANTENNA__5394__B1 _5644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5521_ _5521_/A _5521_/B vssd1 vssd1 vccd1 vccd1 _5521_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_81_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5452_ _6478_/Q _4863_/X _5593_/S vssd1 vssd1 vccd1 vccd1 _5453_/C sky130_fd_sc_hd__mux2_1
XANTENNA__4601__A _5767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6464__RESET_B fanout181/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5383_ _6032_/B _5382_/Y _5513_/S vssd1 vssd1 vccd1 vccd1 _5383_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5416__B _5478_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4403_ hold126/X hold75/X hold55/X hold57/X _4420_/S _5731_/C1 vssd1 vssd1 vccd1
+ vccd1 _5637_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_10_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3217__A _5388_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4334_ _6429_/Q _3632_/D _4253_/Y vssd1 vssd1 vccd1 vccd1 _5362_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_10_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4747__S _5232_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4265_ _5605_/B _4261_/Y _4264_/X _3219_/B _4281_/B vssd1 vssd1 vccd1 vccd1 _4265_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_5_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6528__A _6529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6004_ _4404_/X hold250/X _6011_/S vssd1 vssd1 vccd1 vccd1 _6004_/X sky130_fd_sc_hd__mux2_1
X_4196_ _4196_/A _5158_/B vssd1 vssd1 vccd1 vccd1 _4196_/Y sky130_fd_sc_hd__nand2_1
X_3216_ _3229_/A _3216_/B _5388_/A vssd1 vssd1 vccd1 vccd1 _5364_/A sky130_fd_sc_hd__and3_4
XANTENNA__4672__A2 _4714_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3147_ _5369_/B vssd1 vssd1 vccd1 vccd1 _5124_/C sky130_fd_sc_hd__inv_2
XANTENNA__4409__C1 _5731_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3078_ _4150_/A vssd1 vssd1 vccd1 vccd1 _4199_/A sky130_fd_sc_hd__inv_2
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5621__A1 _4325_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4482__S _4482_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_40_wb_clk_i clkbuf_leaf_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6483_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_5719_ _5719_/A _5719_/B vssd1 vssd1 vccd1 vccd1 _5719_/X sky130_fd_sc_hd__or2_1
XANTENNA__5688__A1 _5757_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold271 _6174_/Q vssd1 vssd1 vccd1 vccd1 hold271/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold260 _6177_/Q vssd1 vssd1 vccd1 vccd1 hold260/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 _5383_/X vssd1 vssd1 vccd1 vccd1 _6351_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold293 _4521_/X vssd1 vssd1 vccd1 vccd1 _6227_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_hold652_A _6355_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4663__A2 _4652_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4392__S _4397_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4415__A2 _4462_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3926__A1 _6286_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4351__A1 _5398_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5332__A_N _5757_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4050_ _6115_/Q _3731_/X _3810_/X _6182_/Q _4049_/X vssd1 vssd1 vccd1 vccd1 _4051_/B
+ sky130_fd_sc_hd__a221o_1
Xinput6 io_in[22] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_78_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4952_ _6420_/Q _4793_/Y _4946_/X _4951_/X vssd1 vssd1 vccd1 vccd1 _4952_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_74_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3903_ _3903_/A _3903_/B vssd1 vssd1 vccd1 vccd1 _5302_/A sky130_fd_sc_hd__xnor2_1
X_4883_ _6364_/Q _6365_/Q _4883_/C vssd1 vssd1 vccd1 vccd1 _4922_/C sky130_fd_sc_hd__and3_1
XFILLER_0_52_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3834_ _6239_/Q _3799_/X _3801_/X _6191_/Q vssd1 vssd1 vccd1 vccd1 _3838_/A sky130_fd_sc_hd__a22o_1
X_3765_ _3511_/A _6333_/Q _4595_/B _4217_/A vssd1 vssd1 vccd1 vccd1 _3765_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_54_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4590__A1 _4276_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4590__B2 _3205_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4331__A _5605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3696_ _3699_/A _5344_/B vssd1 vssd1 vccd1 vccd1 _3700_/B sky130_fd_sc_hd__and2_1
XANTENNA__5427__A _6469_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6484_ _6488_/CLK _6484_/D fanout172/X vssd1 vssd1 vccd1 vccd1 _6484_/Q sky130_fd_sc_hd__dfstp_1
X_5504_ _6482_/Q _4942_/B _5593_/S vssd1 vssd1 vccd1 vccd1 _5506_/B sky130_fd_sc_hd__mux2_1
X_5435_ hold570/X _4656_/A _5510_/S vssd1 vssd1 vccd1 vccd1 _5435_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_42_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5366_ _5393_/A1 hold617/X _5368_/S _5365_/X vssd1 vssd1 vccd1 vccd1 _6347_/D sky130_fd_sc_hd__a22o_1
XANTENNA__4342__B2 _4782_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4893__A2 _5816_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5297_ _5294_/X _5299_/C _5757_/B vssd1 vssd1 vccd1 vccd1 _5297_/X sky130_fd_sc_hd__a21o_1
X_4317_ _4319_/B _4316_/Y _5232_/S vssd1 vssd1 vccd1 vccd1 _4317_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4477__S _4482_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4248_ _6430_/Q _4248_/B _4248_/C vssd1 vssd1 vccd1 vccd1 _4249_/B sky130_fd_sc_hd__and3_1
XANTENNA__6095__A1 _6101_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6095__B2 _6036_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4645__A2 _5268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5842__A1 _6365_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4179_ _4438_/A _5304_/B _4178_/Y _3701_/B vssd1 vssd1 vccd1 vccd1 _4179_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_77_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5101__S _5101_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4581__A1 _5767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6490__SET_B fanout176/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4884__A2 _6364_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6086__A1 _4366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3304__B _3304_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6107__S _6107_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3320__A _5605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4151__A _6290_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4572__A1 _6337_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3550_ _5605_/B _3652_/B _5388_/A vssd1 vssd1 vccd1 vccd1 _3550_/X sky130_fd_sc_hd__and3_1
XFILLER_0_3_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3481_ _3489_/B _3481_/B _3488_/B vssd1 vssd1 vccd1 vccd1 _3492_/A sky130_fd_sc_hd__and3_1
X_5220_ hold636/X _5219_/X _5489_/S vssd1 vssd1 vccd1 vccd1 _6335_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_51_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6275__SET_B fanout183/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5151_ _5289_/S _5151_/B vssd1 vssd1 vccd1 vccd1 _5151_/Y sky130_fd_sc_hd__nor2_1
X_4102_ _6289_/Q _6290_/Q _4101_/B _5268_/A vssd1 vssd1 vccd1 vccd1 _4104_/B sky130_fd_sc_hd__o31a_1
X_5082_ _6315_/Q _4963_/B _6101_/C _4796_/Y vssd1 vssd1 vccd1 vccd1 _5082_/X sky130_fd_sc_hd__a22o_1
X_4033_ _6221_/Q _3804_/X _3807_/X _6137_/Q vssd1 vssd1 vccd1 vccd1 _4033_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3835__B1 _3795_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6017__S _6019_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5984_ _3786_/A _3636_/B _3635_/Y _5983_/Y vssd1 vssd1 vccd1 vccd1 _6429_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_74_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4935_ _6126_/Q _4934_/X _5016_/S vssd1 vssd1 vccd1 vccd1 _4935_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6001__A1 _5384_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4866_ _6364_/Q _4883_/C vssd1 vssd1 vccd1 vccd1 _4867_/C sky130_fd_sc_hd__or2_1
XANTENNA__4012__B1 _6287_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4797_ _4802_/D _4802_/B _4802_/C vssd1 vssd1 vccd1 vccd1 _4963_/B sky130_fd_sc_hd__and3b_4
XFILLER_0_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3817_ hold61/A _3884_/S _3818_/C vssd1 vssd1 vccd1 vccd1 _3817_/X sky130_fd_sc_hd__and3_1
X_3748_ _4150_/A _3747_/X _3748_/S vssd1 vssd1 vccd1 vccd1 _3750_/B sky130_fd_sc_hd__mux2_1
XANTENNA__4563__A1 _6312_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5760__A0 _6311_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3679_ _5146_/C _3667_/X _3678_/X vssd1 vssd1 vccd1 vccd1 _5296_/A sky130_fd_sc_hd__o21ai_4
X_6467_ _6467_/CLK _6467_/D fanout177/X vssd1 vssd1 vccd1 vccd1 _6467_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__5591__S _6104_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5418_ _5418_/A _5418_/B _5418_/C vssd1 vssd1 vccd1 vccd1 _5510_/S sky130_fd_sc_hd__and3_4
XANTENNA__5512__A0 _6465_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6398_ _6399_/CLK hold26/X vssd1 vssd1 vccd1 vccd1 hold25/A sky130_fd_sc_hd__dfxtp_1
X_5349_ _3326_/B _3297_/B _5347_/X _5348_/X vssd1 vssd1 vccd1 vccd1 _5350_/B sky130_fd_sc_hd__o31a_1
XANTENNA__6068__A1 _4366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3124__B _3168_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4935__S _5016_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3794__B _3883_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5503__B1 _5492_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4306__A1 _4310_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4857__A2 _4844_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5806__B2 _5976_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4845__S _5105_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4720_ _5866_/A _5124_/C _4720_/C _6021_/S vssd1 vssd1 vccd1 vccd1 _4720_/X sky130_fd_sc_hd__or4_4
X_4651_ _5995_/C _4324_/B _5567_/B vssd1 vssd1 vccd1 vccd1 _4652_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_71_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3602_ _6529_/A _3602_/B vssd1 vssd1 vccd1 vccd1 _3665_/B sky130_fd_sc_hd__or2_1
X_4582_ _5757_/B _4582_/B vssd1 vssd1 vccd1 vccd1 _4582_/Y sky130_fd_sc_hd__nor2_2
XANTENNA__4312__C _5418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3533_ _6447_/Q _5309_/A _5774_/A _5370_/B vssd1 vssd1 vccd1 vccd1 _3534_/D sky130_fd_sc_hd__a211o_1
XFILLER_0_3_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6321_ _6407_/CLK _6321_/D fanout170/X vssd1 vssd1 vccd1 vccd1 _6321_/Q sky130_fd_sc_hd__dfrtp_1
X_3464_ _3464_/A _3464_/B _3464_/C _3464_/D vssd1 vssd1 vccd1 vccd1 _3465_/B sky130_fd_sc_hd__or4_1
X_6252_ _6472_/CLK _6252_/D vssd1 vssd1 vccd1 vccd1 _6252_/Q sky130_fd_sc_hd__dfxtp_1
X_5203_ _4115_/A _5189_/X _5195_/Y _3770_/A vssd1 vssd1 vccd1 vccd1 _5206_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_58_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6183_ _6223_/CLK _6183_/D vssd1 vssd1 vccd1 vccd1 _6183_/Q sky130_fd_sc_hd__dfxtp_1
X_3395_ _3326_/B _5314_/S _3376_/B vssd1 vssd1 vccd1 vccd1 _3617_/B sky130_fd_sc_hd__o21a_1
X_5134_ hold306/X _5290_/S _5133_/X vssd1 vssd1 vccd1 vccd1 _5134_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_58_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5065_ _6488_/Q _5104_/A2 _4963_/B _6314_/Q _5064_/Y vssd1 vssd1 vccd1 vccd1 _5065_/X
+ sky130_fd_sc_hd__a221o_1
X_4016_ _4016_/A _4016_/B vssd1 vssd1 vccd1 vccd1 _4016_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_2_2__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_2__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
X_5967_ _5977_/S _5966_/X _5784_/X hold546/X vssd1 vssd1 vccd1 vccd1 _5967_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_90_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4490__S _4491_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4918_ _6208_/Q hold89/A _6455_/Q _6232_/Q _6360_/Q _6129_/Q vssd1 vssd1 vccd1 vccd1
+ _4918_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_62_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5898_ _5976_/S _5898_/B vssd1 vssd1 vccd1 vccd1 _5898_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_35_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4849_ _6363_/Q _4847_/B _4924_/C vssd1 vssd1 vccd1 vccd1 _4850_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_7_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_23_wb_clk_i_A _6448_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3119__B _3168_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5321__A1_N _3205_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout99_A _4791_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3578__A2 _5146_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4775__A1 _5866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5525__A _5593_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3180_ _3304_/B _3180_/B vssd1 vssd1 vccd1 vccd1 _3185_/A sky130_fd_sc_hd__or2_1
XANTENNA__3502__A2 _6019_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5821_ _5866_/A _6461_/Q _5866_/C vssd1 vssd1 vccd1 vccd1 _5822_/C sky130_fd_sc_hd__or3_1
XFILLER_0_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5752_ hold15/X _4036_/B _6104_/S vssd1 vssd1 vccd1 vccd1 hold16/A sky130_fd_sc_hd__mux2_1
XANTENNA__4604__A _5767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4703_ _6285_/Q _4702_/X _4712_/S vssd1 vssd1 vccd1 vccd1 _4703_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_60_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4861__S1 _5078_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5683_ _5683_/A _5683_/B vssd1 vssd1 vccd1 vccd1 _5683_/X sky130_fd_sc_hd__or2_1
X_4634_ _4602_/Y _4631_/X _4633_/X vssd1 vssd1 vccd1 vccd1 _4634_/X sky130_fd_sc_hd__a21o_1
Xhold612 _6345_/Q vssd1 vssd1 vccd1 vccd1 hold612/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold601 _6366_/Q vssd1 vssd1 vccd1 vccd1 hold601/X sky130_fd_sc_hd__dlygate4sd3_1
X_4565_ hold454/X _6314_/Q _4575_/S vssd1 vssd1 vccd1 vccd1 _4565_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_8_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3516_ _3513_/X _3515_/X _5322_/A vssd1 vssd1 vccd1 vccd1 _3516_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_69_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6304_ _6307_/CLK _6304_/D fanout183/X vssd1 vssd1 vccd1 vccd1 _6304_/Q sky130_fd_sc_hd__dfrtp_1
Xhold634 _6339_/Q vssd1 vssd1 vccd1 vccd1 _3064_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold645 _6334_/Q vssd1 vssd1 vccd1 vccd1 hold645/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold623 _3650_/Y vssd1 vssd1 vccd1 vccd1 _6474_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout101_A _5499_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold656 _6296_/Q vssd1 vssd1 vccd1 vccd1 hold656/X sky130_fd_sc_hd__dlygate4sd3_1
X_4496_ _4435_/X hold123/X _4500_/S vssd1 vssd1 vccd1 vccd1 _4496_/X sky130_fd_sc_hd__mux2_1
X_3447_ _3587_/B _3619_/C vssd1 vssd1 vccd1 vccd1 _4328_/A sky130_fd_sc_hd__nor2_2
X_6235_ _6237_/CLK hold84/X vssd1 vssd1 vccd1 vccd1 hold83/A sky130_fd_sc_hd__dfxtp_1
X_3378_ _3786_/A _6432_/Q _3557_/B _5317_/B vssd1 vssd1 vccd1 vccd1 _3379_/D sky130_fd_sc_hd__or4_1
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6166_ _6166_/CLK _6169_/D fanout177/X vssd1 vssd1 vccd1 vccd1 _6166_/Q sky130_fd_sc_hd__dfstp_1
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5117_ _5117_/A _6033_/B _4670_/C vssd1 vssd1 vccd1 vccd1 _6073_/A sky130_fd_sc_hd__or3b_1
XANTENNA__4485__S _4491_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6097_ _6097_/A _6107_/S vssd1 vssd1 vccd1 vccd1 _6097_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__5170__A _6284_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5048_ _5086_/C _5047_/Y _5108_/S vssd1 vssd1 vccd1 vccd1 _5048_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__3402__B _3489_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4454__B1 _4463_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4233__B _4406_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5064__B _5064_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4693__A0 _6385_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3496__A1 _5757_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4395__S _4397_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5945__A0 _6407_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4843__S1 _5078_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4350_ _3278_/A _4251_/B _5605_/D _5605_/C vssd1 vssd1 vccd1 vccd1 _4350_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_1_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3301_ _5387_/A _3639_/C vssd1 vssd1 vccd1 vccd1 _5369_/D sky130_fd_sc_hd__nor2_2
X_4281_ _4281_/A _4281_/B _4281_/C _4262_/B vssd1 vssd1 vccd1 vccd1 _4282_/B sky130_fd_sc_hd__or4b_2
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3232_ _4557_/C _3376_/B _3232_/C _4248_/C vssd1 vssd1 vccd1 vccd1 _3232_/X sky130_fd_sc_hd__or4_1
X_6020_ _4325_/A hold185/X _3374_/Y _3620_/X _3704_/B vssd1 vssd1 vccd1 vccd1 _6020_/X
+ sky130_fd_sc_hd__o32a_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4684__B1 _4714_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3163_ _3163_/A _3414_/B vssd1 vssd1 vccd1 vccd1 _5600_/B sky130_fd_sc_hd__nor2_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3094_ _6363_/Q vssd1 vssd1 vccd1 vccd1 _3094_/Y sky130_fd_sc_hd__inv_2
XANTENNA__5633__C1 _5731_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5804_ _5804_/A _5804_/B vssd1 vssd1 vccd1 vccd1 _5813_/B sky130_fd_sc_hd__nor2_1
Xci2406_z80_195 vssd1 vssd1 vccd1 vccd1 ci2406_z80_195/HI io_oeb[10] sky130_fd_sc_hd__conb_1
XANTENNA_fanout149_A _6297_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3996_ _3734_/X _5303_/A _3995_/Y vssd1 vssd1 vccd1 vccd1 _3996_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_17_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5735_ _6420_/Q _5646_/X _5734_/X _5632_/Y vssd1 vssd1 vccd1 vccd1 _5735_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_95_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5666_ _6335_/Q _5628_/X _5643_/X _6423_/Q vssd1 vssd1 vccd1 vccd1 _5674_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_44_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4617_ _6460_/Q _4606_/X _4607_/X _6311_/Q vssd1 vssd1 vccd1 vccd1 _4617_/X sky130_fd_sc_hd__a22o_1
Xhold420 _5738_/X vssd1 vssd1 vccd1 vccd1 _6385_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5597_ hold539/X _5596_/X _6070_/A vssd1 vssd1 vccd1 vccd1 _5597_/X sky130_fd_sc_hd__mux2_1
Xhold453 _4610_/X vssd1 vssd1 vccd1 vccd1 _6284_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold431 _6435_/Q vssd1 vssd1 vccd1 vccd1 _4324_/A sky130_fd_sc_hd__clkbuf_2
X_4548_ _3954_/X hold239/X _4554_/S vssd1 vssd1 vccd1 vccd1 _6260_/D sky130_fd_sc_hd__mux2_1
Xhold442 _6479_/Q vssd1 vssd1 vccd1 vccd1 hold442/X sky130_fd_sc_hd__buf_1
XFILLER_0_40_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold486 _4573_/X vssd1 vssd1 vccd1 vccd1 _6280_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold475 _5807_/X vssd1 vssd1 vccd1 vccd1 _6414_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4479_ hold211/X _4441_/X _4482_/S vssd1 vssd1 vccd1 vccd1 _4479_/X sky130_fd_sc_hd__mux2_1
Xhold464 _6126_/Q vssd1 vssd1 vccd1 vccd1 _4320_/A sky130_fd_sc_hd__buf_1
Xhold497 _5987_/X vssd1 vssd1 vccd1 vccd1 _6430_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6218_ _6489_/CLK _6218_/D vssd1 vssd1 vccd1 vccd1 _6218_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6149_ _6490_/CLK _6149_/D vssd1 vssd1 vccd1 vccd1 _6149_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_95_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5078__S1 _5078_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5059__B _5101_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4902__A1 _6366_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5615__C1 _5364_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3850_ _3712_/Y _3715_/Y _3725_/X _3728_/X _6252_/Q vssd1 vssd1 vccd1 vccd1 _3850_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_46_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3781_ hold489/X _4087_/B _3780_/X vssd1 vssd1 vccd1 vccd1 _6076_/A sky130_fd_sc_hd__a21oi_4
XFILLER_0_39_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3944__A2 _3793_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5520_ _6101_/A _5520_/B vssd1 vssd1 vccd1 vccd1 _5521_/B sky130_fd_sc_hd__or2_1
XFILLER_0_81_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4601__B _4605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5451_ _5757_/A _6461_/Q vssd1 vssd1 vccd1 vccd1 _5453_/B sky130_fd_sc_hd__or2_1
X_5382_ _4605_/B _5377_/Y _6021_/S vssd1 vssd1 vccd1 vccd1 _5382_/Y sky130_fd_sc_hd__a21oi_1
X_4402_ _6386_/Q _4462_/A2 _3783_/Y _4401_/Y _3698_/Y vssd1 vssd1 vccd1 vccd1 _4402_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA__3217__B _5314_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4333_ _3396_/B _3412_/B _5370_/D _4338_/A _4332_/X vssd1 vssd1 vccd1 vccd1 _4333_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_10_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4264_ _4675_/A _4264_/B _4264_/C vssd1 vssd1 vccd1 vccd1 _4264_/X sky130_fd_sc_hd__and3_2
X_3215_ _5315_/A _3281_/A _5360_/A vssd1 vssd1 vccd1 vccd1 _4289_/B sky130_fd_sc_hd__and3_2
XFILLER_0_66_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6003_ _6003_/A _6003_/B vssd1 vssd1 vccd1 vccd1 _6011_/S sky130_fd_sc_hd__or2_4
X_4195_ _4196_/A _5158_/B vssd1 vssd1 vccd1 vccd1 _4195_/X sky130_fd_sc_hd__or2_1
XFILLER_0_66_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3146_ _3247_/A _3282_/A vssd1 vssd1 vccd1 vccd1 _5369_/B sky130_fd_sc_hd__nor2_2
X_3077_ _6343_/Q vssd1 vssd1 vccd1 vccd1 _3740_/B sky130_fd_sc_hd__inv_2
XFILLER_0_77_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4763__S _5289_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5621__A2 _4595_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5082__B1 _6101_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5385__A1 _6023_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4188__A2 _3731_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3979_ _3979_/A _5163_/A vssd1 vssd1 vccd1 vccd1 _3991_/B sky130_fd_sc_hd__nand2_1
X_5718_ hold97/A _6355_/Q _4420_/S hold71/A _3908_/X vssd1 vssd1 vccd1 vccd1 _5719_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_72_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5649_ hold417/X _5629_/X _5641_/X _5648_/X vssd1 vssd1 vccd1 vccd1 _5649_/X sky130_fd_sc_hd__a211o_1
XANTENNA__4345__C1 _5605_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3127__B _4557_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold250 _6449_/Q vssd1 vssd1 vccd1 vccd1 hold250/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold261 _4464_/X vssd1 vssd1 vccd1 vccd1 _6177_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold283 _6134_/Q vssd1 vssd1 vccd1 vccd1 hold283/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold294 _6451_/Q vssd1 vssd1 vccd1 vccd1 hold294/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold272 _6228_/Q vssd1 vssd1 vccd1 vccd1 hold272/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold645_A _6334_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5860__A2 _4791_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5769__S _5769_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5679__A2 _4406_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4887__A0 _4881_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput7 io_in[23] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__buf_1
XFILLER_0_36_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4951_ _5109_/A1 _4948_/X _4950_/X vssd1 vssd1 vccd1 vccd1 _4951_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_86_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3500__B _3501_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4882_ _4361_/B _4881_/X _5771_/A vssd1 vssd1 vccd1 vccd1 _4882_/X sky130_fd_sc_hd__a21o_1
X_3902_ _3901_/A _3901_/B _3903_/A vssd1 vssd1 vccd1 vccd1 _3902_/Y sky130_fd_sc_hd__o21bai_2
XFILLER_0_6_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3833_ _4460_/A _4451_/A vssd1 vssd1 vccd1 vccd1 _3898_/A sky130_fd_sc_hd__and2_1
XFILLER_0_74_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3764_ _6345_/Q _3772_/B _6346_/Q vssd1 vssd1 vccd1 vccd1 _4115_/A sky130_fd_sc_hd__and3b_4
XFILLER_0_27_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4331__B _5315_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3695_ _3665_/A _5418_/A _3624_/Y _6036_/A _3694_/X vssd1 vssd1 vccd1 vccd1 _3695_/Y
+ sky130_fd_sc_hd__o2111ai_4
XANTENNA__5427__B _5427_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6483_ _6483_/CLK _6483_/D fanout176/X vssd1 vssd1 vccd1 vccd1 _6483_/Q sky130_fd_sc_hd__dfstp_1
X_5503_ _5757_/A _6465_/Q _5492_/A vssd1 vssd1 vccd1 vccd1 _5531_/A sky130_fd_sc_hd__o21a_1
X_5434_ hold570/X _5520_/B _5433_/Y _5415_/X vssd1 vssd1 vccd1 vccd1 _5434_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_42_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4758__S _4770_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5365_ _5600_/A _5362_/X _5364_/X _4289_/C _5391_/A vssd1 vssd1 vccd1 vccd1 _5365_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_58_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5296_ _5296_/A _5296_/B _5296_/C _3694_/X vssd1 vssd1 vccd1 vccd1 _5299_/C sky130_fd_sc_hd__or4b_4
X_4316_ _3093_/Y _4310_/S _4315_/X vssd1 vssd1 vccd1 vccd1 _4316_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_10_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4247_ _4247_/A _4247_/B vssd1 vssd1 vccd1 vccd1 _4249_/A sky130_fd_sc_hd__or2_1
X_4178_ _4438_/A _6067_/A vssd1 vssd1 vccd1 vccd1 _4178_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_97_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4493__S _4500_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5589__S _6070_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3129_ _3639_/C _3163_/A vssd1 vssd1 vccd1 vccd1 _4335_/C sky130_fd_sc_hd__nor2_4
XANTENNA__5055__A0 _6462_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5358__B2 _5757_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3908__A2 _4418_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4581__A2 _4605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3138__A _4268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold595_A _6365_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4869__A0 _4863_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5499__S _5499_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3844__A1 _3883_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5800__B _5867_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3320__B _6430_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3480_ _6432_/Q _3480_/B vssd1 vssd1 vccd1 vccd1 _3569_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_51_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5150_ _6276_/Q _4555_/Y _5123_/A _5149_/X vssd1 vssd1 vccd1 vccd1 _5150_/X sky130_fd_sc_hd__o22a_1
X_4101_ _6289_/Q _4101_/B vssd1 vssd1 vccd1 vccd1 _4106_/A sky130_fd_sc_hd__nor2_1
X_5081_ _5102_/A _6101_/C vssd1 vssd1 vccd1 vccd1 _5081_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__6077__A2 _6107_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5285__A0 _6340_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4032_ hold73/A _3799_/X _3801_/X _6145_/Q _4031_/X vssd1 vssd1 vccd1 vccd1 _4035_/A
+ sky130_fd_sc_hd__a221o_1
Xclkbuf_2_1__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_9_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__4607__A _4611_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5983_ _5995_/C _5981_/X _5982_/Y _5978_/Y vssd1 vssd1 vccd1 vccd1 _5983_/Y sky130_fd_sc_hd__a31oi_1
XFILLER_0_59_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5588__B2 _5415_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4934_ _6367_/Q _4933_/X _5863_/S vssd1 vssd1 vccd1 vccd1 _4934_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_86_171 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_19_wb_clk_i _6448_/CLK vssd1 vssd1 vccd1 vccd1 _6340_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_19_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4865_ _6364_/Q _4883_/C vssd1 vssd1 vccd1 vccd1 _4867_/B sky130_fd_sc_hd__nand2_1
XANTENNA__4012__A1 _6285_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout131_A _4276_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4796_ _5064_/A vssd1 vssd1 vccd1 vccd1 _4796_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_27_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3816_ _6217_/Q _3816_/B _3885_/A _3865_/S vssd1 vssd1 vccd1 vccd1 _3816_/X sky130_fd_sc_hd__and4_1
XANTENNA__4061__B _6382_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3747_ _6343_/Q _4150_/A vssd1 vssd1 vccd1 vccd1 _3747_/X sky130_fd_sc_hd__xor2_1
XANTENNA_clkbuf_leaf_13_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__3771__A0 _6378_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3678_ _3670_/Y _3675_/X _3677_/X _3669_/Y vssd1 vssd1 vccd1 vccd1 _3678_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_70_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6466_ _6467_/CLK hold46/X fanout177/X vssd1 vssd1 vccd1 vccd1 _6466_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_0_15_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4488__S _4491_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5417_ _6101_/A _5485_/S vssd1 vssd1 vccd1 vccd1 _5417_/Y sky130_fd_sc_hd__nor2_1
X_6397_ _6455_/CLK hold16/X vssd1 vssd1 vccd1 vccd1 hold15/A sky130_fd_sc_hd__dfxtp_1
X_5348_ _3057_/Y _3161_/B _3304_/B _3235_/B _3272_/B vssd1 vssd1 vccd1 vccd1 _5348_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_10_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5279_ _6459_/Q _6458_/Q _5279_/C _5279_/D vssd1 vssd1 vccd1 vccd1 _5279_/X sky130_fd_sc_hd__or4_1
XANTENNA__3421__A _4289_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4937__S0 _5404_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5503__A1 _5757_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3914__A_N _4150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5806__A2 _5786_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3331__A _4273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4760__A1_N _6315_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5990__A1 _3489_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4650_ _4650_/A _4668_/B vssd1 vssd1 vccd1 vccd1 _4650_/X sky130_fd_sc_hd__and2_1
XFILLER_0_71_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput10 io_in[26] vssd1 vssd1 vccd1 vccd1 _4658_/A sky130_fd_sc_hd__clkbuf_2
X_3601_ _3603_/A _3600_/X _3665_/A vssd1 vssd1 vccd1 vccd1 _6167_/D sky130_fd_sc_hd__mux2_1
XANTENNA__3202__C1 _6435_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4581_ _5767_/A _4605_/B _5384_/B vssd1 vssd1 vccd1 vccd1 _4582_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6320_ _6409_/CLK _6320_/D fanout170/X vssd1 vssd1 vccd1 vccd1 _6320_/Q sky130_fd_sc_hd__dfrtp_1
X_3532_ _5617_/B _4784_/B _5777_/A vssd1 vssd1 vccd1 vccd1 _3534_/C sky130_fd_sc_hd__and3b_1
XFILLER_0_12_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3463_ _3461_/X _3462_/X _3464_/C vssd1 vssd1 vccd1 vccd1 _6025_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_12_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6089__A _6089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6251_ _6449_/CLK _6251_/D vssd1 vssd1 vccd1 vccd1 _6251_/Q sky130_fd_sc_hd__dfxtp_1
X_5202_ _5202_/A vssd1 vssd1 vccd1 vccd1 _5202_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_58_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3506__A _5769_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6182_ _6400_/CLK _6182_/D vssd1 vssd1 vccd1 vccd1 _6182_/Q sky130_fd_sc_hd__dfxtp_1
X_3394_ _3394_/A _3609_/C vssd1 vssd1 vccd1 vccd1 _5372_/A sky130_fd_sc_hd__or2_1
X_5133_ _6333_/Q _5132_/X _5128_/Y _4957_/S vssd1 vssd1 vccd1 vccd1 _5133_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_58_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5064_ _5064_/A _5064_/B vssd1 vssd1 vccd1 vccd1 _5064_/Y sky130_fd_sc_hd__nor2_1
X_4015_ _3933_/Y _4014_/X _6334_/Q vssd1 vssd1 vccd1 vccd1 _4016_/B sky130_fd_sc_hd__a21o_1
XANTENNA_fanout179_A fanout180/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4771__S _5232_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5966_ _5095_/Y _5786_/Y _5965_/X _5961_/Y _5976_/S vssd1 vssd1 vccd1 vccd1 _5966_/X
+ sky130_fd_sc_hd__a32o_1
X_5897_ hold588/X _6023_/A _5976_/S vssd1 vssd1 vccd1 vccd1 _5897_/X sky130_fd_sc_hd__o21ba_1
X_4917_ hold51/X hold53/X hold97/X hold71/A _6360_/Q _6129_/Q vssd1 vssd1 vccd1 vccd1
+ _4917_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_74_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4848_ _6477_/Q _4794_/Y _4796_/Y _4844_/X _4793_/Y vssd1 vssd1 vccd1 vccd1 _4852_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_7_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4779_ _4778_/X _4777_/X _4919_/S vssd1 vssd1 vccd1 vccd1 _5413_/B sky130_fd_sc_hd__mux2_4
XFILLER_0_15_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5733__A1 _5655_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6449_ _6449_/CLK _6449_/D vssd1 vssd1 vccd1 vccd1 _6449_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold558_A _6442_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3151__A _5605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5421__A0 _6458_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4775__A2 _4774_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3983__A0 _6380_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6370__RESET_B fanout172/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5724__A1 _6464_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5488__A0 _6463_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5525__B _5525_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3699__C _5344_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5820_ _5977_/S _5819_/X _5784_/X hold397/X vssd1 vssd1 vccd1 vccd1 _5820_/X sky130_fd_sc_hd__o2bb2a_1
XANTENNA__5412__B1 _5413_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5751_ hold17/X _3962_/B _6104_/S vssd1 vssd1 vccd1 vccd1 hold18/A sky130_fd_sc_hd__mux2_1
XANTENNA__4604__B _4605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4702_ _6383_/Q _6379_/Q _4711_/S vssd1 vssd1 vccd1 vccd1 _4702_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6458__RESET_B fanout181/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5682_ _6137_/Q _5721_/A2 _5721_/B1 _6181_/Q _5721_/C1 vssd1 vssd1 vccd1 vccd1 _5683_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_4_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4633_ hold498/X _4604_/X _4605_/X hold468/X _4632_/X vssd1 vssd1 vccd1 vccd1 _4633_/X
+ sky130_fd_sc_hd__a221o_1
Xhold602 _5489_/X vssd1 vssd1 vccd1 vccd1 _6366_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3726__B1 _4463_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4564_ hold458/X _6313_/Q _4575_/S vssd1 vssd1 vccd1 vccd1 _4564_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_12_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3515_ _4332_/B _3379_/A _3541_/B _3307_/A _3514_/X vssd1 vssd1 vccd1 vccd1 _3515_/X
+ sky130_fd_sc_hd__o221a_1
X_6303_ _6308_/CLK _6303_/D fanout185/X vssd1 vssd1 vccd1 vccd1 _6303_/Q sky130_fd_sc_hd__dfrtp_1
Xhold613 _6340_/Q vssd1 vssd1 vccd1 vccd1 hold613/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold624 _6461_/Q vssd1 vssd1 vccd1 vccd1 hold624/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold635 _6311_/Q vssd1 vssd1 vccd1 vccd1 hold635/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold646 _6295_/Q vssd1 vssd1 vccd1 vccd1 hold646/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold657 _6347_/Q vssd1 vssd1 vccd1 vccd1 _4226_/S sky130_fd_sc_hd__dlygate4sd3_1
X_6234_ _6237_/CLK hold58/X vssd1 vssd1 vccd1 vccd1 hold57/A sky130_fd_sc_hd__dfxtp_1
X_4495_ _4428_/X hold130/X _4500_/S vssd1 vssd1 vccd1 vccd1 _4495_/X sky130_fd_sc_hd__mux2_1
X_3446_ _3691_/B _5777_/B vssd1 vssd1 vccd1 vccd1 _3446_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_85_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3377_ _5777_/A _3557_/B vssd1 vssd1 vccd1 vccd1 _4588_/A sky130_fd_sc_hd__nor2_1
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6165_ _6165_/CLK _6168_/D fanout177/X vssd1 vssd1 vccd1 vccd1 _6165_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA__5451__A _5757_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6096_ _6101_/A _6095_/X _6107_/S vssd1 vssd1 vccd1 vccd1 _6096_/X sky130_fd_sc_hd__o21a_1
X_5116_ _5115_/X hold409/X _5116_/S vssd1 vssd1 vccd1 vccd1 _5116_/X sky130_fd_sc_hd__mux2_1
X_5047_ _6373_/Q _5047_/B vssd1 vssd1 vccd1 vccd1 _5047_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_79_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_34_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6426_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__5597__S _6070_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5949_ _5951_/A _5970_/A vssd1 vssd1 vccd1 vccd1 _5952_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_35_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4233__C _4441_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4142__B1 _3807_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5945__A1 _6426_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3300_ _3300_/A _3300_/B _3632_/D _3300_/D vssd1 vssd1 vccd1 vccd1 _3310_/A sky130_fd_sc_hd__or4_1
XFILLER_0_1_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4280_ _4276_/A _4259_/X _4273_/X _4264_/X _5398_/A vssd1 vssd1 vccd1 vccd1 _4281_/C
+ sky130_fd_sc_hd__a32o_1
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3231_ _3268_/B _4268_/A _3249_/B vssd1 vssd1 vccd1 vccd1 _3231_/X sky130_fd_sc_hd__or3b_1
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4684__A1 _4713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3162_ _3642_/C _4359_/C vssd1 vssd1 vccd1 vccd1 _3557_/B sky130_fd_sc_hd__nand2_4
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3503__B _3503_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3093_ _6314_/Q vssd1 vssd1 vccd1 vccd1 _3093_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_49_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5803_ _5804_/A _5804_/B vssd1 vssd1 vccd1 vccd1 _5805_/A sky130_fd_sc_hd__and2_1
Xci2406_z80_196 vssd1 vssd1 vccd1 vccd1 ci2406_z80_196/HI io_oeb[11] sky130_fd_sc_hd__conb_1
XANTENNA__6292__RESET_B fanout185/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3995_ _4438_/A _6085_/A _3700_/Y vssd1 vssd1 vccd1 vccd1 _3995_/Y sky130_fd_sc_hd__o21ai_1
X_5734_ _5733_/X _4239_/X _5734_/S vssd1 vssd1 vccd1 vccd1 _5734_/X sky130_fd_sc_hd__mux2_1
X_5665_ _6460_/Q _5645_/X _5646_/X hold397/X vssd1 vssd1 vccd1 vccd1 _5674_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_88_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4616_ _3892_/B _3962_/B _4641_/B vssd1 vssd1 vccd1 vccd1 _4616_/X sky130_fd_sc_hd__mux2_1
X_5596_ hold539/X _5520_/B _5595_/Y _5415_/X vssd1 vssd1 vccd1 vccd1 _5596_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_25_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold410 _5116_/X vssd1 vssd1 vccd1 vccd1 _6332_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold432 _3485_/X vssd1 vssd1 vccd1 vccd1 hold432/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold454 _6272_/Q vssd1 vssd1 vccd1 vccd1 hold454/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold421 _6413_/Q vssd1 vssd1 vccd1 vccd1 _5792_/A sky130_fd_sc_hd__buf_1
XFILLER_0_13_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4547_ _3911_/X hold220/X _4554_/S vssd1 vssd1 vccd1 vccd1 _4547_/X sky130_fd_sc_hd__mux2_1
Xhold443 _6060_/X vssd1 vssd1 vccd1 vccd1 _6479_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold487 _6288_/Q vssd1 vssd1 vccd1 vccd1 hold487/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold476 _6270_/Q vssd1 vssd1 vccd1 vccd1 hold476/X sky130_fd_sc_hd__dlygate4sd3_1
X_4478_ hold81/X _4435_/X _4482_/S vssd1 vssd1 vccd1 vccd1 hold82/A sky130_fd_sc_hd__mux2_1
Xhold465 _4323_/X vssd1 vssd1 vccd1 vccd1 _6126_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3429_ _4324_/B _3457_/B vssd1 vssd1 vccd1 vccd1 _3431_/B sky130_fd_sc_hd__nand2_1
XANTENNA__4124__B1 _3795_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold498 _6480_/Q vssd1 vssd1 vccd1 vccd1 hold498/X sky130_fd_sc_hd__dlygate4sd3_1
X_6217_ _6456_/CLK _6217_/D vssd1 vssd1 vccd1 vccd1 _6217_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4496__S _4500_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6148_ _6400_/CLK _6148_/D vssd1 vssd1 vccd1 vccd1 _6148_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6079_ _6101_/B _4982_/B _5534_/Y _6036_/X vssd1 vssd1 vccd1 vccd1 _6079_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold423_A _6383_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4902__A2 _4790_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5863__A0 _6367_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5710__S0 _5655_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6040__B1 _4366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3929__B1 _6379_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3780_ _6347_/Q _6458_/Q _4227_/S _3779_/X vssd1 vssd1 vccd1 vccd1 _3780_/X sky130_fd_sc_hd__o211a_1
XANTENNA__5394__A2 _4948_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5450_ hold583/X _5449_/X _5489_/S vssd1 vssd1 vccd1 vccd1 _5450_/X sky130_fd_sc_hd__mux2_1
X_4401_ _4414_/A _4401_/B vssd1 vssd1 vccd1 vccd1 _4401_/Y sky130_fd_sc_hd__nor2_1
X_5381_ _6032_/A _5380_/Y _5769_/S vssd1 vssd1 vccd1 vccd1 _5381_/X sky130_fd_sc_hd__mux2_1
X_4332_ _5374_/B _4332_/B _5522_/D vssd1 vssd1 vccd1 vccd1 _4332_/X sky130_fd_sc_hd__and3_1
XFILLER_0_10_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4263_ _4263_/A _4328_/A vssd1 vssd1 vccd1 vccd1 _4281_/B sky130_fd_sc_hd__or2_1
XFILLER_0_10_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6097__A _6097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4657__A1 _4782_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3214_ _3986_/A _3514_/B vssd1 vssd1 vccd1 vccd1 _3214_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_66_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6002_ _6447_/Q _3638_/C _3648_/B hold298/X vssd1 vssd1 vccd1 vccd1 _6002_/X sky130_fd_sc_hd__a22o_1
X_4194_ _6344_/Q _6385_/Q vssd1 vssd1 vccd1 vccd1 _5158_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_66_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3145_ _3323_/A _3168_/B _3229_/A vssd1 vssd1 vccd1 vccd1 _3282_/A sky130_fd_sc_hd__nand3_4
XFILLER_0_96_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3076_ _6346_/Q vssd1 vssd1 vccd1 vccd1 _3774_/A sky130_fd_sc_hd__inv_2
XFILLER_0_89_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5082__A1 _6315_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5909__B2 _5977_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3978_ _3080_/Y _4156_/A _3972_/B _3977_/X vssd1 vssd1 vccd1 vccd1 _5163_/A sky130_fd_sc_hd__a31o_1
XFILLER_0_92_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5717_ _6455_/Q _6355_/Q _4420_/S _6232_/Q _3909_/Y vssd1 vssd1 vccd1 vccd1 _5719_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_72_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4080__A _6093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5648_ _6333_/Q _5628_/X _5630_/X _6309_/Q vssd1 vssd1 vccd1 vccd1 _5648_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_5_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5579_ hold562/X _5578_/X _6070_/A vssd1 vssd1 vccd1 vccd1 _5579_/X sky130_fd_sc_hd__mux2_1
Xhold251 _6004_/X vssd1 vssd1 vccd1 vccd1 _6449_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold240 _6224_/Q vssd1 vssd1 vccd1 vccd1 hold240/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold262 _6230_/Q vssd1 vssd1 vccd1 vccd1 hold262/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4440__S0 _5721_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold284 _6217_/Q vssd1 vssd1 vccd1 vccd1 hold284/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold273 _4522_/X vssd1 vssd1 vccd1 vccd1 _6228_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold295 _6006_/X vssd1 vssd1 vccd1 vccd1 _6451_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3424__A _4289_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4648__A1 _4653_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5115__S _6070_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout74_A _5731_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5781__C1 _6434_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3318__B _5314_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput8 io_in[24] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_2_0__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_1_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_78_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4811__A1 _4924_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4811__B2 _5109_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4950_ _6482_/Q _5104_/A2 _4963_/B _6465_/Q _4949_/Y vssd1 vssd1 vccd1 vccd1 _4950_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__6013__A0 _4656_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4881_ _4880_/X _4879_/X _5101_/S vssd1 vssd1 vccd1 vccd1 _4881_/X sky130_fd_sc_hd__mux2_4
X_3901_ _3901_/A _3901_/B vssd1 vssd1 vccd1 vccd1 _3903_/B sky130_fd_sc_hd__or2_1
XFILLER_0_74_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3832_ _4052_/A _4636_/A vssd1 vssd1 vccd1 vccd1 _4451_/A sky130_fd_sc_hd__xnor2_1
X_3763_ _4217_/A _3740_/B _4557_/C _3761_/B _6378_/Q vssd1 vssd1 vccd1 vccd1 _3763_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_54_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5502_ _5494_/B _5496_/B _5494_/A vssd1 vssd1 vccd1 vccd1 _5508_/A sky130_fd_sc_hd__o21ba_1
X_3694_ _5607_/B2 _3689_/Y _3693_/X vssd1 vssd1 vccd1 vccd1 _3694_/X sky130_fd_sc_hd__o21a_1
X_6482_ _6483_/CLK _6482_/D fanout176/X vssd1 vssd1 vccd1 vccd1 _6482_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA__5146__D _5146_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5433_ _5433_/A vssd1 vssd1 vccd1 vccd1 _5433_/Y sky130_fd_sc_hd__inv_2
X_5364_ _5364_/A _5364_/B _5364_/C vssd1 vssd1 vccd1 vccd1 _5364_/X sky130_fd_sc_hd__or3_1
XFILLER_0_2_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4315_ _4322_/B _4315_/B _4315_/C vssd1 vssd1 vccd1 vccd1 _4315_/X sky130_fd_sc_hd__or3_1
XFILLER_0_2_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5295_ _5295_/A _5295_/B vssd1 vssd1 vccd1 vccd1 _5296_/C sky130_fd_sc_hd__and2_1
XFILLER_0_10_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4059__B _6382_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4246_ _5124_/C _5757_/C vssd1 vssd1 vccd1 vccd1 _4247_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_93_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4177_ _6067_/A vssd1 vssd1 vccd1 vccd1 _4177_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_97_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3128_ _5124_/A _4273_/A _3326_/B vssd1 vssd1 vccd1 vccd1 _3163_/A sky130_fd_sc_hd__or3_2
XFILLER_0_96_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3605__A2 _5146_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3059_ _5605_/C vssd1 vssd1 vccd1 vccd1 _5315_/A sky130_fd_sc_hd__inv_6
XANTENNA_clkbuf_leaf_42_wb_clk_i_A clkbuf_leaf_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_37_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3369__A1 _6339_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4030__A2 _6089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3138__B _4273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold588_A _6421_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4713__A _4713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5349__A2 _3297_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4100_ _6288_/Q _4105_/C vssd1 vssd1 vccd1 vccd1 _4101_/B sky130_fd_sc_hd__and2_1
X_5080_ _5079_/X _5078_/X _5101_/S vssd1 vssd1 vccd1 vccd1 _6101_/C sky130_fd_sc_hd__mux2_2
XFILLER_0_47_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4031_ _6262_/Q _3793_/X _3795_/X _6197_/Q vssd1 vssd1 vccd1 vccd1 _4031_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3835__A2 _3793_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5982_ _5995_/D _5988_/B _5995_/B vssd1 vssd1 vccd1 vccd1 _5982_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__5588__A2 _5520_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4933_ _5817_/A _4932_/X _4920_/X vssd1 vssd1 vccd1 vccd1 _4933_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_86_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4864_ _5102_/A _4863_/X _4776_/Y vssd1 vssd1 vccd1 vccd1 _4864_/X sky130_fd_sc_hd__a21o_1
XANTENNA__4012__A2 _6286_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4795_ _4802_/B _4802_/D vssd1 vssd1 vccd1 vccd1 _5064_/A sky130_fd_sc_hd__or2_4
XFILLER_0_6_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3815_ _4052_/A _4600_/A vssd1 vssd1 vccd1 vccd1 _3903_/A sky130_fd_sc_hd__xnor2_1
X_3746_ _6343_/Q _6344_/Q vssd1 vssd1 vccd1 vccd1 _3772_/B sky130_fd_sc_hd__nor2_1
XANTENNA_fanout124_A hold526/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3771__A1 _6382_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6465_ _6465_/CLK _6465_/D fanout181/X vssd1 vssd1 vccd1 vccd1 _6465_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__4769__S _5289_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3677_ _3674_/A _3411_/A _5617_/A _3671_/B _3676_/X vssd1 vssd1 vccd1 vccd1 _3677_/X
+ sky130_fd_sc_hd__o221a_2
XFILLER_0_70_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5416_ _6434_/Q _5478_/S vssd1 vssd1 vccd1 vccd1 _5485_/S sky130_fd_sc_hd__nand2_4
XANTENNA_clkbuf_leaf_9_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_6396_ _6481_/CLK hold18/X vssd1 vssd1 vccd1 vccd1 hold17/A sky130_fd_sc_hd__dfxtp_1
X_5347_ _4273_/A _3206_/Y _3204_/X _3193_/X vssd1 vssd1 vccd1 vccd1 _5347_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_10_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5278_ _6461_/Q _6460_/Q _6465_/Q _6464_/Q vssd1 vssd1 vccd1 vccd1 _5279_/D sky130_fd_sc_hd__or4_1
XANTENNA__5276__A1 _6409_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4229_ _4438_/A _5304_/C _4228_/X vssd1 vssd1 vccd1 vccd1 _4229_/X sky130_fd_sc_hd__a21o_1
XANTENNA__4236__C1 _5731_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5200__A1 _6382_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5364__A _5364_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4937__S1 _5078_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5503__A2 _6465_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4711__A0 _6385_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4742__A2_N _4720_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput11 io_in[27] vssd1 vssd1 vccd1 vccd1 _4668_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4580_ _4289_/C _4576_/X _4578_/X _6159_/Q vssd1 vssd1 vccd1 vccd1 _4605_/C sky130_fd_sc_hd__a22o_1
XANTENNA__3059__A _5605_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3600_ _4653_/A _3602_/B vssd1 vssd1 vccd1 vccd1 _3600_/X sky130_fd_sc_hd__or2_1
X_3531_ _4325_/A _4784_/B _3609_/C _3413_/Y _3530_/X vssd1 vssd1 vccd1 vccd1 _3531_/X
+ sky130_fd_sc_hd__a2111o_1
XANTENNA__4950__B1 _4963_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3462_ hold77/X _3700_/A _3464_/B vssd1 vssd1 vccd1 vccd1 _3462_/X sky130_fd_sc_hd__mux2_1
X_6250_ _6452_/CLK hold80/X vssd1 vssd1 vccd1 vccd1 hold79/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6089__B _6107_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3393_ _3570_/B _5774_/B _3393_/C vssd1 vssd1 vccd1 vccd1 _3399_/B sky130_fd_sc_hd__or3_1
XANTENNA__4702__A0 _6383_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5201_ _6346_/Q _5233_/B vssd1 vssd1 vccd1 vccd1 _5202_/A sky130_fd_sc_hd__and2_2
XFILLER_0_58_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3506__B _3506_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6181_ _6223_/CLK _6181_/D vssd1 vssd1 vccd1 vccd1 _6181_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__6246__RESET_B fanout180/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5132_ _5288_/S _5132_/B vssd1 vssd1 vccd1 vccd1 _5132_/X sky130_fd_sc_hd__or2_1
X_5063_ _5102_/A _5063_/B vssd1 vssd1 vccd1 vccd1 _5063_/Y sky130_fd_sc_hd__nand2_1
X_4014_ _6285_/Q _6286_/Q _6287_/Q vssd1 vssd1 vccd1 vccd1 _4014_/X sky130_fd_sc_hd__or3_1
XFILLER_0_74_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5626__A1_N _3172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5430__A1 _5492_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5965_ _5081_/Y _5964_/Y _5771_/A vssd1 vssd1 vccd1 vccd1 _5965_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_90_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5896_ _6458_/Q _5771_/A _5895_/Y _6021_/S vssd1 vssd1 vccd1 vccd1 _5896_/X sky130_fd_sc_hd__a211o_1
X_4916_ _4915_/X hold351/X _5098_/S vssd1 vssd1 vccd1 vccd1 _4916_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_90_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4847_ _6363_/Q _4847_/B vssd1 vssd1 vccd1 vccd1 _4883_/C sky130_fd_sc_hd__and2_1
XFILLER_0_23_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4778_ hold75/A _6449_/Q _6210_/Q _6226_/Q _5078_/S1 _5404_/A0 vssd1 vssd1 vccd1
+ vccd1 _4778_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_43_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3729_ _3714_/S _3717_/B _3726_/Y _3727_/Y vssd1 vssd1 vccd1 vccd1 _3886_/S sky130_fd_sc_hd__a31o_1
XANTENNA__4499__S _4500_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6448_ _6448_/CLK _6448_/D fanout185/X vssd1 vssd1 vccd1 vccd1 hold1/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6379_ _6465_/CLK _6379_/D vssd1 vssd1 vccd1 vccd1 _6379_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__5497__B2 _5415_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5249__A1 _6338_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3151__B _5315_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold620_A _6463_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3432__B1 _4325_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3983__A1 _6384_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_4_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6452_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5660__A1 _6334_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5099__S0 _5100_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5412__A1 _5757_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5750_ hold23/X _3948_/B _6104_/S vssd1 vssd1 vccd1 vccd1 hold24/A sky130_fd_sc_hd__mux2_1
XFILLER_0_29_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4701_ _6097_/A _4714_/S vssd1 vssd1 vccd1 vccd1 _4701_/Y sky130_fd_sc_hd__nor2_1
X_5681_ _6221_/Q _5721_/A2 _5721_/B1 _6114_/Q _5730_/C1 vssd1 vssd1 vccd1 vccd1 _5683_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_60_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4632_ _6463_/Q _4606_/X _4607_/X _6314_/Q vssd1 vssd1 vccd1 vccd1 _4632_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4901__A _5102_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4563_ hold476/X _6312_/Q _4575_/S vssd1 vssd1 vccd1 vccd1 _4563_/X sky130_fd_sc_hd__mux2_1
Xhold603 _6336_/Q vssd1 vssd1 vccd1 vccd1 hold603/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6427__RESET_B fanout172/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4923__B1 _6367_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold625 _6300_/Q vssd1 vssd1 vccd1 vccd1 hold625/X sky130_fd_sc_hd__dlygate4sd3_1
X_3514_ _3652_/B _3514_/B _4338_/B vssd1 vssd1 vccd1 vccd1 _3514_/X sky130_fd_sc_hd__or3_1
X_6302_ _6308_/CLK _6302_/D fanout185/X vssd1 vssd1 vccd1 vccd1 _6302_/Q sky130_fd_sc_hd__dfrtp_1
Xhold614 _5293_/X vssd1 vssd1 vccd1 vccd1 _6340_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold636 _6335_/Q vssd1 vssd1 vccd1 vccd1 hold636/X sky130_fd_sc_hd__buf_1
X_4494_ _4416_/X hold171/X _4500_/S vssd1 vssd1 vccd1 vccd1 _4494_/X sky130_fd_sc_hd__mux2_1
Xhold647 _6296_/Q vssd1 vssd1 vccd1 vccd1 hold647/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold658 _6150_/Q vssd1 vssd1 vccd1 vccd1 hold658/X sky130_fd_sc_hd__dlygate4sd3_1
X_3445_ _3258_/B _3685_/A _3673_/B vssd1 vssd1 vccd1 vccd1 _3449_/A sky130_fd_sc_hd__a21oi_1
X_6233_ _6456_/CLK _6233_/D vssd1 vssd1 vccd1 vccd1 _6233_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5732__A _5732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3376_ _5522_/A _3376_/B _4325_/C _4253_/A vssd1 vssd1 vccd1 vccd1 _3379_/C sky130_fd_sc_hd__and4_1
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6164_ _6470_/CLK _6167_/D fanout179/X vssd1 vssd1 vccd1 vccd1 _6164_/Q sky130_fd_sc_hd__dfstp_1
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6095_ _6101_/B _5063_/B _5577_/Y _6036_/X vssd1 vssd1 vccd1 vccd1 _6095_/X sky130_fd_sc_hd__o22a_1
X_5115_ _6409_/Q _5114_/X _6070_/A vssd1 vssd1 vccd1 vccd1 _5115_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5451__B _6461_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5046_ _6373_/Q _5047_/B vssd1 vssd1 vccd1 vccd1 _5086_/C sky130_fd_sc_hd__and2_1
XFILLER_0_33_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5878__S _5974_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4454__A2 _4462_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5651__A1 _6421_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5948_ _6463_/Q _5947_/X _5974_/S vssd1 vssd1 vccd1 vccd1 _5948_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_90_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5879_ _5878_/X hold518/X _6021_/S vssd1 vssd1 vccd1 vccd1 _5879_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4914__A0 _6366_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3427__A _5314_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4957__S _4957_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5642__A _5644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4692__S _4711_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3230_ _3230_/A vssd1 vssd1 vccd1 vccd1 _3230_/Y sky130_fd_sc_hd__inv_2
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3161_ _3240_/B _3161_/B vssd1 vssd1 vccd1 vccd1 _5371_/B sky130_fd_sc_hd__nor2_1
XANTENNA__4168__A _4332_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3072__A _5105_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3092_ _6312_/Q vssd1 vssd1 vccd1 vccd1 _3092_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_55_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3800__A _3884_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5802_ _5813_/A _5802_/B vssd1 vssd1 vccd1 vccd1 _5804_/B sky130_fd_sc_hd__or2_1
XANTENNA__4819__S0 _5078_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xci2406_z80_197 vssd1 vssd1 vccd1 vccd1 ci2406_z80_197/HI io_oeb[12] sky130_fd_sc_hd__conb_1
Xci2406_z80_186 vssd1 vssd1 vccd1 vccd1 ci2406_z80_186/HI io_oeb[0] sky130_fd_sc_hd__conb_1
X_3994_ _6085_/A vssd1 vssd1 vccd1 vccd1 _3994_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_29_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5733_ _5655_/B _4458_/X _5730_/X _5732_/X vssd1 vssd1 vccd1 vccd1 _5733_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_29_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5664_ _5757_/B _3081_/A _5611_/Y _5663_/X vssd1 vssd1 vccd1 vccd1 _5664_/X sky130_fd_sc_hd__a22o_1
X_4615_ _5393_/A1 hold564/X _4582_/Y _4614_/X vssd1 vssd1 vccd1 vccd1 _4615_/X sky130_fd_sc_hd__a22o_1
X_5595_ _5595_/A _5595_/B vssd1 vssd1 vccd1 vccd1 _5595_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_25_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold400 _5727_/X vssd1 vssd1 vccd1 vccd1 _6384_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold411 _6329_/Q vssd1 vssd1 vccd1 vccd1 hold411/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4546_ _4546_/A _4546_/B vssd1 vssd1 vccd1 vccd1 _4554_/S sky130_fd_sc_hd__or2_4
Xhold433 _3486_/X vssd1 vssd1 vccd1 vccd1 _6437_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold422 _5795_/X vssd1 vssd1 vccd1 vccd1 _6413_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold444 _6483_/Q vssd1 vssd1 vccd1 vccd1 hold444/X sky130_fd_sc_hd__buf_1
Xhold477 _4563_/X vssd1 vssd1 vccd1 vccd1 _6270_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold455 _4565_/X vssd1 vssd1 vccd1 vccd1 _6272_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold466 _6267_/Q vssd1 vssd1 vccd1 vccd1 hold466/X sky130_fd_sc_hd__dlygate4sd3_1
X_4477_ hold189/X _4428_/X _4482_/S vssd1 vssd1 vccd1 vccd1 _6188_/D sky130_fd_sc_hd__mux2_1
X_3428_ _4313_/A _3428_/B vssd1 vssd1 vccd1 vccd1 _3457_/B sky130_fd_sc_hd__nor2_1
Xhold488 _4630_/X vssd1 vssd1 vccd1 vccd1 _6288_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6216_ _6393_/CLK hold90/X vssd1 vssd1 vccd1 vccd1 hold89/A sky130_fd_sc_hd__dfxtp_1
Xhold499 _6064_/X vssd1 vssd1 vccd1 vccd1 _6480_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3359_ _3511_/A _3986_/A _4217_/A vssd1 vssd1 vccd1 vccd1 _4116_/A sky130_fd_sc_hd__and3b_2
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6147_ _6265_/CLK _6147_/D vssd1 vssd1 vccd1 vccd1 _6147_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6078_ _4366_/A _6075_/X _6076_/Y _6077_/Y hold444/X vssd1 vssd1 vccd1 vccd1 _6078_/X
+ sky130_fd_sc_hd__o32a_1
X_5029_ _6461_/Q _5028_/Y _5108_/S vssd1 vssd1 vccd1 vccd1 _5029_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_95_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6349__RESET_B fanout176/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5637__A _5732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3157__A _4268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4687__S _4712_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5615__A1 _4675_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4716__A _4716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5710__S1 _5734_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5394__A3 _5645_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4400_ _4400_/A _6003_/B vssd1 vssd1 vccd1 vccd1 _4464_/S sky130_fd_sc_hd__nor2_4
X_5380_ _5767_/A _5377_/Y _6021_/S vssd1 vssd1 vccd1 vccd1 _5380_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_22_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4331_ _5605_/A _5315_/A _5374_/B vssd1 vssd1 vccd1 vccd1 _5370_/D sky130_fd_sc_hd__and3_1
XFILLER_0_22_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4262_ _5364_/A _4262_/B vssd1 vssd1 vccd1 vccd1 _4328_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_1_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4657__A2 _4652_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3213_ _5605_/A _3281_/A _5360_/A _4595_/B vssd1 vssd1 vccd1 vccd1 _3213_/X sky130_fd_sc_hd__and4_1
X_6001_ _5384_/A _3469_/B hold1/X vssd1 vssd1 vccd1 vccd1 hold2/A sky130_fd_sc_hd__o21a_1
XFILLER_0_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6097__B _6107_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4193_ _5268_/A _4193_/B vssd1 vssd1 vccd1 vccd1 _4196_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_66_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3144_ _4782_/A _3172_/A _3284_/B vssd1 vssd1 vccd1 vccd1 _3281_/A sky130_fd_sc_hd__and3_2
XANTENNA__5606__A1 _5777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4409__A2 _4406_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3075_ _6347_/Q vssd1 vssd1 vccd1 vccd1 _5294_/A sky130_fd_sc_hd__inv_2
XANTENNA__5606__B2 _4595_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3530__A _3530_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_32_wb_clk_i_A clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__5082__A2 _4963_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4814__C1 _5102_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5241__A2_N _5292_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5909__A2 _5785_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3977_ _4156_/A _3975_/Y _3976_/X vssd1 vssd1 vccd1 vccd1 _3977_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_45_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4593__A1 _4675_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6442__RESET_B fanout181/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4361__A _6100_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5716_ _6339_/Q _5628_/X _5643_/X _6427_/Q vssd1 vssd1 vccd1 vccd1 _5726_/B sky130_fd_sc_hd__a22o_1
XANTENNA__5790__B1 _5867_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5647_ _6483_/Q _5653_/B _5645_/C vssd1 vssd1 vccd1 vccd1 _5647_/X sky130_fd_sc_hd__a21o_1
X_5578_ hold562/X _5520_/B _5577_/Y _5415_/X vssd1 vssd1 vccd1 vccd1 _5578_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_5_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold230 _6342_/Q vssd1 vssd1 vccd1 vccd1 hold230/X sky130_fd_sc_hd__dlygate4sd3_1
X_4529_ hold57/X _4404_/X _4536_/S vssd1 vssd1 vccd1 vccd1 hold58/A sky130_fd_sc_hd__mux2_1
XANTENNA__4896__A2 _5783_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold241 _4517_/X vssd1 vssd1 vccd1 vccd1 _6224_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold252 _6115_/Q vssd1 vssd1 vccd1 vccd1 hold252/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4440__S1 _5721_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold285 _6114_/Q vssd1 vssd1 vccd1 vccd1 hold285/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold263 _6175_/Q vssd1 vssd1 vccd1 vccd1 hold263/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6098__A1 _4366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold296 _6453_/Q vssd1 vssd1 vccd1 vccd1 hold296/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold274 _6410_/Q vssd1 vssd1 vccd1 vccd1 hold274/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5845__A1 _5887_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5845__B2 _5786_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4970__S _5108_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4033__B1 _3807_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4584__A1 _4276_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4336__A1 _4782_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5836__A1 _5867_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5117__C_N _4670_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput9 io_in[25] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_59_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5976__S _5976_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3152__A_N _5605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3709__C_N _4670_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4880_ _6206_/Q _6214_/Q _6453_/Q _6230_/Q _5100_/S0 _5100_/S1 vssd1 vssd1 vccd1
+ vccd1 _4880_/X sky130_fd_sc_hd__mux4_1
X_3900_ _4190_/A _4641_/A _3898_/A _4451_/C _4459_/A vssd1 vssd1 vccd1 vccd1 _3901_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_86_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3831_ _4190_/A _4636_/A vssd1 vssd1 vccd1 vccd1 _4459_/A sky130_fd_sc_hd__and2_1
X_3762_ _4168_/B vssd1 vssd1 vccd1 vccd1 _3762_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4575__A1 _6340_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4291__C_N _4768_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5772__B1 _3503_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5501_ hold590/X _5500_/X _5513_/S vssd1 vssd1 vccd1 vccd1 _5501_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_27_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3693_ _3693_/A _3693_/B _3693_/C vssd1 vssd1 vccd1 vccd1 _3693_/X sky130_fd_sc_hd__or3_2
X_6481_ _6481_/CLK _6481_/D fanout176/X vssd1 vssd1 vccd1 vccd1 _6481_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA__4327__A1 _5315_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5432_ _5432_/A _5432_/B vssd1 vssd1 vccd1 vccd1 _5433_/A sky130_fd_sc_hd__xnor2_1
X_5363_ hold655/X _3278_/A _4328_/A _4281_/A vssd1 vssd1 vccd1 vccd1 _5364_/C sky130_fd_sc_hd__a211o_1
XFILLER_0_2_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3525__A _5384_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4314_ _4313_/A _4319_/D _4319_/B vssd1 vssd1 vccd1 vccd1 _4315_/C sky130_fd_sc_hd__a21oi_1
XFILLER_0_10_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3244__B _3304_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5294_ _5294_/A _5294_/B vssd1 vssd1 vccd1 vccd1 _5294_/X sky130_fd_sc_hd__or2_1
XFILLER_0_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4245_ _5314_/S _4251_/B _3219_/A vssd1 vssd1 vccd1 vccd1 _5388_/B sky130_fd_sc_hd__o21a_1
X_4176_ _3083_/Y _4175_/Y _4227_/S vssd1 vssd1 vccd1 vccd1 _6067_/A sky130_fd_sc_hd__mux2_4
X_3127_ _5387_/A _4557_/C _3627_/B vssd1 vssd1 vccd1 vccd1 _3617_/A sky130_fd_sc_hd__or3_2
X_3058_ _3511_/A vssd1 vssd1 vccd1 vccd1 _5124_/A sky130_fd_sc_hd__inv_2
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4015__B1 _6334_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4091__A _6289_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4566__A1 _6315_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5763__A0 _6314_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6337__SET_B fanout183/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4318__A1 _4313_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4965__S _5105_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3829__B1 _3804_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3170__A _5344_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6364__RESET_B fanout181/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5809__B _5867_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3780__A2 _6458_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5036__S _6070_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4030_ _3734_/X _6089_/A _3700_/Y vssd1 vssd1 vccd1 vccd1 _4030_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__3080__A _6286_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5981_ _5995_/D _5988_/B _5995_/B vssd1 vssd1 vccd1 vccd1 _5981_/X sky130_fd_sc_hd__or3_1
XFILLER_0_63_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4932_ _4931_/X _6367_/Q _5861_/S vssd1 vssd1 vccd1 vccd1 _4932_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_59_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4863_ _4862_/X _4861_/X _5101_/S vssd1 vssd1 vccd1 vccd1 _4863_/X sky130_fd_sc_hd__mux2_2
X_4794_ _4802_/D _4802_/C _4802_/B vssd1 vssd1 vccd1 vccd1 _4794_/Y sky130_fd_sc_hd__nor3b_2
X_3814_ _4600_/A vssd1 vssd1 vccd1 vccd1 _3814_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_27_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3239__B _3632_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3745_ _6345_/Q _6333_/Q vssd1 vssd1 vccd1 vccd1 _3748_/S sky130_fd_sc_hd__and2b_1
XFILLER_0_6_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6464_ _6465_/CLK _6464_/D fanout181/X vssd1 vssd1 vccd1 vccd1 _6464_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_42_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3676_ _5406_/B _4267_/B _5777_/A _5387_/C vssd1 vssd1 vccd1 vccd1 _3676_/X sky130_fd_sc_hd__a211o_1
X_5415_ _6434_/Q _6469_/Q vssd1 vssd1 vccd1 vccd1 _5415_/X sky130_fd_sc_hd__and2_2
XFILLER_0_2_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout117_A _6108_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_28_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6417_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_6395_ _6490_/CLK hold24/X vssd1 vssd1 vccd1 vccd1 hold23/A sky130_fd_sc_hd__dfxtp_1
X_5346_ _5346_/A _5346_/B _5346_/C _5346_/D vssd1 vssd1 vccd1 vccd1 _5346_/X sky130_fd_sc_hd__or4_1
X_5277_ _5271_/X _5276_/X _5290_/S vssd1 vssd1 vccd1 vccd1 _5277_/X sky130_fd_sc_hd__mux2_1
X_4228_ _4414_/A _4227_/X _3701_/B vssd1 vssd1 vccd1 vccd1 _4228_/X sky130_fd_sc_hd__a21o_1
XANTENNA__3702__B _4150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5681__C1 _5730_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4159_ _5136_/A _6290_/Q _6384_/Q _4060_/B _4158_/X vssd1 vssd1 vccd1 vccd1 _5160_/A
+ sky130_fd_sc_hd__o41a_2
XFILLER_0_38_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5645__A _5645_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4711__A1 _6381_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4724__A _5605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput12 io_in[28] vssd1 vssd1 vccd1 vccd1 _4656_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_83_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3202__A1 _6430_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3530_ _3530_/A _3530_/B _3307_/B vssd1 vssd1 vccd1 vccd1 _3530_/X sky130_fd_sc_hd__or3b_1
XFILLER_0_24_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4950__B2 _6465_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3461_ hold45/X _3464_/B _3460_/X vssd1 vssd1 vccd1 vccd1 _3461_/X sky130_fd_sc_hd__a21o_1
X_3392_ _3497_/B _4335_/C _5369_/A _5369_/B vssd1 vssd1 vccd1 vccd1 _3393_/C sky130_fd_sc_hd__or4_1
XANTENNA__4702__A1 _6379_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5200_ _6382_/Q _4073_/A _5196_/X _5199_/X vssd1 vssd1 vccd1 vccd1 _5200_/X sky130_fd_sc_hd__a211o_1
X_6180_ _6263_/CLK _6180_/D vssd1 vssd1 vccd1 vccd1 _6180_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4804__B_N _5777_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5131_ _5288_/S _5132_/B vssd1 vssd1 vccd1 vccd1 _5131_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_58_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5062_ _5064_/B vssd1 vssd1 vccd1 vccd1 _5063_/B sky130_fd_sc_hd__inv_2
X_4013_ _6285_/Q _6286_/Q _6287_/Q _4107_/B vssd1 vssd1 vccd1 vccd1 _4013_/Y sky130_fd_sc_hd__a31oi_1
XFILLER_0_74_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5964_ _5964_/A _5964_/B vssd1 vssd1 vccd1 vccd1 _5964_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_90_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5895_ _4962_/Y _5894_/Y _5771_/A vssd1 vssd1 vccd1 vccd1 _5895_/Y sky130_fd_sc_hd__a21oi_1
X_4915_ _4319_/B _4914_/X _5016_/S vssd1 vssd1 vccd1 vccd1 _4915_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3992__A2 _6460_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4846_ _4844_/X _4845_/X _4948_/S vssd1 vssd1 vccd1 vccd1 _4846_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_35_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4777_ hold57/A hold65/A hold55/A hold87/A _5078_/S1 _5404_/A0 vssd1 vssd1 vccd1
+ vccd1 _4777_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_7_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3728_ _5295_/A _3711_/Y _5296_/A _4948_/S vssd1 vssd1 vccd1 vccd1 _3728_/X sky130_fd_sc_hd__a211o_1
XANTENNA__5795__A1_N _5977_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3659_ _6166_/Q _3657_/Y _3658_/X _6169_/Q vssd1 vssd1 vccd1 vccd1 _3659_/X sky130_fd_sc_hd__o22a_4
X_6447_ _6474_/CLK _6447_/D fanout179/X vssd1 vssd1 vccd1 vccd1 _6447_/Q sky130_fd_sc_hd__dfrtp_2
X_6378_ _6462_/CLK _6378_/D vssd1 vssd1 vccd1 vccd1 _6378_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__5497__A2 _5520_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5329_ _3219_/A _5360_/A _3428_/B vssd1 vssd1 vccd1 vccd1 _5329_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_11_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold613_A _6340_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_2_3__f_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4932__A1 _6367_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5822__B _5867_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5314__S _5314_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6109__2 _6439_/CLK vssd1 vssd1 vccd1 vccd1 _6166_/CLK sky130_fd_sc_hd__inv_2
XANTENNA__5948__A0 _6463_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5099__S1 _5100_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4700_ _4715_/B2 _4696_/Y _4699_/X hold320/X _4672_/Y vssd1 vssd1 vccd1 vccd1 _4700_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_0_29_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5680_ _5680_/A _5680_/B vssd1 vssd1 vccd1 vccd1 _5680_/X sky130_fd_sc_hd__or2_1
XANTENNA__4604__D _4641_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4631_ _3839_/B _4131_/B _4641_/B vssd1 vssd1 vccd1 vccd1 _4631_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4901__B _4901_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3726__A2 _3701_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4562_ hold462/X _6311_/Q _4575_/S vssd1 vssd1 vccd1 vccd1 _4562_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_8_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4923__A1 _6366_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold615 _6299_/Q vssd1 vssd1 vccd1 vccd1 hold615/X sky130_fd_sc_hd__dlygate4sd3_1
X_3513_ _6300_/Q _4248_/C _3333_/C _3986_/A vssd1 vssd1 vccd1 vccd1 _3513_/X sky130_fd_sc_hd__o2bb2a_1
X_6301_ _6340_/CLK _6301_/D fanout183/X vssd1 vssd1 vccd1 vccd1 _6301_/Q sky130_fd_sc_hd__dfrtp_1
Xhold604 _6161_/Q vssd1 vssd1 vccd1 vccd1 hold604/X sky130_fd_sc_hd__clkbuf_2
Xhold626 _6460_/Q vssd1 vssd1 vccd1 vccd1 hold626/X sky130_fd_sc_hd__dlygate4sd3_1
X_4493_ _4404_/X hold75/X _4500_/S vssd1 vssd1 vccd1 vccd1 hold76/A sky130_fd_sc_hd__mux2_1
Xhold648 _6297_/Q vssd1 vssd1 vccd1 vccd1 hold648/X sky130_fd_sc_hd__dlygate4sd3_1
X_3444_ _4325_/A _5777_/B vssd1 vssd1 vccd1 vccd1 _3444_/Y sky130_fd_sc_hd__nand2_1
Xhold659 _6440_/Q vssd1 vssd1 vccd1 vccd1 hold659/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold637 _6315_/Q vssd1 vssd1 vccd1 vccd1 hold637/X sky130_fd_sc_hd__dlygate4sd3_1
X_6232_ _6455_/CLK _6232_/D vssd1 vssd1 vccd1 vccd1 _6232_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4687__A0 _6384_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3375_ _3668_/A _5770_/B _3617_/A vssd1 vssd1 vccd1 vccd1 _3375_/X sky130_fd_sc_hd__a21o_1
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6163_ _6426_/CLK _6163_/D fanout171/X vssd1 vssd1 vccd1 vccd1 _6163_/Q sky130_fd_sc_hd__dfstp_1
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6094_ _4366_/A _6092_/X _6093_/Y hold535/X _6077_/Y vssd1 vssd1 vccd1 vccd1 _6094_/X
+ sky130_fd_sc_hd__o32a_1
X_5114_ _6465_/Q _5113_/X _5974_/S vssd1 vssd1 vccd1 vccd1 _5114_/X sky130_fd_sc_hd__mux2_1
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5045_ _5041_/B _5044_/X _5106_/S vssd1 vssd1 vccd1 vccd1 _5045_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_18_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5636__C1 _5730_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout184_A fanout185/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5947_ _5964_/A _5946_/X _5063_/Y vssd1 vssd1 vccd1 vccd1 _5947_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_63_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5878_ _6368_/Q _5877_/X _5974_/S vssd1 vssd1 vccd1 vccd1 _5878_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_62_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4829_ _6361_/Q _5108_/S _6362_/Q vssd1 vssd1 vccd1 vccd1 _4830_/B sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_43_wb_clk_i clkbuf_leaf_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6490_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_90_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3427__B _5360_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4678__A0 _6382_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5642__B _5734_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4142__A2 _3804_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3653__A1 _6023_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3337__B _3685_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6107__A0 _4227_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5044__S _5105_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3160_ _4247_/A _5345_/B vssd1 vssd1 vccd1 vccd1 _5369_/C sky130_fd_sc_hd__or2_1
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1 hold1/A vssd1 vssd1 vccd1 vccd1 hold1/X sky130_fd_sc_hd__clkbuf_2
X_3091_ _4303_/C vssd1 vssd1 vccd1 vccd1 _3091_/Y sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_22_wb_clk_i_A _6448_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5633__A2 _4406_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4398__C_N _4670_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4841__B1 _4789_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3800__B _3818_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5397__A1 _6434_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5801_ _5867_/B _5800_/C _6414_/Q vssd1 vssd1 vccd1 vccd1 _5802_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__4819__S1 _5404_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xci2406_z80_187 vssd1 vssd1 vccd1 vccd1 ci2406_z80_187/HI io_oeb[1] sky130_fd_sc_hd__conb_1
X_3993_ _3969_/B _3992_/Y _4227_/S vssd1 vssd1 vccd1 vccd1 _6085_/A sky130_fd_sc_hd__mux2_4
XFILLER_0_57_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xci2406_z80_198 vssd1 vssd1 vccd1 vccd1 ci2406_z80_198/HI io_oeb[13] sky130_fd_sc_hd__conb_1
X_5732_ _5732_/A _5732_/B vssd1 vssd1 vccd1 vccd1 _5732_/X sky130_fd_sc_hd__or2_1
XFILLER_0_84_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5149__A1 _6334_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5219__S _5292_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5663_ _5663_/A _5663_/B _5663_/C vssd1 vssd1 vccd1 vccd1 _5663_/X sky130_fd_sc_hd__or3_1
XFILLER_0_72_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5594_ _5594_/A _5594_/B vssd1 vssd1 vccd1 vccd1 _5595_/B sky130_fd_sc_hd__xor2_1
X_4614_ hold460/X _4604_/X _4605_/X hold520/X _4613_/X vssd1 vssd1 vccd1 vccd1 _4614_/X
+ sky130_fd_sc_hd__a221o_1
Xhold401 _6447_/Q vssd1 vssd1 vccd1 vccd1 _3373_/B sky130_fd_sc_hd__clkbuf_2
X_4545_ hold277/X _4463_/X _4545_/S vssd1 vssd1 vccd1 vccd1 _4545_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_40_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold434 _6274_/Q vssd1 vssd1 vccd1 vccd1 hold434/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold423 _6383_/Q vssd1 vssd1 vccd1 vccd1 _4087_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold412 _5057_/X vssd1 vssd1 vccd1 vccd1 _6329_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold445 _6078_/X vssd1 vssd1 vccd1 vccd1 _6483_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold478 _6439_/Q vssd1 vssd1 vccd1 vccd1 _5995_/B sky130_fd_sc_hd__clkbuf_2
Xhold467 _4560_/X vssd1 vssd1 vccd1 vccd1 _6267_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4476_ hold199/X _4416_/X _4482_/S vssd1 vssd1 vccd1 vccd1 _4476_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_13_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold456 _6403_/Q vssd1 vssd1 vccd1 vccd1 hold456/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3427_ _5314_/S _5360_/C vssd1 vssd1 vccd1 vccd1 _3428_/B sky130_fd_sc_hd__nor2_1
Xhold489 _6378_/Q vssd1 vssd1 vccd1 vccd1 hold489/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__4124__A2 _3793_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6215_ _6455_/CLK hold68/X vssd1 vssd1 vccd1 vccd1 hold67/A sky130_fd_sc_hd__dfxtp_1
X_3358_ _5605_/B _4716_/A vssd1 vssd1 vccd1 vccd1 _4720_/C sky130_fd_sc_hd__nand2b_2
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6146_ _6263_/CLK _6146_/D vssd1 vssd1 vccd1 vccd1 _6146_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3289_ _4335_/B _5777_/A vssd1 vssd1 vccd1 vccd1 _3674_/A sky130_fd_sc_hd__nor2_4
XANTENNA__5085__A0 _6101_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6077_ _6039_/Y _6107_/S _4366_/A vssd1 vssd1 vccd1 vccd1 _6077_/Y sky130_fd_sc_hd__a21oi_4
X_5028_ _5047_/B _5028_/B vssd1 vssd1 vccd1 vccd1 _5028_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_95_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold409_A _6332_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5312__A1 _5387_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5076__A0 _6407_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4716__B _5124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4330_ _3668_/A _5370_/B _5362_/A _5315_/A vssd1 vssd1 vccd1 vccd1 _4330_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_10_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4261_ _4261_/A _5145_/D vssd1 vssd1 vccd1 vccd1 _4261_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_10_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3212_ _5124_/A _5315_/A vssd1 vssd1 vccd1 vccd1 _3297_/B sky130_fd_sc_hd__nor2_2
X_6000_ _4653_/A _3638_/C _3650_/B vssd1 vssd1 vccd1 vccd1 _6000_/X sky130_fd_sc_hd__a21o_1
XANTENNA__5897__B1_N _5976_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4192_ _4155_/A _4155_/B _4157_/B vssd1 vssd1 vccd1 vccd1 _4193_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_66_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3143_ _3639_/C _3639_/D vssd1 vssd1 vccd1 vccd1 _5369_/A sky130_fd_sc_hd__nor2_2
X_3074_ _6436_/Q vssd1 vssd1 vccd1 vccd1 _3074_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_82_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3976_ _5136_/B _3971_/Y _3975_/A _3753_/X vssd1 vssd1 vccd1 vccd1 _3976_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_64_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4042__B2 _4441_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4361__B _4361_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5715_ _6481_/Q _5629_/X _5646_/X _6419_/Q vssd1 vssd1 vccd1 vccd1 _5726_/A sky130_fd_sc_hd__a22o_1
XANTENNA__5790__A1 _5866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5646_ _5644_/A _5646_/B _5734_/S vssd1 vssd1 vccd1 vccd1 _5646_/X sky130_fd_sc_hd__and3b_2
XFILLER_0_5_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5577_ _5577_/A vssd1 vssd1 vccd1 vccd1 _5577_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_13_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold220 _6259_/Q vssd1 vssd1 vccd1 vccd1 hold220/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold231 _5333_/X vssd1 vssd1 vccd1 vccd1 _6342_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold253 _6377_/Q vssd1 vssd1 vccd1 vccd1 _5601_/A sky130_fd_sc_hd__buf_1
X_4528_ _4528_/A _6003_/B vssd1 vssd1 vccd1 vccd1 _4536_/S sky130_fd_sc_hd__nor2_4
Xhold242 _6225_/Q vssd1 vssd1 vccd1 vccd1 hold242/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3705__B _4713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold286 _6253_/Q vssd1 vssd1 vccd1 vccd1 hold286/X sky130_fd_sc_hd__dlygate4sd3_1
X_4459_ _4459_/A _4459_/B vssd1 vssd1 vccd1 vccd1 _4460_/B sky130_fd_sc_hd__nor2_1
Xhold275 _5766_/X vssd1 vssd1 vccd1 vccd1 _6410_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold264 _6251_/Q vssd1 vssd1 vccd1 vccd1 hold264/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold297 _6222_/Q vssd1 vssd1 vccd1 vccd1 hold297/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6129_ _6481_/CLK _6129_/D vssd1 vssd1 vccd1 vccd1 _6129_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4584__A2 _4595_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3168__A _4782_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4698__S _4712_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5297__B1 _5757_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4272__A1 _4675_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4024__A1 _6381_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3830_ _3830_/A _3830_/B _3830_/C vssd1 vssd1 vccd1 vccd1 _4636_/A sky130_fd_sc_hd__or3_2
XFILLER_0_39_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3761_ _6343_/Q _3761_/B vssd1 vssd1 vccd1 vccd1 _4168_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_54_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5772__A1 _4957_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3078__A _4150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5500_ _6464_/Q _5499_/X _5512_/S vssd1 vssd1 vccd1 vccd1 _5500_/X sky130_fd_sc_hd__mux2_1
X_3692_ _4386_/A _3691_/X _3674_/A vssd1 vssd1 vccd1 vccd1 _3693_/C sky130_fd_sc_hd__a21oi_1
XFILLER_0_42_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6480_ _6480_/CLK _6480_/D fanout175/X vssd1 vssd1 vccd1 vccd1 _6480_/Q sky130_fd_sc_hd__dfstp_1
X_5431_ _5429_/X _5431_/B vssd1 vssd1 vccd1 vccd1 _5432_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_2_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5362_ _5362_/A _5388_/B _5362_/C _5362_/D vssd1 vssd1 vccd1 vccd1 _5362_/X sky130_fd_sc_hd__or4_1
XANTENNA__3597__A_N _5362_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4313_ _4313_/A _4319_/B _4319_/D vssd1 vssd1 vccd1 vccd1 _4315_/B sky130_fd_sc_hd__and3_1
XFILLER_0_2_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5293_ hold613/X _5292_/X _5489_/S vssd1 vssd1 vccd1 vccd1 _5293_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5288__A0 _6340_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4244_ _4244_/A vssd1 vssd1 vccd1 vccd1 _4244_/Y sky130_fd_sc_hd__inv_2
X_4175_ _5294_/A _6464_/Q _4174_/X vssd1 vssd1 vccd1 vccd1 _4175_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__5232__S _5232_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3126_ _5387_/A _4557_/C _3627_/B vssd1 vssd1 vccd1 vccd1 _5309_/A sky130_fd_sc_hd__nor3_4
X_3057_ _4217_/A vssd1 vssd1 vccd1 vccd1 _3057_/Y sky130_fd_sc_hd__inv_2
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3959_ _6220_/Q _3804_/X _3807_/X _6136_/Q vssd1 vssd1 vccd1 vccd1 _3959_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_18_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5515__A1 _4962_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5629_ _5644_/A _5653_/A _5734_/S vssd1 vssd1 vccd1 vccd1 _5629_/X sky130_fd_sc_hd__and3b_2
XFILLER_0_60_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5818__A2 _5771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold643_A _6333_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3170__B _4556_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4981__S _5101_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4254__A1 _4313_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3765__B1 _4595_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5754__A1 _4131_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3517__B1 _4324_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4245__A1 _5314_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5980_ _5980_/A _5995_/B vssd1 vssd1 vccd1 vccd1 _5980_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_86_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5993__A1 _5995_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4931_ _5892_/S _4929_/X _4930_/X _4921_/X vssd1 vssd1 vccd1 vccd1 _4931_/X sky130_fd_sc_hd__a31o_1
X_4862_ hold123/X _6213_/Q _6452_/Q _6229_/Q _5404_/A0 _5078_/S1 vssd1 vssd1 vccd1
+ vccd1 _4862_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_74_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3813_ _3813_/A _3813_/B vssd1 vssd1 vccd1 vccd1 _4600_/A sky130_fd_sc_hd__nand2_2
X_4793_ _4930_/B vssd1 vssd1 vccd1 vccd1 _4793_/Y sky130_fd_sc_hd__inv_4
XFILLER_0_6_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3744_ _6284_/Q _3744_/B vssd1 vssd1 vccd1 vccd1 _3750_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_82_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4920__A _5102_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3675_ _4344_/A _3673_/B _3674_/B _3674_/A _3557_/B vssd1 vssd1 vccd1 vccd1 _3675_/X
+ sky130_fd_sc_hd__o221a_2
X_6463_ _6465_/CLK _6463_/D fanout181/X vssd1 vssd1 vccd1 vccd1 _6463_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_88_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5414_ _5478_/S _5413_/Y _5432_/A vssd1 vssd1 vccd1 vccd1 _5414_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_88_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6394_ _6489_/CLK hold10/X vssd1 vssd1 vccd1 vccd1 hold9/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5345_ _5345_/A _5345_/B _5345_/C _5345_/D vssd1 vssd1 vccd1 vccd1 _5346_/D sky130_fd_sc_hd__or4_1
XFILLER_0_56_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5276_ _6409_/Q _4723_/X _5275_/X _5273_/Y vssd1 vssd1 vccd1 vccd1 _5276_/X sky130_fd_sc_hd__o31a_1
X_4227_ hold419/X _4226_/X _4227_/S vssd1 vssd1 vccd1 vccd1 _4227_/X sky130_fd_sc_hd__mux2_4
XANTENNA__5681__B1 _5721_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4158_ _3753_/X _4155_/A _4157_/X _5136_/B _4156_/Y vssd1 vssd1 vccd1 vccd1 _4158_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_69_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4089_ _5136_/A _6383_/Q vssd1 vssd1 vccd1 vccd1 _4091_/C sky130_fd_sc_hd__and2_1
X_3109_ _4782_/B _5605_/A _3547_/C vssd1 vssd1 vccd1 vccd1 _3652_/B sky130_fd_sc_hd__and3_2
XFILLER_0_77_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5629__C _5734_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5736__B2 _6465_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4976__S _5974_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5424__B1 _4300_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4724__B _6469_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6479__SET_B fanout176/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5727__A1 _4300_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput13 io_in[29] vssd1 vssd1 vccd1 vccd1 _4650_/A sky130_fd_sc_hd__buf_2
XFILLER_0_12_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3460_ _3464_/B _3464_/D _5478_/S vssd1 vssd1 vccd1 vccd1 _3460_/X sky130_fd_sc_hd__and3b_1
XFILLER_0_12_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3391_ _5109_/A1 _3388_/X _4948_/S _3072_/Y vssd1 vssd1 vccd1 vccd1 _4800_/S sky130_fd_sc_hd__o211a_4
XFILLER_0_20_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4886__S _5105_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5130_ _6021_/S _5783_/A vssd1 vssd1 vccd1 vccd1 _5786_/A sky130_fd_sc_hd__or2_2
X_5061_ _5101_/S _5060_/X _5059_/Y vssd1 vssd1 vccd1 vccd1 _5064_/B sky130_fd_sc_hd__o21ai_4
X_4012_ _6285_/Q _6286_/Q _6287_/Q vssd1 vssd1 vccd1 vccd1 _4107_/C sky130_fd_sc_hd__a21o_1
XANTENNA__3522__C _6442_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4218__A1 _5605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5963_ _6375_/Q _5848_/S _5972_/B1 _5962_/X vssd1 vssd1 vccd1 vccd1 _5964_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_87_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5966__B2 _5976_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4914_ _6366_/Q _4913_/X _5863_/S vssd1 vssd1 vccd1 vccd1 _4914_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_90_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5894_ _5964_/A _5894_/B vssd1 vssd1 vccd1 vccd1 _5894_/Y sky130_fd_sc_hd__nand2_1
X_4845_ _6415_/Q _6363_/Q _5105_/S vssd1 vssd1 vccd1 vccd1 _4845_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4650__A _4650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4776_ _5866_/A _4774_/Y _3644_/C vssd1 vssd1 vccd1 vccd1 _4776_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_55_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3727_ _5295_/A _3711_/Y _5296_/A _4948_/S vssd1 vssd1 vccd1 vccd1 _3727_/Y sky130_fd_sc_hd__a211oi_2
XFILLER_0_7_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6446_ _6446_/CLK _6446_/D fanout185/X vssd1 vssd1 vccd1 vccd1 _6446_/Q sky130_fd_sc_hd__dfrtp_1
X_3658_ input3/X input2/X vssd1 vssd1 vccd1 vccd1 _3658_/X sky130_fd_sc_hd__and2b_1
X_3589_ _5317_/A _5387_/C vssd1 vssd1 vccd1 vccd1 _4281_/A sky130_fd_sc_hd__nor2_1
X_6377_ _6377_/CLK _6377_/D fanout176/X vssd1 vssd1 vccd1 vccd1 _6377_/Q sky130_fd_sc_hd__dfrtp_1
X_5328_ _3221_/C _5350_/A _4217_/A _4313_/A vssd1 vssd1 vccd1 vccd1 _5328_/X sky130_fd_sc_hd__o2bb2a_1
XANTENNA__4809__B _5108_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5259_ _3368_/S _6354_/Q _5258_/X _6346_/Q vssd1 vssd1 vccd1 vccd1 _5259_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_97_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xwire92 wire92/A vssd1 vssd1 vccd1 vccd1 wire92/X sky130_fd_sc_hd__buf_2
XFILLER_0_65_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4448__B2 _4441_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_12_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_88_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3408__C1 _3632_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3959__B1 _3807_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4620__B2 _4619_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4630_ _5393_/A1 hold487/X _4582_/Y _4629_/X vssd1 vssd1 vccd1 vccd1 _4630_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_56_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6300_ _6446_/CLK _6300_/D fanout184/X vssd1 vssd1 vccd1 vccd1 _6300_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_52_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4561_ hold436/X _6310_/Q _4575_/S vssd1 vssd1 vccd1 vccd1 _4561_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3086__A _6458_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold605 _5353_/X vssd1 vssd1 vccd1 vccd1 hold605/X sky130_fd_sc_hd__dlygate4sd3_1
X_3512_ _4276_/A _3512_/B _3512_/C vssd1 vssd1 vccd1 vccd1 _3541_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_69_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold627 _6464_/Q vssd1 vssd1 vccd1 vccd1 hold627/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold616 _6458_/Q vssd1 vssd1 vccd1 vccd1 hold616/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4492_ _4546_/B _6003_/B vssd1 vssd1 vccd1 vccd1 _4500_/S sky130_fd_sc_hd__or2_4
Xhold649 _6293_/Q vssd1 vssd1 vccd1 vccd1 hold649/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3443_ _5145_/A _3443_/B vssd1 vssd1 vccd1 vccd1 _5777_/B sky130_fd_sc_hd__nand2_4
Xhold638 _6429_/Q vssd1 vssd1 vccd1 vccd1 hold638/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4136__B1 _4463_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6231_ _6454_/CLK _6231_/D vssd1 vssd1 vccd1 vccd1 _6231_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6162_ _6377_/CLK _6162_/D fanout179/X vssd1 vssd1 vccd1 vccd1 _6162_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3374_ _5770_/B vssd1 vssd1 vccd1 vccd1 _3374_/Y sky130_fd_sc_hd__inv_2
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5113_ _5964_/A _5112_/X _5102_/Y vssd1 vssd1 vccd1 vccd1 _5113_/X sky130_fd_sc_hd__a21bo_1
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6093_ _6093_/A _6107_/S vssd1 vssd1 vccd1 vccd1 _6093_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__4439__B2 _4462_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5044_ _6425_/Q _6373_/Q _5105_/S vssd1 vssd1 vccd1 vccd1 _5044_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_79_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout177_A fanout180/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5946_ _6374_/Q _5848_/S _5972_/B1 _5945_/X vssd1 vssd1 vccd1 vccd1 _5946_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_34_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5877_ _5964_/A _5876_/X _4942_/Y vssd1 vssd1 vccd1 vccd1 _5877_/X sky130_fd_sc_hd__a21bo_1
X_4828_ _6361_/Q _6362_/Q _5108_/S vssd1 vssd1 vccd1 vccd1 _4847_/B sky130_fd_sc_hd__and3_1
XFILLER_0_90_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4759_ hold639/X _4758_/X _5232_/S vssd1 vssd1 vccd1 vccd1 _6314_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_7_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6429_ _6444_/CLK _6429_/D fanout178/X vssd1 vssd1 vccd1 vccd1 _6429_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA__4127__B1 _3810_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_12_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6248_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__5875__A0 _6368_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold389_A _6434_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6100__A _6100_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4555__A _6159_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4290__A _5124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_max_cap91_A wire92/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2 hold2/A vssd1 vssd1 vccd1 vccd1 hold2/X sky130_fd_sc_hd__dlygate4sd3_1
X_3090_ _6309_/Q vssd1 vssd1 vccd1 vccd1 _3090_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_55_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5094__A1 _5102_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3992_ _5294_/A _6460_/Q _3991_/X vssd1 vssd1 vccd1 vccd1 _3992_/Y sky130_fd_sc_hd__a21oi_1
X_5800_ _6414_/Q _5867_/B _5800_/C vssd1 vssd1 vccd1 vccd1 _5813_/A sky130_fd_sc_hd__and3_1
Xci2406_z80_188 vssd1 vssd1 vccd1 vccd1 ci2406_z80_188/HI io_oeb[2] sky130_fd_sc_hd__conb_1
Xci2406_z80_199 vssd1 vssd1 vccd1 vccd1 ci2406_z80_199/HI io_oeb[14] sky130_fd_sc_hd__conb_1
X_5731_ _6177_/Q _4406_/B _4420_/S _6256_/Q _5731_/C1 vssd1 vssd1 vccd1 vccd1 _5732_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_57_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5662_ _6310_/Q _5630_/X _5646_/X _6414_/Q vssd1 vssd1 vccd1 vccd1 _5663_/C sky130_fd_sc_hd__a22o_1
X_5593_ _6490_/Q _5102_/B _5593_/S vssd1 vssd1 vccd1 vccd1 _5594_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4613_ _6459_/Q _4606_/X _4607_/X _6310_/Q _4612_/X vssd1 vssd1 vccd1 vccd1 _4613_/X
+ sky130_fd_sc_hd__a221o_1
Xhold402 _4647_/X vssd1 vssd1 vccd1 vccd1 _6292_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4544_ hold71/X _4456_/X _4545_/S vssd1 vssd1 vccd1 vccd1 hold72/A sky130_fd_sc_hd__mux2_1
Xhold424 _5714_/X vssd1 vssd1 vccd1 vccd1 _6383_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold435 _4567_/X vssd1 vssd1 vccd1 vccd1 _6274_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold413 _6349_/Q vssd1 vssd1 vccd1 vccd1 _6033_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_96_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold446 _6282_/Q vssd1 vssd1 vccd1 vccd1 hold446/X sky130_fd_sc_hd__dlygate4sd3_1
X_4475_ hold55/X _4404_/X _4482_/S vssd1 vssd1 vccd1 vccd1 hold56/A sky130_fd_sc_hd__mux2_1
Xhold468 _6488_/Q vssd1 vssd1 vccd1 vccd1 hold468/X sky130_fd_sc_hd__dlygate4sd3_1
X_6214_ _6454_/CLK _6214_/D vssd1 vssd1 vccd1 vccd1 _6214_/Q sky130_fd_sc_hd__dfxtp_1
Xhold457 _5759_/X vssd1 vssd1 vccd1 vccd1 _6403_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3426_ _4335_/B _3426_/B vssd1 vssd1 vccd1 vccd1 _5360_/C sky130_fd_sc_hd__nand2_2
Xhold479 _5998_/X vssd1 vssd1 vccd1 vccd1 hold479/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3357_ _4217_/A _4268_/A _5315_/A vssd1 vssd1 vccd1 vccd1 _4022_/B sky130_fd_sc_hd__and3_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6145_ _6239_/CLK _6145_/D vssd1 vssd1 vccd1 vccd1 _6145_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6076_ _6076_/A _6107_/S vssd1 vssd1 vccd1 vccd1 _6076_/Y sky130_fd_sc_hd__nor2_1
X_3288_ _3587_/B _5317_/B _3285_/Y vssd1 vssd1 vccd1 vccd1 _3288_/X sky130_fd_sc_hd__o21a_1
X_5027_ _6371_/Q _5026_/C _6372_/Q vssd1 vssd1 vccd1 vccd1 _5028_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_67_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6034__B1 _5418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5929_ _5928_/X _5922_/A _6021_/S vssd1 vssd1 vccd1 vccd1 _5929_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_0_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4716__C _6159_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3626__A2 _5757_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4823__A1 _5101_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3629__A _4325_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4434__S0 _5731_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5055__S _5974_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4260_ _4338_/A _4260_/B _4325_/C vssd1 vssd1 vccd1 vccd1 _5145_/D sky130_fd_sc_hd__or3_1
XFILLER_0_5_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3211_ _3323_/A _3211_/B _3326_/A _3514_/B vssd1 vssd1 vccd1 vccd1 _3352_/B sky130_fd_sc_hd__or4_4
X_4191_ _4191_/A _4191_/B vssd1 vssd1 vccd1 vccd1 _5304_/C sky130_fd_sc_hd__xnor2_1
X_3142_ _3497_/B _4358_/B vssd1 vssd1 vccd1 vccd1 _5371_/A sky130_fd_sc_hd__or2_1
X_3073_ _6025_/A vssd1 vssd1 vccd1 vccd1 _3464_/A sky130_fd_sc_hd__inv_2
XANTENNA__6016__A0 input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3975_ _3975_/A _3975_/B vssd1 vssd1 vccd1 vccd1 _3975_/Y sky130_fd_sc_hd__xnor2_1
X_5714_ _4300_/A _4087_/A _5611_/Y _5713_/X vssd1 vssd1 vccd1 vccd1 _5714_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_72_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5645_ _5645_/A _5645_/B _5645_/C vssd1 vssd1 vccd1 vccd1 _5645_/X sky130_fd_sc_hd__and3_2
XFILLER_0_86_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3553__A1 _3525_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold210 _5305_/X vssd1 vssd1 vccd1 vccd1 _6341_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5576_ _5576_/A _5576_/B vssd1 vssd1 vccd1 vccd1 _5577_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_13_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold232 _6112_/Q vssd1 vssd1 vccd1 vccd1 hold232/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold221 _4547_/X vssd1 vssd1 vccd1 vccd1 _6259_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold243 _4518_/X vssd1 vssd1 vccd1 vccd1 _6225_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4527_ _4463_/X hold290/X _4527_/S vssd1 vssd1 vccd1 vccd1 _6233_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_40_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4089__B _6383_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold254 _5601_/X vssd1 vssd1 vccd1 vccd1 _6377_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold287 _6113_/Q vssd1 vssd1 vccd1 vccd1 hold287/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold276 _6194_/Q vssd1 vssd1 vccd1 vccd1 hold276/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold265 _6254_/Q vssd1 vssd1 vccd1 vccd1 hold265/X sky130_fd_sc_hd__dlygate4sd3_1
X_4458_ hold284/X hold215/X hold255/X hold61/X _5731_/C1 _4420_/S vssd1 vssd1 vccd1
+ vccd1 _4458_/X sky130_fd_sc_hd__mux4_1
X_3409_ _3786_/A _5522_/D vssd1 vssd1 vccd1 vccd1 _3409_/Y sky130_fd_sc_hd__nor2_1
Xhold298 _6292_/Q vssd1 vssd1 vccd1 vccd1 hold298/X sky130_fd_sc_hd__buf_1
X_6128_ _6481_/CLK _6128_/D vssd1 vssd1 vccd1 vccd1 _6128_/Q sky130_fd_sc_hd__dfxtp_1
X_4389_ _4546_/A _4528_/A vssd1 vssd1 vccd1 vccd1 _4397_/S sky130_fd_sc_hd__nor2_4
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6059_ _6093_/A _6071_/S vssd1 vssd1 vccd1 vccd1 _6059_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_95_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4033__A2 _3804_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3168__B _3168_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3883__S _3883_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3184__A _5315_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5049__A1 _6462_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3760_ _4217_/A _4557_/C vssd1 vssd1 vccd1 vccd1 _3760_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_6_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3691_ _4338_/A _3691_/B vssd1 vssd1 vccd1 vccd1 _3691_/X sky130_fd_sc_hd__or2_1
X_5430_ _5492_/A _5429_/B _5429_/C vssd1 vssd1 vccd1 vccd1 _5431_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_42_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3535__A1 _3205_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5361_ _5359_/X _5360_/Y hold604/X vssd1 vssd1 vccd1 vccd1 _5391_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_2_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3806__B _3885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5292_ _4227_/X _5291_/X _5292_/S vssd1 vssd1 vccd1 vccd1 _5292_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_2_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4312_ _4312_/A _4312_/B _5418_/A _4312_/D vssd1 vssd1 vccd1 vccd1 _4319_/D sky130_fd_sc_hd__and4_1
X_4243_ _5388_/A _3296_/Y _4261_/A _5322_/A vssd1 vssd1 vccd1 vccd1 _4244_/A sky130_fd_sc_hd__a31o_1
XFILLER_0_10_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3299__B1 _4248_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4174_ _3738_/X _5160_/A _4173_/X _6347_/Q vssd1 vssd1 vccd1 vccd1 _4174_/X sky130_fd_sc_hd__o211a_1
X_3125_ _3323_/A _3168_/B _3229_/A _3205_/B vssd1 vssd1 vccd1 vccd1 _3627_/B sky130_fd_sc_hd__or4_4
X_3056_ _3229_/A vssd1 vssd1 vccd1 vccd1 _3326_/A sky130_fd_sc_hd__inv_2
XFILLER_0_96_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5460__A1 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4653__A _4653_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3958_ _6261_/Q _3793_/X _3795_/X _6196_/Q _3957_/X vssd1 vssd1 vccd1 vccd1 _3961_/A
+ sky130_fd_sc_hd__a221o_1
X_3889_ _3816_/B _3883_/X _3885_/Y _3887_/Y vssd1 vssd1 vccd1 vccd1 _5299_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_33_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5628_ _5644_/A _5653_/A _5630_/D vssd1 vssd1 vccd1 vccd1 _5628_/X sky130_fd_sc_hd__and3_2
XANTENNA__3526__B2 _3525_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3526__A1 _5384_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5559_ _6487_/Q _5041_/B _5593_/S vssd1 vssd1 vccd1 vccd1 _5561_/B sky130_fd_sc_hd__mux2_1
XANTENNA__3829__A2 _3731_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3732__A _3852_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4254__A2 _5387_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold636_A _6335_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3179__A _3304_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4411__C1 _5655_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4502__S _4509_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4714__A0 _4227_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6373__RESET_B fanout172/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6302__RESET_B fanout185/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5690__A1 _6337_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5690__B2 _6425_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_13 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5442__A1 _5492_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4930_ _6419_/Q _4930_/B vssd1 vssd1 vccd1 vccd1 _4930_/X sky130_fd_sc_hd__or2_1
XFILLER_0_47_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4861_ hold151/X hold81/X _6173_/Q hold206/X _5404_/A0 _5078_/S1 vssd1 vssd1 vccd1
+ vccd1 _4861_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_86_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3812_ _6111_/Q _4519_/A _4537_/A _6178_/Q _3809_/X vssd1 vssd1 vccd1 vccd1 _3813_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_27_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4792_ _4792_/A _4802_/C _4802_/D vssd1 vssd1 vccd1 vccd1 _4930_/B sky130_fd_sc_hd__or3b_4
XANTENNA__4953__A0 _6368_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3743_ _4150_/A _3743_/B vssd1 vssd1 vccd1 vccd1 _3743_/X sky130_fd_sc_hd__or2_1
XFILLER_0_12_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4920__B _4920_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3674_ _3674_/A _3674_/B vssd1 vssd1 vccd1 vccd1 _5603_/C sky130_fd_sc_hd__nor2_1
X_6462_ _6462_/CLK _6462_/D fanout181/X vssd1 vssd1 vccd1 vccd1 _6462_/Q sky130_fd_sc_hd__dfrtp_4
X_5413_ _6458_/Q _5413_/B vssd1 vssd1 vccd1 vccd1 _5413_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_42_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6393_ _6393_/CLK hold14/X vssd1 vssd1 vccd1 vccd1 hold13/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5344_ _5369_/A _5344_/B _4344_/A vssd1 vssd1 vccd1 vccd1 _5345_/D sky130_fd_sc_hd__or3b_1
XFILLER_0_88_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5275_ _6407_/Q _6406_/Q _6408_/Q _5275_/D vssd1 vssd1 vccd1 vccd1 _5275_/X sky130_fd_sc_hd__or4_1
X_4226_ _6465_/Q _4225_/X _4226_/S vssd1 vssd1 vccd1 vccd1 _4226_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_49_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4157_ _6344_/Q _4157_/B vssd1 vssd1 vccd1 vccd1 _4157_/X sky130_fd_sc_hd__or2_1
X_3108_ _3323_/A _3211_/B vssd1 vssd1 vccd1 vccd1 _3229_/C sky130_fd_sc_hd__nand2_2
XANTENNA__3692__B1 _3674_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4088_ _5136_/A _6383_/Q vssd1 vssd1 vccd1 vccd1 _4091_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_78_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4236__A2 _4406_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5479__A _5492_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_37_wb_clk_i clkbuf_leaf_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6488_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_93_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3446__B _5777_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4172__A1 _4332_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4172__B2 _6384_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold586_A _6423_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4558__A wire92/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5672__A1 _6311_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3683__B1 _5607_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5424__A1 _4957_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5188__B1 _5600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput14 io_in[30] vssd1 vssd1 vccd1 vccd1 _6445_/D sky130_fd_sc_hd__buf_1
XANTENNA__3202__A3 _4248_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3356__B _6333_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_41_wb_clk_i_A clkbuf_leaf_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_3390_ _6359_/Q _3390_/B vssd1 vssd1 vccd1 vccd1 _3390_/X sky130_fd_sc_hd__or2_2
XFILLER_0_20_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5060_ _6264_/Q _6199_/Q _6223_/Q _6116_/Q _5100_/S0 _5100_/S1 vssd1 vssd1 vccd1
+ vccd1 _5060_/X sky130_fd_sc_hd__mux4_2
XFILLER_0_20_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4011_ _4199_/A _6287_/Q _6381_/Q _4060_/B _4010_/X vssd1 vssd1 vccd1 vccd1 _5256_/B
+ sky130_fd_sc_hd__o41a_2
XANTENNA__4218__A2 _6290_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5962_ _6408_/Q _6427_/Q _5971_/S vssd1 vssd1 vccd1 vccd1 _5962_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5966__A2 _5786_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4913_ _5817_/A _4912_/X _4901_/Y vssd1 vssd1 vccd1 vccd1 _4913_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_90_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5893_ _6369_/Q _5861_/S _5972_/B1 _5892_/X vssd1 vssd1 vccd1 vccd1 _5894_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_62_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5718__A2 _6355_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4844_ _4843_/X _4842_/X _5101_/S vssd1 vssd1 vccd1 vccd1 _4844_/X sky130_fd_sc_hd__mux2_2
XANTENNA__4650__B _4668_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4775_ _5866_/A _4774_/Y _3644_/C vssd1 vssd1 vccd1 vccd1 _5863_/S sky130_fd_sc_hd__o21a_4
XFILLER_0_7_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4926__A0 _4920_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3726_ hold41/A _3701_/B _4463_/S vssd1 vssd1 vccd1 vccd1 _3726_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_70_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6445_ _6446_/CLK _6445_/D fanout184/X vssd1 vssd1 vccd1 vccd1 _6445_/Q sky130_fd_sc_hd__dfrtp_1
X_3657_ input2/X input3/X vssd1 vssd1 vccd1 vccd1 _3657_/Y sky130_fd_sc_hd__nor2_1
X_3588_ _4276_/A _4676_/A vssd1 vssd1 vccd1 vccd1 _3588_/Y sky130_fd_sc_hd__nand2_1
X_6376_ _6376_/CLK _6376_/D fanout172/X vssd1 vssd1 vccd1 vccd1 _6376_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_2_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5327_ _5327_/A _5327_/B _5327_/C _5327_/D vssd1 vssd1 vccd1 vccd1 _5350_/A sky130_fd_sc_hd__and4_1
XFILLER_0_2_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6485__SET_B fanout172/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5258_ _5160_/A _5160_/B _5257_/X _5284_/S vssd1 vssd1 vccd1 vccd1 _5258_/X sky130_fd_sc_hd__o31a_1
XANTENNA__5654__B2 _6459_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5654__A1 _6422_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5189_ _5866_/A _6335_/Q _5187_/Y _5188_/X vssd1 vssd1 vccd1 vccd1 _5189_/X sky130_fd_sc_hd__o22a_1
X_4209_ _4209_/A _4209_/B vssd1 vssd1 vccd1 vccd1 _4211_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_3_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4317__S _5232_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5002__A _5102_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4090__B1 _6289_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5590__A0 _6464_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4288__A _4289_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout180 input18/X vssd1 vssd1 vccd1 vccd1 fanout180/X sky130_fd_sc_hd__buf_4
XFILLER_0_88_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_8_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__4081__B1 _4462_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4560_ hold466/X _6309_/Q _4575_/S vssd1 vssd1 vccd1 vccd1 _4560_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_4_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold606 _5354_/X vssd1 vssd1 vccd1 vccd1 _6344_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3511_ _3511_/A _3511_/B vssd1 vssd1 vccd1 vccd1 _3512_/C sky130_fd_sc_hd__nand2_1
Xhold617 _6347_/Q vssd1 vssd1 vccd1 vccd1 hold617/X sky130_fd_sc_hd__buf_1
X_4491_ _4240_/X hold167/X _4491_/S vssd1 vssd1 vccd1 vccd1 _4491_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_100_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3442_ _3489_/B _3477_/A vssd1 vssd1 vccd1 vccd1 _3443_/B sky130_fd_sc_hd__nor2_1
Xhold628 _6465_/Q vssd1 vssd1 vccd1 vccd1 hold628/X sky130_fd_sc_hd__buf_1
Xhold639 _6314_/Q vssd1 vssd1 vccd1 vccd1 hold639/X sky130_fd_sc_hd__dlygate4sd3_1
X_6230_ _6454_/CLK _6230_/D vssd1 vssd1 vccd1 vccd1 _6230_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4198__A _5268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3373_ _6442_/Q _3373_/B vssd1 vssd1 vccd1 vccd1 _5770_/B sky130_fd_sc_hd__or2_4
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6161_ _6470_/CLK _6161_/D fanout179/X vssd1 vssd1 vccd1 vccd1 _6161_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5112_ _6376_/Q _5848_/S _5972_/B1 _5111_/X vssd1 vssd1 vccd1 vccd1 _5112_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_20_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6092_ _6101_/A _6091_/X _6107_/S vssd1 vssd1 vccd1 vccd1 _6092_/X sky130_fd_sc_hd__o21a_1
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5043_ _6487_/Q _5104_/A2 _5042_/X vssd1 vssd1 vccd1 vccd1 _5043_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_18_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6061__B2 _6036_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6061__A1 _6101_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5945_ _6407_/Q _6426_/Q _5971_/S vssd1 vssd1 vccd1 vccd1 _5945_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5757__A _5757_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5876_ _6368_/Q _5861_/S _5972_/B1 _5875_/X vssd1 vssd1 vccd1 vccd1 _5876_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_90_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4827_ _4822_/X _4826_/X _4948_/S vssd1 vssd1 vccd1 vccd1 _4827_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_47_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4758_ _4122_/Y _4757_/X _4770_/S vssd1 vssd1 vccd1 vccd1 _4758_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_43_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4689_ _4713_/A _4687_/X _4714_/S vssd1 vssd1 vccd1 vccd1 _4689_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_70_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3709_ _3709_/A _4398_/B _4670_/C vssd1 vssd1 vccd1 vccd1 _3709_/X sky130_fd_sc_hd__or3b_1
XANTENNA__5492__A _5492_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6428_ _6428_/CLK _6428_/D fanout172/X vssd1 vssd1 vccd1 vccd1 _6428_/Q sky130_fd_sc_hd__dfrtp_2
X_6359_ _6377_/CLK _6359_/D fanout179/X vssd1 vssd1 vccd1 vccd1 _6359_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_0_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4555__B _4556_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6052__A1 _4366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4290__B _5478_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4118__B2 _6383_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4669__A2 _4652_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3 hold3/A vssd1 vssd1 vccd1 vccd1 hold3/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3237__D_N _4268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4841__A2 _4790_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3991_ _6347_/Q _3991_/B _3991_/C vssd1 vssd1 vccd1 vccd1 _3991_/X sky130_fd_sc_hd__and3_1
XFILLER_0_29_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xci2406_z80_189 vssd1 vssd1 vccd1 vccd1 ci2406_z80_189/HI io_oeb[3] sky130_fd_sc_hd__conb_1
X_5730_ _6456_/Q _4406_/B _4420_/S _6233_/Q _5730_/C1 vssd1 vssd1 vccd1 vccd1 _5730_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_72_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5661_ _6476_/Q _5629_/X _5632_/Y _5659_/X vssd1 vssd1 vccd1 vccd1 _5663_/B sky130_fd_sc_hd__a22o_1
X_5592_ _5587_/A _5587_/B _5585_/A vssd1 vssd1 vccd1 vccd1 _5595_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_25_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4612_ _3948_/B _4611_/B _4602_/Y _4611_/Y vssd1 vssd1 vccd1 vccd1 _4612_/X sky130_fd_sc_hd__o211a_1
X_4543_ hold265/X _4448_/X _4545_/S vssd1 vssd1 vccd1 vccd1 _6254_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_20_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold425 _6379_/Q vssd1 vssd1 vccd1 vccd1 _3081_/A sky130_fd_sc_hd__buf_1
Xhold414 _5379_/X vssd1 vssd1 vccd1 vccd1 _6349_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold436 _6268_/Q vssd1 vssd1 vccd1 vccd1 hold436/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold403 _6404_/Q vssd1 vssd1 vccd1 vccd1 hold403/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold447 _4575_/X vssd1 vssd1 vccd1 vccd1 _6282_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold458 _6271_/Q vssd1 vssd1 vccd1 vccd1 hold458/X sky130_fd_sc_hd__dlygate4sd3_1
X_6213_ _6452_/CLK _6213_/D vssd1 vssd1 vccd1 vccd1 _6213_/Q sky130_fd_sc_hd__dfxtp_1
X_4474_ _4474_/A _6003_/B vssd1 vssd1 vccd1 vccd1 _4482_/S sky130_fd_sc_hd__nor2_4
Xhold469 _6098_/X vssd1 vssd1 vccd1 vccd1 _6488_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3425_ _3786_/A _3421_/Y _5146_/C vssd1 vssd1 vccd1 vccd1 _3425_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3356_ _4217_/A _6333_/Q vssd1 vssd1 vccd1 vccd1 _3511_/B sky130_fd_sc_hd__xnor2_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6144_ _6263_/CLK hold96/X vssd1 vssd1 vccd1 vccd1 hold95/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__4656__A _4656_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3287_ _4276_/A _3489_/B vssd1 vssd1 vccd1 vccd1 _5317_/B sky130_fd_sc_hd__or2_4
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6075_ _6101_/A _6074_/X _6107_/S vssd1 vssd1 vccd1 vccd1 _6075_/X sky130_fd_sc_hd__o21a_1
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5026_ _6371_/Q _6372_/Q _5026_/C vssd1 vssd1 vccd1 vccd1 _5047_/B sky130_fd_sc_hd__and3_1
XFILLER_0_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4293__B1 _4310_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4596__B2 _4276_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5928_ _6461_/Q _5927_/X _5974_/S vssd1 vssd1 vccd1 vccd1 _5928_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_75_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5859_ _5852_/A _5785_/Y _5858_/X _5874_/S vssd1 vssd1 vccd1 vccd1 _5859_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_16_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5848__A1 _6366_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5950__A _6426_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4285__B _5767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4716__D _5369_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4505__S _4509_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5784__B1 _5977_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4339__A1 _4782_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5536__A0 _6459_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3210_ _4675_/A _5317_/A vssd1 vssd1 vccd1 vccd1 _5323_/A sky130_fd_sc_hd__nor2_1
X_4190_ _4190_/A _4190_/B vssd1 vssd1 vccd1 vccd1 _4191_/B sky130_fd_sc_hd__xnor2_1
X_3141_ _3497_/B _4358_/B vssd1 vssd1 vccd1 vccd1 _5522_/B sky130_fd_sc_hd__nor2_1
X_3072_ _5105_/S vssd1 vssd1 vccd1 vccd1 _3072_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_89_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4578__A1 _4276_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3974_ _3974_/A _3974_/B vssd1 vssd1 vccd1 vccd1 _3975_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5713_ _5713_/A _5713_/B _5713_/C vssd1 vssd1 vccd1 vccd1 _5713_/X sky130_fd_sc_hd__or3_1
XFILLER_0_45_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5790__A3 _5866_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5527__B1 _4300_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5644_ _5644_/A _5734_/S vssd1 vssd1 vccd1 vccd1 _5645_/C sky130_fd_sc_hd__and2_1
XFILLER_0_79_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold200 _4476_/X vssd1 vssd1 vccd1 vccd1 _6187_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5575_ _5562_/B _5565_/B _5562_/A vssd1 vssd1 vccd1 vccd1 _5576_/B sky130_fd_sc_hd__o21ba_1
XFILLER_0_25_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold211 _6190_/Q vssd1 vssd1 vccd1 vccd1 hold211/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold244 _6352_/Q vssd1 vssd1 vccd1 vccd1 _3088_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold222 _6223_/Q vssd1 vssd1 vccd1 vccd1 hold222/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold233 _3955_/X vssd1 vssd1 vccd1 vccd1 _6112_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4526_ _4456_/X hold228/X _4527_/S vssd1 vssd1 vccd1 vccd1 _4526_/X sky130_fd_sc_hd__mux2_1
Xhold277 _6256_/Q vssd1 vssd1 vccd1 vccd1 hold277/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold255 _6209_/Q vssd1 vssd1 vccd1 vccd1 hold255/X sky130_fd_sc_hd__dlygate4sd3_1
X_4457_ hold97/X _4456_/X _4464_/S vssd1 vssd1 vccd1 vccd1 hold98/A sky130_fd_sc_hd__mux2_1
Xhold266 _6450_/Q vssd1 vssd1 vccd1 vccd1 hold266/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3408_ _3308_/B _5522_/D _3407_/X _5309_/A _3632_/D vssd1 vssd1 vccd1 vccd1 _3408_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5770__A _6436_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold299 _6002_/X vssd1 vssd1 vccd1 vccd1 _6447_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold288 _6350_/Q vssd1 vssd1 vccd1 vccd1 _6032_/A sky130_fd_sc_hd__dlygate4sd3_1
X_4388_ hold306/X _4387_/X _5232_/S vssd1 vssd1 vccd1 vccd1 _6150_/D sky130_fd_sc_hd__mux2_1
X_6127_ _6412_/CLK _6127_/D vssd1 vssd1 vccd1 vccd1 _6127_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3339_ _3489_/B _6432_/Q _5145_/A vssd1 vssd1 vccd1 vccd1 _3673_/B sky130_fd_sc_hd__o21ai_4
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6058_ _6101_/A _6057_/X _6071_/S vssd1 vssd1 vccd1 vccd1 _6058_/X sky130_fd_sc_hd__o21a_1
X_5009_ _5109_/A1 _5006_/X _5008_/X _4924_/C vssd1 vssd1 vccd1 vccd1 _5009_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4018__A0 _6381_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4569__A1 _6334_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5766__A0 _6316_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5781__A3 _5317_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3544__A2 _3525_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5297__A2 _5299_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5049__A2 _5108_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3783__A2 _6076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3690_ _5146_/B _5405_/B _5317_/B _5777_/A vssd1 vssd1 vccd1 vccd1 _3693_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_54_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5066__S _5105_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5360_ _5360_/A _5360_/B _5360_/C vssd1 vssd1 vccd1 vccd1 _5360_/Y sky130_fd_sc_hd__nor3_1
XFILLER_0_2_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5291_ _6465_/Q _5290_/X _5291_/S vssd1 vssd1 vccd1 vccd1 _5291_/X sky130_fd_sc_hd__mux2_1
X_4311_ _4312_/B _4306_/X _4310_/X _5581_/S vssd1 vssd1 vccd1 vccd1 _4311_/X sky130_fd_sc_hd__a22o_1
X_4242_ _4276_/A _4338_/B vssd1 vssd1 vccd1 vccd1 _4261_/A sky130_fd_sc_hd__nand2_1
X_4173_ _3773_/Y _5171_/A _4170_/X _4172_/X vssd1 vssd1 vccd1 vccd1 _4173_/X sky130_fd_sc_hd__a211o_1
X_3124_ _3323_/A _3168_/B _3229_/A vssd1 vssd1 vccd1 vccd1 _4260_/B sky130_fd_sc_hd__or3_4
XFILLER_0_93_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3055_ _3168_/B vssd1 vssd1 vccd1 vccd1 _3211_/B sky130_fd_sc_hd__inv_2
XFILLER_0_77_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3957_ hold93/A _3799_/X _3801_/X hold95/A vssd1 vssd1 vccd1 vccd1 _3957_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_18_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3984__S _4716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4971__A1 _5109_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3888_ _3885_/Y _3887_/Y _3816_/B _3883_/X vssd1 vssd1 vccd1 vccd1 _4401_/B sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_5_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4971__B2 _4924_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3285__A _3352_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5627_ _5734_/S vssd1 vssd1 vccd1 vccd1 _5630_/D sky130_fd_sc_hd__inv_2
XFILLER_0_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3596__A1_N _3632_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5558_ hold556/X _5557_/X _6104_/S vssd1 vssd1 vccd1 vccd1 _5558_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4509_ _4463_/X hold284/X _4509_/S vssd1 vssd1 vccd1 vccd1 _6217_/D sky130_fd_sc_hd__mux2_1
X_5489_ hold601/X _5488_/X _5489_/S vssd1 vssd1 vccd1 vccd1 _5489_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3732__B _3885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_hold629_A _6316_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3765__A2 _6333_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3907__B _4463_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_31_wb_clk_i_A clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_7_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6470_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__3642__B _5478_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3361__C _6335_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4754__A2_N _4720_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_25 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3453__B2 _3674_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4860_ _4859_/Y hold340/X _5098_/S vssd1 vssd1 vccd1 vccd1 _4860_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_74_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3811_ _3865_/S _3811_/B vssd1 vssd1 vccd1 vccd1 _4537_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_67_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4791_ _6431_/Q _6442_/Q _6257_/Q vssd1 vssd1 vccd1 vccd1 _4791_/Y sky130_fd_sc_hd__nand3_2
XFILLER_0_55_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3742_ _6284_/Q _3744_/B vssd1 vssd1 vccd1 vccd1 _3743_/B sky130_fd_sc_hd__and2_1
XANTENNA__3756__A2 _6284_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3673_ _4344_/A _3673_/B vssd1 vssd1 vccd1 vccd1 _5603_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_70_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6461_ _6465_/CLK _6461_/D fanout181/X vssd1 vssd1 vccd1 vccd1 _6461_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_15_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3817__B _3884_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4705__A1 _4715_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5412_ _5757_/A _6475_/Q _5413_/B _5411_/Y vssd1 vssd1 vccd1 vccd1 _5432_/A sky130_fd_sc_hd__a22o_1
X_6392_ _6452_/CLK hold32/X vssd1 vssd1 vccd1 vccd1 hold31/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5343_ _5364_/A _5339_/X _5342_/X _4289_/C vssd1 vssd1 vccd1 vccd1 _5343_/X sky130_fd_sc_hd__o31a_1
XFILLER_0_2_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5274_ _6403_/Q _6402_/Q _6405_/Q _6404_/Q vssd1 vssd1 vccd1 vccd1 _5275_/D sky130_fd_sc_hd__or4_1
X_4225_ _3979_/A _5160_/B _4216_/Y _4224_/X vssd1 vssd1 vccd1 vccd1 _4225_/X sky130_fd_sc_hd__a211o_1
X_4156_ _4156_/A _4156_/B vssd1 vssd1 vccd1 vccd1 _4156_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__5681__A2 _5721_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3107_ _3168_/B _3323_/A vssd1 vssd1 vccd1 vccd1 _3547_/C sky130_fd_sc_hd__and2b_2
XANTENNA__4664__A input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4087_ _4087_/A _4087_/B vssd1 vssd1 vccd1 vccd1 _4087_/X sky130_fd_sc_hd__and2_1
XANTENNA__3995__A2 _6085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5197__A1 _6383_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5197__B2 _6378_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4989_ _5026_/C _4988_/Y _5108_/S vssd1 vssd1 vccd1 vccd1 _4989_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_73_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3743__A _4150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold579_A _6424_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5657__C1 _5731_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3181__C _3205_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3435__A1 _3632_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4513__S _4518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput15 io_in[31] vssd1 vssd1 vccd1 vccd1 _3099_/A sky130_fd_sc_hd__buf_1
XANTENNA__4699__B1 _4714_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5852__B _5867_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5896__C1 _6021_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3371__B1 _3674_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4010_ _4007_/X _4008_/Y _4009_/X vssd1 vssd1 vccd1 vccd1 _4010_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_28_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5961_ _5961_/A _5961_/B vssd1 vssd1 vccd1 vccd1 _5961_/Y sky130_fd_sc_hd__xnor2_1
X_4912_ _4911_/X _6366_/Q _5848_/S vssd1 vssd1 vccd1 vccd1 _4912_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5179__A1 _6334_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5892_ _6402_/Q _6421_/Q _5892_/S vssd1 vssd1 vccd1 vccd1 _5892_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_90_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4843_ _6204_/Q _6212_/Q _6451_/Q _6228_/Q _5404_/A0 _5078_/S1 vssd1 vssd1 vccd1
+ vccd1 _4843_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_90_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4774_ _3305_/B _3404_/B _3522_/X _3786_/Y _4773_/X vssd1 vssd1 vccd1 vccd1 _4774_/Y
+ sky130_fd_sc_hd__a221oi_4
XFILLER_0_74_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3725_ hold41/A _3701_/B _4463_/S vssd1 vssd1 vccd1 vccd1 _3725_/X sky130_fd_sc_hd__o21a_1
X_6444_ _6444_/CLK hold2/X fanout178/X vssd1 vssd1 vccd1 vccd1 _6444_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3656_ _6164_/Q _6167_/Q input1/X vssd1 vssd1 vccd1 vccd1 _3656_/X sky130_fd_sc_hd__mux2_4
XANTENNA_fanout115_A _5489_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5254__S _5489_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3587_ _5605_/A _3587_/B vssd1 vssd1 vccd1 vccd1 _4676_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_61_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6375_ _6376_/CLK _6375_/D fanout172/X vssd1 vssd1 vccd1 vccd1 _6375_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_0_2_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5326_ _3240_/B _3228_/C _3204_/X _3219_/Y vssd1 vssd1 vccd1 vccd1 _5327_/D sky130_fd_sc_hd__a31o_1
X_5257_ _5257_/A _5257_/B _5257_/C vssd1 vssd1 vccd1 vccd1 _5257_/X sky130_fd_sc_hd__or3_1
XANTENNA__5103__A1 _6316_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4208_ _6290_/Q _4207_/C _6291_/Q vssd1 vssd1 vccd1 vccd1 _4209_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_48_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5188_ _5187_/A _5187_/B _5600_/A vssd1 vssd1 vccd1 vccd1 _5188_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_97_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4139_ _4138_/X hold223/X _4241_/S vssd1 vssd1 vccd1 vccd1 _6116_/D sky130_fd_sc_hd__mux2_1
XANTENNA__5002__B _5002_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5342__A1 _5605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout181 fanout185/X vssd1 vssd1 vccd1 vccd1 fanout181/X sky130_fd_sc_hd__clkbuf_8
Xfanout170 fanout171/X vssd1 vssd1 vccd1 vccd1 fanout170/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__4508__S _4509_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3959__A2 _3804_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4908__A1 _6463_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4908__B2 _5109_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3510_ _3699_/A _3503_/Y _3638_/B hold575/X _3509_/X vssd1 vssd1 vccd1 vccd1 _3510_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold618 _6459_/Q vssd1 vssd1 vccd1 vccd1 hold618/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold607 _6364_/Q vssd1 vssd1 vccd1 vccd1 hold607/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4490_ _4182_/X hold138/X _4491_/S vssd1 vssd1 vccd1 vccd1 _6200_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_100_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3441_ _3432_/X _3440_/X _5522_/A vssd1 vssd1 vccd1 vccd1 _3441_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__5333__A1 _5757_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold629 _6316_/Q vssd1 vssd1 vccd1 vccd1 hold629/X sky130_fd_sc_hd__buf_1
XANTENNA__4136__A2 _4462_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3372_ _3372_/A vssd1 vssd1 vccd1 vccd1 _3372_/Y sky130_fd_sc_hd__inv_2
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6160_ _6474_/CLK _6160_/D fanout179/X vssd1 vssd1 vccd1 vccd1 _6160_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__4198__B _6385_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5111_ _6409_/Q _5110_/X _5971_/S vssd1 vssd1 vccd1 vccd1 _5111_/X sky130_fd_sc_hd__mux2_1
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5097__A0 _6408_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6091_ _5565_/Y _6037_/B _6101_/B _5041_/B vssd1 vssd1 vccd1 vccd1 _6091_/X sky130_fd_sc_hd__o2bb2a_1
XANTENNA__5636__A2 _5721_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5042_ _6313_/Q _4963_/B _5041_/B _4796_/Y vssd1 vssd1 vccd1 vccd1 _5042_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_79_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6061__A2 _4901_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5944_ _5933_/A _5943_/X _5977_/S vssd1 vssd1 vccd1 vccd1 _5944_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4942__A _5102_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5757__B _5757_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5875_ _6368_/Q _6420_/Q _5892_/S vssd1 vssd1 vccd1 vccd1 _5875_/X sky130_fd_sc_hd__mux2_1
X_4826_ _6414_/Q _6362_/Q _5105_/S vssd1 vssd1 vccd1 vccd1 _4826_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_35_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3277__B _4324_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4757_ _4755_/X _4756_/X _5289_/S vssd1 vssd1 vccd1 vccd1 _4757_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_31_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4688_ _6085_/A _4714_/S vssd1 vssd1 vccd1 vccd1 _4688_/Y sky130_fd_sc_hd__nor2_1
X_3708_ _6352_/Q _6033_/B _4670_/D vssd1 vssd1 vccd1 vccd1 _4398_/B sky130_fd_sc_hd__or3_1
XFILLER_0_31_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3639_ _5605_/A _5322_/A _3639_/C _3639_/D vssd1 vssd1 vccd1 vccd1 _3640_/C sky130_fd_sc_hd__or4_2
XANTENNA__5324__A1 _4675_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4127__A2 _3731_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6427_ _6428_/CLK _6427_/D fanout172/X vssd1 vssd1 vccd1 vccd1 _6427_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_31_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6276__SET_B fanout183/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6358_ _6470_/CLK _6358_/D fanout179/X vssd1 vssd1 vccd1 vccd1 _6358_/Q sky130_fd_sc_hd__dfrtp_1
X_5309_ _5309_/A _5345_/A _5345_/B _5309_/D vssd1 vssd1 vccd1 vccd1 _5311_/C sky130_fd_sc_hd__or4_1
X_6289_ _6465_/CLK _6289_/D vssd1 vssd1 vccd1 vccd1 _6289_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__5088__B1 _5108_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_21_wb_clk_i _6448_/CLK vssd1 vssd1 vccd1 vccd1 _6312_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_93_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3468__A _6021_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4290__C _4768_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5618__A2 _4332_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4 hold4/A vssd1 vssd1 vccd1 vccd1 hold4/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3990_ _3759_/Y _3987_/B _3989_/X _3985_/X vssd1 vssd1 vccd1 vccd1 _3991_/C sky130_fd_sc_hd__a211o_1
XFILLER_0_69_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5069__S _5108_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5660_ _6334_/Q _5628_/X _5653_/X _6484_/Q _5654_/X vssd1 vssd1 vccd1 vccd1 _5663_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_72_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4611_ _4611_/A _4611_/B vssd1 vssd1 vccd1 vccd1 _4611_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__5003__B1 _5002_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5591_ hold531/X _5590_/X _6104_/S vssd1 vssd1 vccd1 vccd1 _5591_/X sky130_fd_sc_hd__mux2_1
X_4542_ hold286/X _4441_/X _4545_/S vssd1 vssd1 vccd1 vccd1 _6253_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_25_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5306__A1 _3205_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold426 _5664_/X vssd1 vssd1 vccd1 vccd1 _6379_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold404 _5760_/X vssd1 vssd1 vccd1 vccd1 _6404_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold415 _6325_/Q vssd1 vssd1 vccd1 vccd1 hold415/X sky130_fd_sc_hd__dlygate4sd3_1
X_4473_ hold145/X _4240_/X _4473_/S vssd1 vssd1 vccd1 vccd1 _4473_/X sky130_fd_sc_hd__mux2_1
X_3424_ _4289_/B _3424_/B _3424_/C _3423_/X vssd1 vssd1 vccd1 vccd1 _3424_/X sky130_fd_sc_hd__or4b_1
Xhold448 _6277_/Q vssd1 vssd1 vccd1 vccd1 hold448/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold437 _4561_/X vssd1 vssd1 vccd1 vccd1 _6268_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold459 _4564_/X vssd1 vssd1 vccd1 vccd1 _6271_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6212_ _6456_/CLK _6212_/D vssd1 vssd1 vccd1 vccd1 _6212_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3355_ _5600_/A _5323_/C _3355_/C _3355_/D vssd1 vssd1 vccd1 vccd1 _3355_/X sky130_fd_sc_hd__and4bb_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6143_ _6490_/CLK hold92/X vssd1 vssd1 vccd1 vccd1 hold91/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__4656__B _4668_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3286_ _4335_/B _3489_/B vssd1 vssd1 vccd1 vccd1 _5387_/C sky130_fd_sc_hd__nor2_4
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6074_ _5519_/Y _6037_/B _6101_/B _4962_/B vssd1 vssd1 vccd1 vccd1 _6074_/X sky130_fd_sc_hd__o2bb2a_1
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5025_ _5021_/B _5024_/X _5106_/S vssd1 vssd1 vccd1 vccd1 _5025_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout182_A fanout183/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5927_ _5964_/A _5926_/X _5021_/Y vssd1 vssd1 vccd1 vccd1 _5927_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_75_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5858_ _5786_/Y _5850_/X _5857_/Y _5887_/S vssd1 vssd1 vccd1 vccd1 _5858_/X sky130_fd_sc_hd__a22o_1
X_4809_ _6361_/Q _5108_/S vssd1 vssd1 vccd1 vccd1 _4809_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__4979__S0 _5100_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5789_ _6361_/Q _5771_/A _4780_/X _5788_/X vssd1 vssd1 vccd1 vccd1 _5789_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_0_90_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5950__B _5970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4058__S _4716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4582__A _5757_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6367__RESET_B fanout175/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5784__A1 _6023_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4339__A2 _5314_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4521__S _4527_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3140_ _3414_/B _3639_/D vssd1 vssd1 vccd1 vccd1 _4358_/B sky130_fd_sc_hd__nor2_2
XANTENNA__4275__A1 _5398_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3071_ hold1/X vssd1 vssd1 vccd1 vccd1 _3469_/A sky130_fd_sc_hd__inv_2
XFILLER_0_15_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5775__A1 _6430_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4578__A2 _4595_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3973_ _3973_/A _3973_/B vssd1 vssd1 vccd1 vccd1 _3975_/A sky130_fd_sc_hd__and2_1
XFILLER_0_85_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5712_ _6314_/Q _5630_/X _5653_/X _6488_/Q _5711_/X vssd1 vssd1 vccd1 vccd1 _5713_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_85_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5643_ _5646_/B _5653_/B vssd1 vssd1 vccd1 vccd1 _5643_/X sky130_fd_sc_hd__and2_2
XANTENNA__5527__A1 _5593_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5574_ _5574_/A _5574_/B vssd1 vssd1 vccd1 vccd1 _5576_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_5_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold201 _6229_/Q vssd1 vssd1 vccd1 vccd1 hold201/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4525_ _4448_/X hold270/X _4527_/S vssd1 vssd1 vccd1 vccd1 _6231_/D sky130_fd_sc_hd__mux2_1
Xhold223 _6116_/Q vssd1 vssd1 vccd1 vccd1 hold223/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold212 _4479_/X vssd1 vssd1 vccd1 vccd1 _6190_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold234 _6118_/Q vssd1 vssd1 vccd1 vccd1 hold234/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold245 _5385_/X vssd1 vssd1 vccd1 vccd1 _6352_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold278 _4545_/X vssd1 vssd1 vccd1 vccd1 _6256_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4456_ _4453_/X _4454_/X _4455_/X _4441_/S vssd1 vssd1 vccd1 vccd1 _4456_/X sky130_fd_sc_hd__a22o_2
Xhold256 _4500_/X vssd1 vssd1 vccd1 vccd1 _6209_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold267 _6005_/X vssd1 vssd1 vccd1 vccd1 _6450_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3407_ _5777_/A _5770_/B _3406_/Y vssd1 vssd1 vccd1 vccd1 _3407_/X sky130_fd_sc_hd__a21o_1
X_4387_ _5600_/A _4253_/Y _5364_/B _4289_/C vssd1 vssd1 vccd1 vccd1 _4387_/X sky130_fd_sc_hd__a22o_1
Xhold289 _5381_/X vssd1 vssd1 vccd1 vccd1 _6350_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3338_ _3489_/B _6432_/Q _5145_/A vssd1 vssd1 vccd1 vccd1 _3338_/X sky130_fd_sc_hd__o21a_1
XANTENNA__3710__B1 _5384_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6126_ _6419_/CLK _6126_/D fanout173/X vssd1 vssd1 vccd1 vccd1 _6126_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3269_ _3278_/B _5323_/B vssd1 vssd1 vccd1 vccd1 _3685_/A sky130_fd_sc_hd__nor2_2
X_6057_ _6101_/B _4881_/X _5470_/X _6036_/X vssd1 vssd1 vccd1 vccd1 _6057_/X sky130_fd_sc_hd__o22a_1
X_5008_ _6460_/Q _5007_/X _5108_/S vssd1 vssd1 vccd1 vccd1 _5008_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4018__A1 _6385_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6460__RESET_B fanout181/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_21_wb_clk_i_A _6448_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3481__A _3489_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5900__S _5977_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4516__S _4518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6130__RESET_B fanout180/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5509__B2 _5485_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5290_ _5287_/X _5289_/X _5290_/S vssd1 vssd1 vccd1 vccd1 _5290_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_2_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4310_ _6313_/Q _4309_/Y _4310_/S vssd1 vssd1 vccd1 vccd1 _4310_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_77_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4241_ _4240_/X hold234/X _4241_/S vssd1 vssd1 vccd1 vccd1 _4241_/X sky130_fd_sc_hd__mux2_1
X_4172_ _4332_/B _3759_/Y _4171_/X _6384_/Q vssd1 vssd1 vccd1 vccd1 _4172_/X sky130_fd_sc_hd__a22o_1
X_3123_ _3323_/A _3168_/B vssd1 vssd1 vccd1 vccd1 _3216_/B sky130_fd_sc_hd__nor2_1
X_3054_ _5995_/C vssd1 vssd1 vccd1 vccd1 _5980_/A sky130_fd_sc_hd__inv_2
XANTENNA_fanout145_A _5605_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3956_ hold141/X hold95/X hold207/X hold93/X _5721_/C1 _4235_/S vssd1 vssd1 vccd1
+ vccd1 _3956_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_18_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5626_ _3172_/A _5613_/X _5625_/X _6435_/Q vssd1 vssd1 vccd1 vccd1 _5734_/S sky130_fd_sc_hd__o2bb2a_4
X_3887_ _3883_/S _3886_/X _3852_/A vssd1 vssd1 vccd1 vccd1 _3887_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_33_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5557_ _6461_/Q _5556_/X _5598_/S vssd1 vssd1 vccd1 vccd1 _5557_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5920__B2 _5976_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5488_ _6463_/Q _5487_/X _5512_/S vssd1 vssd1 vccd1 vccd1 _5488_/X sky130_fd_sc_hd__mux2_1
X_4508_ _4456_/X hold89/X _4509_/S vssd1 vssd1 vccd1 vccd1 hold90/A sky130_fd_sc_hd__mux2_1
X_4439_ _4081_/X _4438_/Y hold3/X _4462_/A2 vssd1 vssd1 vccd1 vccd1 _4439_/X sky130_fd_sc_hd__o2bb2a_1
XANTENNA__4828__C _5108_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3732__C _3884_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4239__A1 _5732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5021__A _5102_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4411__A1 _5730_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5911__A1 _6421_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output39_A _6331_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4790_ _6431_/Q _6442_/Q _6257_/Q vssd1 vssd1 vccd1 vccd1 _4790_/X sky130_fd_sc_hd__and3_2
X_3810_ _3852_/A _3883_/S _3865_/S vssd1 vssd1 vccd1 vccd1 _3810_/X sky130_fd_sc_hd__and3_4
XFILLER_0_27_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5866__A _5866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3741_ _4150_/A _6378_/Q vssd1 vssd1 vccd1 vccd1 _3744_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_55_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3756__A3 _6378_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3672_ _3674_/A _3411_/A _5617_/A _3671_/B vssd1 vssd1 vccd1 vccd1 _3672_/X sky130_fd_sc_hd__o22a_1
X_6460_ _6465_/CLK _6460_/D fanout181/X vssd1 vssd1 vccd1 vccd1 _6460_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3817__C _3818_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5411_ _5757_/A _5411_/B vssd1 vssd1 vccd1 vccd1 _5411_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__5902__A1 _6421_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6391_ _6399_/CLK hold28/X vssd1 vssd1 vccd1 vccd1 hold27/A sky130_fd_sc_hd__dfxtp_1
X_5342_ _5605_/A _4328_/A _5341_/X _3278_/A _5340_/X vssd1 vssd1 vccd1 vccd1 _5342_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_2_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5273_ _6339_/Q _5288_/S _5272_/X vssd1 vssd1 vccd1 vccd1 _5273_/Y sky130_fd_sc_hd__o21ai_1
X_4224_ _4115_/A _5263_/B _4221_/X _4223_/X vssd1 vssd1 vccd1 vccd1 _4224_/X sky130_fd_sc_hd__a211o_1
X_4155_ _4155_/A _4155_/B vssd1 vssd1 vccd1 vccd1 _4156_/B sky130_fd_sc_hd__xnor2_1
X_3106_ _3106_/A vssd1 vssd1 vccd1 vccd1 _3110_/A sky130_fd_sc_hd__inv_2
XANTENNA__5540__S _5593_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4664__B _4668_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4086_ _4085_/X hold252/X _4241_/S vssd1 vssd1 vccd1 vccd1 _6115_/D sky130_fd_sc_hd__mux2_1
XANTENNA__6091__B1 _6101_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4988_ _6370_/Q _4988_/B vssd1 vssd1 vccd1 vccd1 _4988_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__3296__A _5314_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3939_ _5427_/B _3938_/Y _6347_/Q vssd1 vssd1 vccd1 vccd1 _3939_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_46_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5609_ _5610_/B vssd1 vssd1 vccd1 vccd1 _5645_/B sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_46_wb_clk_i clkbuf_leaf_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6399_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_14_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3683__A2 _5146_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5450__S _5489_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold641_A _6129_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5424__A3 _5520_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4632__A1 _6463_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4632__B2 _6314_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput16 io_in[35] vssd1 vssd1 vccd1 vccd1 _3100_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3934__A _6337_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4699__A1 _4713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3371__A1 _5777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4871__A1 _6461_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5299__C _5299_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5960_ _5950_/Y _5954_/B _5952_/A vssd1 vssd1 vccd1 vccd1 _5961_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_87_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_2_0__f_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5891_ _5890_/A _5890_/B _5889_/Y vssd1 vssd1 vccd1 vccd1 _5912_/A sky130_fd_sc_hd__o21ba_1
X_4911_ _5971_/S _4909_/X _4910_/X _4902_/X vssd1 vssd1 vccd1 vccd1 _4911_/X sky130_fd_sc_hd__a31o_1
XANTENNA__5820__B1 _5784_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4842_ hold69/A _6188_/Q _6172_/Q _6251_/Q _5404_/A0 _5078_/S1 vssd1 vssd1 vccd1
+ vccd1 _4842_/X sky130_fd_sc_hd__mux4_1
X_4773_ _3489_/B _3305_/A _5346_/B _3561_/Y vssd1 vssd1 vccd1 vccd1 _4773_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_62_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3724_ _3712_/Y _3715_/Y _3721_/X _3722_/X vssd1 vssd1 vccd1 vccd1 _3883_/S sky130_fd_sc_hd__o31a_4
XFILLER_0_7_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3655_ _6023_/A _3655_/B vssd1 vssd1 vccd1 vccd1 _6440_/D sky130_fd_sc_hd__nor2_1
X_6443_ _6470_/CLK _6443_/D fanout177/X vssd1 vssd1 vccd1 vccd1 _6443_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3586_ _5367_/B _3586_/B vssd1 vssd1 vccd1 vccd1 _6441_/D sky130_fd_sc_hd__nor2_1
X_6374_ _6376_/CLK _6374_/D fanout172/X vssd1 vssd1 vccd1 vccd1 _6374_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3362__B2 _6335_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5325_ _4675_/A _3590_/A _4676_/A _5324_/X vssd1 vssd1 vccd1 vccd1 _5325_/X sky130_fd_sc_hd__a211o_1
X_5256_ _5256_/A _5256_/B _5163_/A vssd1 vssd1 vccd1 vccd1 _5257_/C sky130_fd_sc_hd__or3b_1
XFILLER_0_54_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5103__A2 _4963_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4207_ _5268_/A _6290_/Q _4207_/C vssd1 vssd1 vccd1 vccd1 _4209_/A sky130_fd_sc_hd__or3_1
XANTENNA__4675__A _4675_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5187_ _5187_/A _5187_/B vssd1 vssd1 vccd1 vccd1 _5187_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_97_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4138_ _4135_/X _4136_/X _4137_/X _4441_/S vssd1 vssd1 vccd1 vccd1 _4138_/X sky130_fd_sc_hd__a22o_2
XFILLER_0_97_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4069_ _3753_/X _4064_/X _4068_/Y _5136_/B _4067_/X vssd1 vssd1 vccd1 vccd1 _4070_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_64_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5878__A0 _6368_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3473__B _4363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout160 _3172_/A vssd1 vssd1 vccd1 vccd1 _3168_/B sky130_fd_sc_hd__buf_4
Xfanout182 fanout183/X vssd1 vssd1 vccd1 vccd1 fanout182/X sky130_fd_sc_hd__clkbuf_8
Xfanout171 fanout172/X vssd1 vssd1 vccd1 vccd1 fanout171/X sky130_fd_sc_hd__buf_4
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4081__A2 _6093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4524__S _4527_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5030__A1 _5109_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4908__A2 _4963_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5030__B2 _4924_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3592__A1 _5777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold608 _5463_/X vssd1 vssd1 vccd1 vccd1 _6364_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold619 _6343_/Q vssd1 vssd1 vccd1 vccd1 hold619/X sky130_fd_sc_hd__dlygate4sd3_1
X_3440_ _3440_/A _3440_/B _3440_/C _3437_/Y vssd1 vssd1 vccd1 vccd1 _3440_/X sky130_fd_sc_hd__or4b_1
XFILLER_0_69_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3371_ _5777_/A _4784_/B _5617_/B _3674_/A vssd1 vssd1 vccd1 vccd1 _3372_/A sky130_fd_sc_hd__a31o_1
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5110_ _6428_/Q _4793_/Y _5104_/X _5109_/X vssd1 vssd1 vccd1 vccd1 _5110_/X sky130_fd_sc_hd__a211o_1
X_6090_ _4366_/A _6088_/X _6089_/Y hold522/X _6077_/Y vssd1 vssd1 vccd1 vccd1 _6090_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_0_85_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5041_ _5102_/A _5041_/B vssd1 vssd1 vccd1 vccd1 _5041_/Y sky130_fd_sc_hd__nand2_1
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
X_5943_ _5942_/X _5937_/X _5976_/S vssd1 vssd1 vccd1 vccd1 _5943_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5757__C _5757_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5874_ hold524/X _5873_/X _5874_/S vssd1 vssd1 vccd1 vccd1 _5874_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_34_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4825_ _6476_/Q _4794_/Y _4963_/B _6459_/Q _4824_/Y vssd1 vssd1 vccd1 vccd1 _4825_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_28_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4455__S0 _5731_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3583__A1 _4313_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4756_ hold502/X _4319_/B _4768_/S vssd1 vssd1 vccd1 vccd1 _4756_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_7_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4687_ _6384_/Q _4686_/X _4712_/S vssd1 vssd1 vccd1 vccd1 _4687_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3574__A _6435_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3707_ _6350_/Q _6351_/Q vssd1 vssd1 vccd1 vccd1 _4670_/D sky130_fd_sc_hd__and2_1
XANTENNA__4780__B1 _5974_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3638_ _5400_/A _3638_/B _3638_/C vssd1 vssd1 vccd1 vccd1 _3648_/B sky130_fd_sc_hd__nor3_1
X_6426_ _6426_/CLK _6426_/D fanout171/X vssd1 vssd1 vccd1 vccd1 _6426_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_31_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3569_ _5317_/B _3569_/B vssd1 vssd1 vccd1 vccd1 _3569_/X sky130_fd_sc_hd__or2_1
X_6357_ _6377_/CLK _6357_/D fanout179/X vssd1 vssd1 vccd1 vccd1 _6357_/Q sky130_fd_sc_hd__dfrtp_1
X_5308_ _5369_/B _5757_/C _3305_/B _3570_/B vssd1 vssd1 vccd1 vccd1 _5309_/D sky130_fd_sc_hd__a211o_1
XFILLER_0_11_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6288_ _6441_/CLK _6288_/D vssd1 vssd1 vccd1 vccd1 _6288_/Q sky130_fd_sc_hd__dfxtp_4
X_5239_ _5783_/A _5239_/B vssd1 vssd1 vccd1 vccd1 _5239_/X sky130_fd_sc_hd__or2_1
XFILLER_0_98_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4771__A0 hold629/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5720__C1 _5730_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5 hold5/A vssd1 vssd1 vccd1 vccd1 hold5/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_71_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4610_ _5757_/B hold452/X _4582_/Y _4609_/X vssd1 vssd1 vccd1 vccd1 _4610_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_44_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5003__A1 _6311_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3565__A1 _4557_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5590_ _6464_/Q _5589_/X _5598_/S vssd1 vssd1 vccd1 vccd1 _5590_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_37_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4541_ hold206/X _4435_/X _4545_/S vssd1 vssd1 vccd1 vccd1 _6252_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_4_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold405 _6354_/Q vssd1 vssd1 vccd1 vccd1 hold405/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold427 _6330_/Q vssd1 vssd1 vccd1 vccd1 hold427/X sky130_fd_sc_hd__dlygate4sd3_1
X_4472_ hold107/X _4182_/X _4473_/S vssd1 vssd1 vccd1 vccd1 _4472_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_13_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold416 _4978_/X vssd1 vssd1 vccd1 vccd1 _6325_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3423_ _3786_/A _3258_/B _5522_/D _3691_/B vssd1 vssd1 vccd1 vccd1 _3423_/X sky130_fd_sc_hd__o31a_1
Xhold449 _4570_/X vssd1 vssd1 vccd1 vccd1 _6277_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold438 _6273_/Q vssd1 vssd1 vccd1 vccd1 hold438/X sky130_fd_sc_hd__dlygate4sd3_1
X_6211_ _6452_/CLK _6211_/D vssd1 vssd1 vccd1 vccd1 _6211_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6142_ _6399_/CLK _6142_/D vssd1 vssd1 vccd1 vccd1 _6142_/Q sky130_fd_sc_hd__dfxtp_1
X_3354_ _5146_/B _4251_/B vssd1 vssd1 vccd1 vccd1 _5323_/C sky130_fd_sc_hd__nor2_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4278__C1 _5600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3285_ _3352_/B _3285_/B _3355_/C _3285_/D vssd1 vssd1 vccd1 vccd1 _3285_/Y sky130_fd_sc_hd__nand4_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6073_ _6073_/A _6073_/B vssd1 vssd1 vccd1 vccd1 _6107_/S sky130_fd_sc_hd__or2_4
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4429__S _4464_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6019__A0 _4668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5024_ _6424_/Q _6372_/Q _5105_/S vssd1 vssd1 vccd1 vccd1 _5024_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4293__A2 _3506_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout175_A fanout176/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3569__A _5317_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5926_ _6372_/Q _5848_/S _5972_/B1 _5925_/X vssd1 vssd1 vccd1 vccd1 _5926_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_8_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5857_ _5857_/A _5872_/B vssd1 vssd1 vccd1 vccd1 _5857_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_35_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_11_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_5788_ _6361_/Q _5861_/S _5842_/B1 _5787_/X _5102_/A vssd1 vssd1 vccd1 vccd1 _5788_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_8_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4979__S1 _5100_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4808_ _5108_/S vssd1 vssd1 vccd1 vccd1 _4808_/Y sky130_fd_sc_hd__inv_2
X_4739_ _4737_/X _4738_/X _5289_/S vssd1 vssd1 vccd1 vccd1 _4739_/X sky130_fd_sc_hd__mux2_1
X_6409_ _6409_/CLK _6409_/D fanout170/X vssd1 vssd1 vccd1 vccd1 _6409_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_31_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout88_A _4360_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold387_A _6327_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold554_A _6380_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_50_wb_clk_i_A clkbuf_leaf_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_94_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5784__A2 _5976_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4103__A _6333_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3070_ _4366_/A vssd1 vssd1 vccd1 vccd1 _6108_/S sky130_fd_sc_hd__inv_2
XFILLER_0_89_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3972_ _6286_/Q _3972_/B _3972_/C vssd1 vssd1 vccd1 vccd1 _3973_/B sky130_fd_sc_hd__or3_1
XFILLER_0_45_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5711_ _6463_/Q _5645_/X _5710_/X _5632_/Y vssd1 vssd1 vccd1 vccd1 _5711_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4983__B1 _4982_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4712__S _4712_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5642_ _5644_/A _5734_/S vssd1 vssd1 vccd1 vccd1 _5653_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_72_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5573_ _5594_/A _5573_/B vssd1 vssd1 vccd1 vccd1 _5574_/B sky130_fd_sc_hd__or2_1
XFILLER_0_5_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold202 _4523_/X vssd1 vssd1 vccd1 vccd1 _6229_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4524_ _4441_/X hold262/X _4527_/S vssd1 vssd1 vccd1 vccd1 _6230_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_40_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold213 _6198_/Q vssd1 vssd1 vccd1 vccd1 hold213/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold235 _4241_/X vssd1 vssd1 vccd1 vccd1 _6118_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold224 _6212_/Q vssd1 vssd1 vccd1 vccd1 hold224/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3852__A _3852_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold257 _6136_/Q vssd1 vssd1 vccd1 vccd1 hold257/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold268 _6178_/Q vssd1 vssd1 vccd1 vccd1 hold268/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold246 _6454_/Q vssd1 vssd1 vccd1 vccd1 hold246/X sky130_fd_sc_hd__dlygate4sd3_1
X_4455_ hold89/X hold53/X hold113/X hold51/X _5731_/C1 _4420_/S vssd1 vssd1 vccd1
+ vccd1 _4455_/X sky130_fd_sc_hd__mux4_1
X_3406_ _5317_/B _5770_/B _3786_/A vssd1 vssd1 vccd1 vccd1 _3406_/Y sky130_fd_sc_hd__a21oi_2
Xhold279 _6244_/Q vssd1 vssd1 vccd1 vccd1 _3493_/A sky130_fd_sc_hd__dlygate4sd3_1
X_4386_ _4386_/A _4386_/B vssd1 vssd1 vccd1 vccd1 _5364_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_0_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3337_ _3786_/A _3685_/A vssd1 vssd1 vccd1 vccd1 _3424_/B sky130_fd_sc_hd__nor2_1
X_6125_ _6316_/CLK _6125_/D fanout174/X vssd1 vssd1 vccd1 vccd1 _6125_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3268_ _5387_/B _3268_/B vssd1 vssd1 vccd1 vccd1 _4386_/A sky130_fd_sc_hd__or2_2
XANTENNA__3998__S _4463_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6056_ _4366_/A _6054_/X _6055_/Y hold483/X _6040_/Y vssd1 vssd1 vccd1 vccd1 _6056_/X
+ sky130_fd_sc_hd__o32a_1
X_3199_ _3326_/A _3229_/C vssd1 vssd1 vccd1 vccd1 _4248_/C sky130_fd_sc_hd__nor2_2
X_5007_ _6371_/Q _5026_/C vssd1 vssd1 vccd1 vccd1 _5007_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_68_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3777__A1 _6378_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4423__C1 _5655_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5909_ _5901_/A _5785_/Y _5908_/X _5977_/S vssd1 vssd1 vccd1 vccd1 _5909_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_36_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3529__A1 _4332_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4821__S0 _5078_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4577__B _4595_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5454__A1 _5492_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4965__A0 _6421_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4532__S _4536_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5390__B1 _5607_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4240_ _4229_/X _4230_/X _4239_/X _4441_/S vssd1 vssd1 vccd1 vccd1 _4240_/X sky130_fd_sc_hd__a22o_2
X_4171_ _4332_/B _4223_/A _4168_/Y _3759_/Y vssd1 vssd1 vccd1 vccd1 _4171_/X sky130_fd_sc_hd__a211o_1
X_3122_ _3530_/A _3497_/B _6434_/Q vssd1 vssd1 vccd1 vccd1 _3122_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_93_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4707__S _4711_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4879__S0 _5100_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6258__RESET_B fanout181/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3955_ _3954_/X hold232/X _4241_/S vssd1 vssd1 vccd1 vccd1 _3955_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4956__A0 _6368_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4442__S _4464_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4708__A0 _6286_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5625_ _3699_/A _5624_/X _5146_/C _5616_/X vssd1 vssd1 vccd1 vccd1 _5625_/X sky130_fd_sc_hd__o2bb2a_1
X_3886_ _6226_/Q _6449_/Q _3886_/S vssd1 vssd1 vccd1 vccd1 _3886_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout138_A _5404_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5556_ hold556/X _5555_/X _6070_/A vssd1 vssd1 vccd1 vccd1 _5556_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_5_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5920__A2 _5786_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5487_ _5485_/X _5486_/X _5567_/B vssd1 vssd1 vccd1 vccd1 _5487_/X sky130_fd_sc_hd__mux2_1
X_4507_ _4448_/X hold67/X _4509_/S vssd1 vssd1 vccd1 vccd1 hold68/A sky130_fd_sc_hd__mux2_1
X_4438_ _4438_/A _5301_/A vssd1 vssd1 vccd1 vccd1 _4438_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_1_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4369_ hold283/X _3911_/X _4376_/S vssd1 vssd1 vccd1 vccd1 _6134_/D sky130_fd_sc_hd__mux2_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6108_ hold594/X _6107_/X _6108_/S vssd1 vssd1 vccd1 vccd1 _6490_/D sky130_fd_sc_hd__mux2_1
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6039_ _6039_/A vssd1 vssd1 vccd1 vccd1 _6039_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_68_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5021__B _5021_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5448__S _5499_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5911__A2 _6422_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5675__A1 _5757_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4527__S _4527_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5212__A _6461_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3989__B2 _6380_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5866__B _6464_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3740_ _6345_/Q _3740_/B vssd1 vssd1 vccd1 vccd1 _5136_/B sky130_fd_sc_hd__and2_4
XANTENNA__6043__A _6076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4402__A2 _4462_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5038__S0 _5404_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3671_ _5617_/A _3671_/B vssd1 vssd1 vccd1 vccd1 _5603_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_42_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5410_ _5410_/A _5410_/B vssd1 vssd1 vccd1 vccd1 _5512_/S sky130_fd_sc_hd__nand2_4
XANTENNA__5902__A2 _5970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6390_ _6393_/CLK hold4/X vssd1 vssd1 vccd1 vccd1 hold3/A sky130_fd_sc_hd__dfxtp_1
X_5341_ _5605_/B _6429_/Q vssd1 vssd1 vccd1 vccd1 _5341_/X sky130_fd_sc_hd__or2_1
XFILLER_0_2_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5115__A0 _6409_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5272_ _6281_/Q _5783_/A _4555_/Y _4723_/X vssd1 vssd1 vccd1 vccd1 _5272_/X sky130_fd_sc_hd__o31a_1
XANTENNA__5666__B2 _6423_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5666__A1 _6335_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4223_ _4223_/A _5199_/A vssd1 vssd1 vccd1 vccd1 _4223_/X sky130_fd_sc_hd__and2_1
X_4154_ _4095_/A _4095_/B _4096_/B vssd1 vssd1 vccd1 vccd1 _4155_/B sky130_fd_sc_hd__a21o_1
X_3105_ _5124_/A _3247_/A vssd1 vssd1 vccd1 vccd1 _3106_/A sky130_fd_sc_hd__or2_2
X_4085_ _4082_/Y _4083_/X _4084_/X _4441_/S vssd1 vssd1 vccd1 vccd1 _4085_/X sky130_fd_sc_hd__a22o_2
XANTENNA__5122__A _6021_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6091__B2 _5041_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4987_ _6370_/Q _4988_/B vssd1 vssd1 vccd1 vccd1 _5026_/C sky130_fd_sc_hd__and2_1
X_3938_ _3938_/A _3938_/B vssd1 vssd1 vccd1 vccd1 _3938_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_46_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3869_ hold159/X hold171/X _3884_/S vssd1 vssd1 vccd1 vccd1 _3869_/X sky130_fd_sc_hd__mux2_1
X_5608_ _5980_/A _5608_/B vssd1 vssd1 vccd1 vccd1 _5610_/B sky130_fd_sc_hd__and2_2
XANTENNA__4900__S _5101_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5539_ _5519_/A _5519_/B _5532_/A _5532_/B _5538_/Y vssd1 vssd1 vccd1 vccd1 _5545_/A
+ sky130_fd_sc_hd__o41a_1
XFILLER_0_41_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_15_wb_clk_i _6448_/CLK vssd1 vssd1 vccd1 vccd1 _6441_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__5409__A1 _6430_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5409__B2 _5600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6082__A1 _4366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold634_A _6339_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3840__B1 _3795_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput17 io_in[4] vssd1 vssd1 vccd1 vccd1 _3501_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__5896__A1 _6458_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5207__A _6463_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5648__A1 _6333_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5648__B2 _6309_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output51_A _3662_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4871__A2 _4963_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5890_ _5890_/A _5890_/B _5889_/Y vssd1 vssd1 vccd1 vccd1 _5898_/B sky130_fd_sc_hd__or3b_1
X_4910_ _6418_/Q _4930_/B vssd1 vssd1 vccd1 vccd1 _4910_/X sky130_fd_sc_hd__or2_1
XFILLER_0_87_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4841_ _6363_/Q _4790_/X _4789_/B vssd1 vssd1 vccd1 vccd1 _4841_/X sky130_fd_sc_hd__a21o_1
XANTENNA__4387__A1 _5600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4772_ _6023_/A _5499_/S _3503_/B vssd1 vssd1 vccd1 vccd1 _5116_/S sky130_fd_sc_hd__o21ai_2
XFILLER_0_7_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3723_ _3712_/Y _3715_/Y _3721_/X _3722_/X vssd1 vssd1 vccd1 vccd1 _3723_/Y sky130_fd_sc_hd__o31ai_2
X_3654_ _4325_/A _3374_/Y _3620_/X hold185/X vssd1 vssd1 vccd1 vccd1 _3654_/X sky130_fd_sc_hd__o22a_1
X_6442_ _6474_/CLK _6442_/D fanout181/X vssd1 vssd1 vccd1 vccd1 _6442_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_3_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5816__S _5816_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3585_ hold636/X _5218_/S _3584_/X _3368_/S _5605_/B vssd1 vssd1 vccd1 vccd1 _3586_/B
+ sky130_fd_sc_hd__o221a_1
X_6373_ _6428_/CLK _6373_/D fanout172/X vssd1 vssd1 vccd1 vccd1 _6373_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_11_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5324_ _4675_/A _4281_/A _5364_/B _5316_/Y _5323_/X vssd1 vssd1 vccd1 vccd1 _5324_/X
+ sky130_fd_sc_hd__o32a_1
X_5255_ _3368_/S _6342_/Q _5162_/A _5162_/B vssd1 vssd1 vccd1 vccd1 _5256_/A sky130_fd_sc_hd__a211o_1
X_4206_ _4206_/A _4206_/B vssd1 vssd1 vccd1 vccd1 _4206_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4311__B2 _5581_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4167__S _6334_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5186_ _5186_/A _5186_/B vssd1 vssd1 vccd1 vccd1 _5187_/B sky130_fd_sc_hd__xnor2_1
X_4137_ hold190/X hold181/X hold208/X hold105/X _5721_/C1 _5721_/B1 vssd1 vssd1 vccd1
+ vccd1 _4137_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_3_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6064__A1 _4366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4068_ _5136_/A _4068_/B vssd1 vssd1 vccd1 vccd1 _4068_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__4691__A _6089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4866__A _6364_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5461__S _5567_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout161 hold649/X vssd1 vssd1 vccd1 vccd1 _3172_/A sky130_fd_sc_hd__buf_4
Xfanout150 _4675_/A vssd1 vssd1 vccd1 vccd1 _3205_/B sky130_fd_sc_hd__buf_4
Xfanout183 fanout185/X vssd1 vssd1 vccd1 vccd1 fanout183/X sky130_fd_sc_hd__clkbuf_8
Xfanout172 fanout175/X vssd1 vssd1 vccd1 vccd1 fanout172/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3577__C1 _5607_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5318__B1 _5605_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4540__S _4545_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold609 _6468_/Q vssd1 vssd1 vccd1 vccd1 _3501_/A sky130_fd_sc_hd__buf_2
XANTENNA__5869__A1 _5867_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3370_ _3370_/A _3370_/B _3370_/C vssd1 vssd1 vccd1 vccd1 _5617_/B sky130_fd_sc_hd__and3_2
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3680__A _5605_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5040_ _5039_/X _5038_/X _5101_/S vssd1 vssd1 vccd1 vccd1 _5041_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_85_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6046__A1 _5567_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5942_ _5941_/X _5933_/A _5975_/S vssd1 vssd1 vccd1 vccd1 _5942_/X sky130_fd_sc_hd__mux2_1
X_5873_ _5976_/S _5884_/B _5872_/X _5865_/X vssd1 vssd1 vccd1 vccd1 _5873_/X sky130_fd_sc_hd__a31o_1
X_4824_ _5064_/A _4835_/B vssd1 vssd1 vccd1 vccd1 _4824_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__5557__A0 _6461_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4755_ _6314_/Q _4719_/A _4754_/X _4957_/S vssd1 vssd1 vccd1 vccd1 _4755_/X sky130_fd_sc_hd__a22o_1
X_3706_ _5294_/A _6346_/Q _5247_/S _3705_/Y vssd1 vssd1 vccd1 vccd1 _4670_/C sky130_fd_sc_hd__o31a_2
XANTENNA__3583__A2 _3581_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4686_ _6380_/Q _6286_/Q _4711_/S vssd1 vssd1 vccd1 vccd1 _4686_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3637_ _6457_/Q _3506_/B _3638_/C _3464_/A vssd1 vssd1 vccd1 vccd1 _3637_/X sky130_fd_sc_hd__o211a_1
X_6425_ _6428_/CLK _6425_/D fanout171/X vssd1 vssd1 vccd1 vccd1 _6425_/Q sky130_fd_sc_hd__dfrtp_4
X_3568_ _5317_/B _3569_/B vssd1 vssd1 vccd1 vccd1 _4264_/C sky130_fd_sc_hd__nor2_1
X_6356_ _6481_/CLK _6356_/D vssd1 vssd1 vccd1 vccd1 _6356_/Q sky130_fd_sc_hd__dfxtp_1
X_5307_ _5345_/C _5523_/A _5307_/C _5346_/C vssd1 vssd1 vccd1 vccd1 _5311_/B sky130_fd_sc_hd__or4_1
XFILLER_0_59_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5281__S _5292_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6287_ _6465_/CLK _6287_/D vssd1 vssd1 vccd1 vccd1 _6287_/Q sky130_fd_sc_hd__dfxtp_4
X_3499_ _5384_/A _5567_/B vssd1 vssd1 vccd1 vccd1 _5600_/C sky130_fd_sc_hd__nor2_1
X_5238_ _5123_/Y _5126_/Y _6279_/Q _4555_/Y vssd1 vssd1 vccd1 vccd1 _5239_/B sky130_fd_sc_hd__o2bb2a_1
X_5169_ _6335_/Q _5168_/X _5284_/S vssd1 vssd1 vccd1 vccd1 _5169_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4048__B1 _3801_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4599__A1 _3172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_40_wb_clk_i_A clkbuf_leaf_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5548__A0 _6460_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_30_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6419_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__5720__B1 _5721_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6 hold6/A vssd1 vssd1 vccd1 vccd1 hold6/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6028__A1 _5478_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4535__S _4536_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5003__A2 _4963_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4540_ hold264/X _4428_/X _4545_/S vssd1 vssd1 vccd1 vccd1 _6251_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_40_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6051__A _6085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold406 _5393_/X vssd1 vssd1 vccd1 vccd1 _6354_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold417 _6475_/Q vssd1 vssd1 vccd1 vccd1 hold417/X sky130_fd_sc_hd__dlygate4sd3_1
X_4471_ hold187/X _4138_/X _4473_/S vssd1 vssd1 vccd1 vccd1 _4471_/X sky130_fd_sc_hd__mux2_1
X_3422_ _3590_/A _3674_/A _3409_/Y _3281_/X _3421_/Y vssd1 vssd1 vccd1 vccd1 _3424_/C
+ sky130_fd_sc_hd__a221o_1
Xhold439 _4566_/X vssd1 vssd1 vccd1 vccd1 _6273_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6210_ _6449_/CLK _6210_/D vssd1 vssd1 vccd1 vccd1 _6210_/Q sky130_fd_sc_hd__dfxtp_1
Xhold428 _5077_/X vssd1 vssd1 vccd1 vccd1 _6330_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5711__B1 _5710_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3722__C1 _4948_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6141_ _6393_/CLK _6141_/D vssd1 vssd1 vccd1 vccd1 _6141_/Q sky130_fd_sc_hd__dfxtp_1
X_3353_ _3691_/B _5405_/B _4251_/B vssd1 vssd1 vccd1 vccd1 _3353_/X sky130_fd_sc_hd__a21o_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3284_ _4782_/A _3284_/B _4325_/C vssd1 vssd1 vccd1 vccd1 _3285_/D sky130_fd_sc_hd__or3_2
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6072_ hold578/X _6040_/Y _6071_/X _4366_/A vssd1 vssd1 vccd1 vccd1 _6482_/D sky130_fd_sc_hd__o22a_1
XFILLER_0_29_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5023_ _6486_/Q _5104_/A2 _5022_/X vssd1 vssd1 vccd1 vccd1 _5023_/X sky130_fd_sc_hd__a21o_1
XANTENNA__6019__A1 hold628/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5130__A _6021_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5778__B1 _5322_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5925_ _6405_/Q _6424_/Q _5971_/S vssd1 vssd1 vccd1 vccd1 _5925_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5856_ _5855_/A _5855_/B _5854_/X vssd1 vssd1 vccd1 vccd1 _5872_/B sky130_fd_sc_hd__o21ba_1
XFILLER_0_90_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4807_ _4264_/B _4676_/B _4806_/X vssd1 vssd1 vccd1 vccd1 _5108_/S sky130_fd_sc_hd__a21o_4
XFILLER_0_61_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5787_ _6361_/Q _6413_/Q _5892_/S vssd1 vssd1 vccd1 vccd1 _5787_/X sky130_fd_sc_hd__mux2_1
X_4738_ hold403/X _4303_/C _4768_/S vssd1 vssd1 vccd1 vccd1 _4738_/X sky130_fd_sc_hd__mux2_1
X_4669_ hold625/X _4652_/X _4654_/Y _4668_/X vssd1 vssd1 vccd1 vccd1 _6300_/D sky130_fd_sc_hd__o22a_1
XFILLER_0_43_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_7_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6408_ _6426_/CLK _6408_/D fanout171/X vssd1 vssd1 vccd1 vccd1 _6408_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_0_12_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6339_ _6465_/CLK _6339_/D fanout185/X vssd1 vssd1 vccd1 vccd1 _6339_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_0_98_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4992__A1 _6422_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5941__A0 _6462_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6376__RESET_B fanout172/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6305__RESET_B fanout183/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4275__A3 _5317_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3483__B2 _5995_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3971_ _5136_/A _3973_/A vssd1 vssd1 vccd1 vccd1 _3971_/Y sky130_fd_sc_hd__nand2_1
X_5710_ _4447_/X _5706_/X _4137_/X _5709_/X _5655_/B _5734_/S vssd1 vssd1 vccd1 vccd1
+ _5710_/X sky130_fd_sc_hd__mux4_2
XANTENNA__4983__A1 _6310_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5527__A3 _5525_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5641_ _5734_/S _5638_/X _5640_/X _5632_/Y vssd1 vssd1 vccd1 vccd1 _5641_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_72_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3538__A2 _3352_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5572_ _5594_/A _5573_/B vssd1 vssd1 vccd1 vccd1 _5574_/A sky130_fd_sc_hd__nand2_1
X_4523_ _4435_/X hold201/X _4527_/S vssd1 vssd1 vccd1 vccd1 _4523_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_5_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold203 _6213_/Q vssd1 vssd1 vccd1 vccd1 hold203/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold214 _6180_/Q vssd1 vssd1 vccd1 vccd1 hold214/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold225 _4504_/X vssd1 vssd1 vccd1 vccd1 _6212_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold247 _6358_/Q vssd1 vssd1 vccd1 vccd1 _3390_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold258 _6162_/Q vssd1 vssd1 vccd1 vccd1 _3554_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold236 _6181_/Q vssd1 vssd1 vccd1 vccd1 hold236/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold269 _4466_/X vssd1 vssd1 vccd1 vccd1 _6178_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4454_ hold31/X _4462_/A2 _4463_/S vssd1 vssd1 vccd1 vccd1 _4454_/X sky130_fd_sc_hd__o21a_1
X_3405_ _3405_/A _3405_/B vssd1 vssd1 vccd1 vccd1 _3440_/A sky130_fd_sc_hd__and2_1
XFILLER_0_0_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4385_ hold121/X _4240_/X _4385_/S vssd1 vssd1 vccd1 vccd1 _4385_/X sky130_fd_sc_hd__mux2_1
X_3336_ _3336_/A _3336_/B _3336_/C vssd1 vssd1 vccd1 vccd1 _4802_/B sky130_fd_sc_hd__nand3_4
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6124_ _6422_/CLK _6124_/D fanout173/X vssd1 vssd1 vccd1 vccd1 _6124_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6055_ _6089_/A _6071_/S vssd1 vssd1 vccd1 vccd1 _6055_/Y sky130_fd_sc_hd__nor2_1
X_3267_ _5387_/B _3268_/B vssd1 vssd1 vccd1 vccd1 _5323_/B sky130_fd_sc_hd__nor2_2
X_5006_ _5002_/B _5005_/X _5106_/S vssd1 vssd1 vccd1 vccd1 _5006_/X sky130_fd_sc_hd__mux2_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3198_ _6300_/Q _6299_/Q vssd1 vssd1 vccd1 vccd1 _3514_/B sky130_fd_sc_hd__nand2b_2
XFILLER_0_95_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4903__S _5105_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5908_ _5976_/S _5903_/Y _5907_/X _5786_/Y vssd1 vssd1 vccd1 vccd1 _5908_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_8_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5839_ _5839_/A _5839_/B _5837_/X vssd1 vssd1 vccd1 vccd1 _5840_/B sky130_fd_sc_hd__or3b_1
XANTENNA__4204__A _5268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4821__S1 _5404_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5734__S _5734_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4577__C _5317_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4257__A3 _5317_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5678__C1 _3909_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4170_ _6290_/Q _3770_/A _5263_/A _4115_/A _3979_/A vssd1 vssd1 vccd1 vccd1 _4170_/X
+ sky130_fd_sc_hd__a221o_1
X_3121_ _3205_/B _3249_/A _3167_/B vssd1 vssd1 vccd1 vccd1 _3497_/B sky130_fd_sc_hd__and3_2
XFILLER_0_93_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4879__S1 _5100_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3954_ _3951_/X _3952_/X _5655_/A _4441_/S vssd1 vssd1 vccd1 vccd1 _3954_/X sky130_fd_sc_hd__a22o_2
XFILLER_0_85_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3885_ _3885_/A _3885_/B vssd1 vssd1 vccd1 vccd1 _3885_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__6103__A2_N _6107_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5624_ _5624_/A _5624_/B _5624_/C _5624_/D vssd1 vssd1 vccd1 vccd1 _5624_/X sky130_fd_sc_hd__or4_1
X_5555_ hold556/X _5520_/B _5554_/Y _5415_/X vssd1 vssd1 vccd1 vccd1 _5555_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_77_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5486_ hold601/X input8/X _5510_/S vssd1 vssd1 vccd1 vccd1 _5486_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_13_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4506_ _4441_/X hold249/X _4509_/S vssd1 vssd1 vccd1 vccd1 _6214_/D sky130_fd_sc_hd__mux2_1
XANTENNA__5133__B2 _4957_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4437_ _4437_/A _4437_/B vssd1 vssd1 vccd1 vccd1 _5301_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_1_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6107_ _4227_/X _6106_/X _6107_/S vssd1 vssd1 vccd1 vccd1 _6107_/X sky130_fd_sc_hd__mux2_1
X_4368_ _4546_/A _4400_/A vssd1 vssd1 vccd1 vccd1 _4376_/S sky130_fd_sc_hd__nor2_4
XANTENNA__4892__A0 _6365_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3319_ _5387_/A _5314_/S vssd1 vssd1 vccd1 vccd1 _3379_/A sky130_fd_sc_hd__or2_2
X_4299_ _4296_/A _4298_/X _5232_/S vssd1 vssd1 vccd1 vccd1 _4299_/X sky130_fd_sc_hd__mux2_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6038_ _6101_/B _6036_/X _6101_/A vssd1 vssd1 vccd1 vccd1 _6039_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_96_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4947__A1 _6368_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3757__B _4150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4175__A2 _6464_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4109__A _6289_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5212__B _6460_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4543__S _4545_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5866__C _5866_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5038__S1 _5078_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3670_ _4268_/A _5369_/D vssd1 vssd1 vccd1 vccd1 _3670_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__5882__B _5970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5340_ _6297_/Q _5317_/B _5323_/A vssd1 vssd1 vccd1 vccd1 _5340_/X sky130_fd_sc_hd__o21a_1
X_5271_ _5259_/X _5266_/X _5270_/X _5202_/A _3368_/S vssd1 vssd1 vccd1 vccd1 _5271_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_50_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4222_ _6385_/Q _5374_/C vssd1 vssd1 vccd1 vccd1 _5199_/A sky130_fd_sc_hd__and2_1
XANTENNA__3677__A1 _3674_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4153_ _4157_/B _4153_/B vssd1 vssd1 vccd1 vccd1 _4155_/A sky130_fd_sc_hd__nor2_1
X_3104_ _6300_/Q _6299_/Q _4273_/A vssd1 vssd1 vccd1 vccd1 _3247_/A sky130_fd_sc_hd__or3b_2
X_4084_ hold213/X hold103/X hold204/X hold177/X _5721_/C1 _4235_/S vssd1 vssd1 vccd1
+ vccd1 _4084_/X sky130_fd_sc_hd__mux4_1
XANTENNA__5122__B wire92/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5549__S _5581_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout150_A _4675_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4986_ _4982_/B _4985_/X _5106_/S vssd1 vssd1 vccd1 vccd1 _4986_/X sky130_fd_sc_hd__mux2_1
X_3937_ _5260_/A _5170_/B _5162_/B _3979_/A vssd1 vssd1 vccd1 vccd1 _3938_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_46_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3868_ _3892_/A _3892_/B vssd1 vssd1 vccd1 vccd1 _5300_/C sky130_fd_sc_hd__nand2_1
XANTENNA__5354__A1 _5757_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5607_ _3699_/A _5604_/X _5606_/X _5607_/B2 vssd1 vssd1 vccd1 vccd1 _5608_/B sky130_fd_sc_hd__a22o_1
X_3799_ _3884_/S _3818_/C vssd1 vssd1 vccd1 vccd1 _3799_/X sky130_fd_sc_hd__and2_2
XFILLER_0_33_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5538_ _5517_/B _5531_/B _5531_/A vssd1 vssd1 vccd1 vccd1 _5538_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__5657__A2 _4406_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5469_ _5455_/B _5457_/B _5455_/A vssd1 vssd1 vccd1 vccd1 _5470_/B sky130_fd_sc_hd__a21bo_1
XANTENNA__4960__S0 _5100_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout63_A _5874_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold627_A _6464_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5459__S _5485_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6480__SET_B fanout175/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5042__B1 _5041_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput18 rst_n vssd1 vssd1 vccd1 vccd1 input18/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__5896__A2 _5771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5207__B _6462_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3371__A3 _5617_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4538__S _4545_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5281__A0 _6067_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4840_ _4839_/X hold367/X _5098_/S vssd1 vssd1 vccd1 vccd1 _4840_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_74_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4771_ hold629/X _4770_/X _5232_/S vssd1 vssd1 vccd1 vccd1 _6316_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_7_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3722_ _5295_/A _3711_/Y _5296_/B _4948_/S vssd1 vssd1 vccd1 vccd1 _3722_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_99_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6441_ _6441_/CLK _6441_/D fanout185/X vssd1 vssd1 vccd1 vccd1 _6441_/Q sky130_fd_sc_hd__dfrtp_1
X_3653_ _6023_/A _6022_/A _5770_/C _3374_/Y hold491/X vssd1 vssd1 vccd1 vccd1 _3653_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_43_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6372_ _6376_/CLK _6372_/D fanout172/X vssd1 vssd1 vccd1 vccd1 _6372_/Q sky130_fd_sc_hd__dfrtp_4
X_5323_ _5323_/A _5323_/B _5323_/C _5323_/D vssd1 vssd1 vccd1 vccd1 _5323_/X sky130_fd_sc_hd__or4_1
X_3584_ _3581_/B _4386_/A _3643_/B _4338_/A vssd1 vssd1 vccd1 vccd1 _3584_/X sky130_fd_sc_hd__a211o_1
X_5254_ hold598/X _5253_/Y _5489_/S vssd1 vssd1 vccd1 vccd1 _6338_/D sky130_fd_sc_hd__mux2_1
X_4205_ _5268_/A _5194_/A _4205_/S vssd1 vssd1 vccd1 vccd1 _4206_/B sky130_fd_sc_hd__mux2_1
X_5185_ _5185_/A _5185_/B vssd1 vssd1 vccd1 vccd1 _5186_/B sky130_fd_sc_hd__xnor2_1
X_4136_ hold21/X _4462_/A2 _4463_/S vssd1 vssd1 vccd1 vccd1 _4136_/X sky130_fd_sc_hd__o21a_1
X_4067_ _4064_/X _4065_/X _4066_/Y vssd1 vssd1 vccd1 vccd1 _4067_/X sky130_fd_sc_hd__o21a_1
XANTENNA__4075__B2 _6382_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_30_wb_clk_i_A clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_3_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4691__B _4714_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3588__A _4276_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5024__A0 _6424_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4183__S _4241_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6242__RESET_B fanout180/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4969_ _4988_/B _4969_/B vssd1 vssd1 vccd1 vccd1 _4969_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_46_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout140 _4354_/A vssd1 vssd1 vccd1 vccd1 _5105_/S sky130_fd_sc_hd__buf_6
Xfanout151 _4675_/A vssd1 vssd1 vccd1 vccd1 _3547_/B sky130_fd_sc_hd__buf_2
Xfanout162 hold650/X vssd1 vssd1 vccd1 vccd1 _5268_/A sky130_fd_sc_hd__buf_4
Xfanout173 fanout175/X vssd1 vssd1 vccd1 vccd1 fanout173/X sky130_fd_sc_hd__clkbuf_8
Xfanout184 fanout185/X vssd1 vssd1 vccd1 vccd1 fanout184/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__5978__A _5995_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5566__B2 _5485_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6338__SET_B fanout183/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3592__A3 _5777_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4122__A _6097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5646__A_N _5644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5941_ _6462_/Q _5940_/X _5974_/S vssd1 vssd1 vccd1 vccd1 _5941_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3201__A _5995_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5006__A0 _5002_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_0_wb_clk_i clkbuf_leaf_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6455_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_5872_ _5872_/A _5872_/B _5870_/X vssd1 vssd1 vccd1 vccd1 _5872_/X sky130_fd_sc_hd__or3b_1
X_4823_ _5101_/S _4821_/X _4820_/Y vssd1 vssd1 vccd1 vccd1 _4835_/B sky130_fd_sc_hd__o21ai_2
XFILLER_0_28_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4754_ _6314_/Q _4720_/X _5224_/A2 hold454/X vssd1 vssd1 vccd1 vccd1 _4754_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_7_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3705_ _5294_/A _4713_/A vssd1 vssd1 vccd1 vccd1 _3705_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_55_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4685_ _4715_/B2 _4681_/Y _4684_/X hold334/X _4672_/Y vssd1 vssd1 vccd1 vccd1 _4685_/X
+ sky130_fd_sc_hd__o32a_1
XANTENNA__4780__A2 _5413_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3574__C _5146_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3636_ _4800_/S _3636_/B _3636_/C vssd1 vssd1 vccd1 vccd1 _3638_/C sky130_fd_sc_hd__or3_2
XANTENNA_fanout113_A _6108_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6424_ _6426_/CLK _6424_/D fanout171/X vssd1 vssd1 vccd1 vccd1 _6424_/Q sky130_fd_sc_hd__dfrtp_4
X_3567_ _4325_/C _3567_/B _3567_/C vssd1 vssd1 vccd1 vccd1 _3567_/X sky130_fd_sc_hd__and3_1
X_6355_ _6377_/CLK _6355_/D vssd1 vssd1 vccd1 vccd1 _6355_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_11_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5306_ _3205_/B _4335_/C _3305_/A _5371_/A vssd1 vssd1 vccd1 vccd1 _5346_/C sky130_fd_sc_hd__a211o_1
X_6286_ _6441_/CLK _6286_/D vssd1 vssd1 vccd1 vccd1 _6286_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_59_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3590__B _5317_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5237_ _4716_/A _5125_/Y _5132_/B _6337_/Q _4719_/Y vssd1 vssd1 vccd1 vccd1 _5237_/X
+ sky130_fd_sc_hd__a311o_1
X_3498_ _4363_/A _3699_/A _3497_/B _5567_/B vssd1 vssd1 vccd1 vccd1 _3503_/A sky130_fd_sc_hd__a31o_1
XFILLER_0_11_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5168_ _4156_/A _5159_/Y _5166_/Y _5167_/X vssd1 vssd1 vccd1 vccd1 _5168_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_75_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4119_ _3979_/A _5257_/B _4113_/X _4118_/X vssd1 vssd1 vccd1 vccd1 _4119_/X sky130_fd_sc_hd__a211o_1
X_5099_ _6158_/Q _6149_/Q _6141_/Q _6185_/Q _5100_/S0 _5100_/S1 vssd1 vssd1 vccd1
+ vccd1 _5099_/X sky130_fd_sc_hd__mux4_1
XANTENNA__4599__A2 _4324_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4207__A _5268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3559__B1 _5387_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6033__D_N _4670_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5472__S _5485_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5484__A0 _5605_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold7 hold7/A vssd1 vssd1 vccd1 vccd1 hold7/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3378__D _5317_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4551__S _4554_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3970__B1 _6286_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold418 _6044_/X vssd1 vssd1 vccd1 vccd1 _6475_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4470_ hold157/X _4085_/X _4473_/S vssd1 vssd1 vccd1 vccd1 _4470_/X sky130_fd_sc_hd__mux2_1
Xhold407 _6405_/Q vssd1 vssd1 vccd1 vccd1 hold407/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3421_ _4289_/B _5316_/B vssd1 vssd1 vccd1 vccd1 _3421_/Y sky130_fd_sc_hd__nor2_1
Xhold429 _6381_/Q vssd1 vssd1 vccd1 vccd1 _4027_/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5711__A1 _6463_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3352_ _4338_/A _3352_/B vssd1 vssd1 vccd1 vccd1 _5405_/B sky130_fd_sc_hd__or2_1
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6140_ _6239_/CLK _6140_/D vssd1 vssd1 vccd1 vccd1 _6140_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3283_ _4386_/A _5405_/A _3587_/B vssd1 vssd1 vccd1 vccd1 _3355_/C sky130_fd_sc_hd__and3_1
XANTENNA__5475__A0 _6462_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6071_ _4227_/X _6070_/Y _6071_/S vssd1 vssd1 vccd1 vccd1 _6071_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_29_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5022_ _6312_/Q _4963_/B _5021_/B _4796_/Y vssd1 vssd1 vccd1 vccd1 _5022_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4726__S _4768_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5411__A _5757_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5130__B _5783_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5924_ _5924_/A _5924_/B vssd1 vssd1 vccd1 vccd1 _5924_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5855_ _5855_/A _5855_/B _5854_/X vssd1 vssd1 vccd1 vccd1 _5857_/A sky130_fd_sc_hd__nor3b_1
X_4806_ _4806_/A _4806_/B _4806_/C _4806_/D vssd1 vssd1 vccd1 vccd1 _4806_/X sky130_fd_sc_hd__and4_1
XFILLER_0_75_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5786_ _5786_/A _5786_/B vssd1 vssd1 vccd1 vccd1 _5786_/Y sky130_fd_sc_hd__nor2_4
XFILLER_0_16_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4737_ _6311_/Q _4719_/A _4736_/X _4957_/S vssd1 vssd1 vccd1 vccd1 _4737_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_43_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4668_ _4668_/A _4668_/B vssd1 vssd1 vccd1 vccd1 _4668_/X sky130_fd_sc_hd__and2_1
XFILLER_0_16_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3619_ _5322_/A _5345_/C _3619_/C _5372_/B vssd1 vssd1 vccd1 vccd1 _3619_/X sky130_fd_sc_hd__or4_1
X_6407_ _6407_/CLK _6407_/D fanout170/X vssd1 vssd1 vccd1 vccd1 _6407_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__5292__S _5292_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4599_ _3172_/A _4324_/B _4592_/X _4597_/X vssd1 vssd1 vccd1 vccd1 _4611_/B sky130_fd_sc_hd__a211o_2
XFILLER_0_101_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6338_ _6340_/CLK _6338_/D fanout183/X vssd1 vssd1 vccd1 vccd1 _6338_/Q sky130_fd_sc_hd__dfstp_2
X_6269_ _6312_/CLK _6269_/D fanout182/X vssd1 vssd1 vccd1 vccd1 _6269_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_0_79_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4371__S _4376_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3952__B1 _4463_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5930__S _5976_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4680__A1 _4715_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3970_ _3972_/B _3972_/C _6286_/Q vssd1 vssd1 vccd1 vccd1 _3973_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_97_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4983__A2 _4963_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5640_ _3910_/X _5732_/A _5630_/D _5639_/X vssd1 vssd1 vccd1 vccd1 _5640_/X sky130_fd_sc_hd__a211o_1
X_5571_ _6488_/Q _5063_/B _5593_/S vssd1 vssd1 vccd1 vccd1 _5573_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_31_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3943__B1 _3801_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4522_ _4428_/X hold272/X _4527_/S vssd1 vssd1 vccd1 vccd1 _4522_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_80_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold204 _6263_/Q vssd1 vssd1 vccd1 vccd1 hold204/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold226 _6195_/Q vssd1 vssd1 vccd1 vccd1 hold226/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold215 _6193_/Q vssd1 vssd1 vccd1 vccd1 hold215/X sky130_fd_sc_hd__dlygate4sd3_1
X_4453_ _4438_/A _5301_/C _4178_/Y _3701_/B vssd1 vssd1 vccd1 vccd1 _4453_/X sky130_fd_sc_hd__a211o_1
X_3404_ _5777_/A _3404_/B vssd1 vssd1 vccd1 vccd1 _3405_/B sky130_fd_sc_hd__nor2_1
XANTENNA__5406__A _5777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold248 _5401_/X vssd1 vssd1 vccd1 vccd1 _6358_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold259 _3554_/X vssd1 vssd1 vccd1 vccd1 _6162_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold237 _6111_/Q vssd1 vssd1 vccd1 vccd1 hold237/X sky130_fd_sc_hd__dlygate4sd3_1
X_4384_ hold114/X _4182_/X _4385_/S vssd1 vssd1 vccd1 vccd1 _4384_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3171__A1 _4273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3335_ _3310_/Y _3317_/X _3329_/X _3334_/X _3298_/X vssd1 vssd1 vccd1 vccd1 _3336_/C
+ sky130_fd_sc_hd__a41o_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6123_ _6419_/CLK _6123_/D fanout173/X vssd1 vssd1 vccd1 vccd1 _6123_/Q sky130_fd_sc_hd__dfrtp_1
X_3266_ _4260_/B _3268_/B vssd1 vssd1 vccd1 vccd1 _5146_/B sky130_fd_sc_hd__or2_2
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6054_ _6101_/A _6053_/X _6071_/S vssd1 vssd1 vccd1 vccd1 _6054_/X sky130_fd_sc_hd__o21a_1
XANTENNA__3459__C1 _5995_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4120__A0 _6463_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5999__B2 _5995_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5005_ _6423_/Q _6371_/Q _5105_/S vssd1 vssd1 vccd1 vccd1 _5005_/X sky130_fd_sc_hd__mux2_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3197_ _6300_/Q _6299_/Q vssd1 vssd1 vccd1 vccd1 _5360_/A sky130_fd_sc_hd__and2b_2
XANTENNA_fanout180_A input18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5907_ _6459_/Q _5906_/X _5974_/S vssd1 vssd1 vccd1 vccd1 _5907_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4423__A1 _5730_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5838_ _5839_/A _5839_/B _5837_/X vssd1 vssd1 vccd1 vccd1 _5855_/B sky130_fd_sc_hd__o21ba_1
XFILLER_0_36_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4204__B _6290_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5769_ hold19/X _4283_/Y _5769_/S vssd1 vssd1 vccd1 vccd1 hold20/A sky130_fd_sc_hd__mux2_1
XFILLER_0_8_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5923__A1 _6423_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4187__B1 _3807_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5316__A _5364_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4220__A _6385_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout93_A _5016_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5750__S _6104_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5611__B1 _4300_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3925__A0 _6379_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3120_ _3284_/B _3172_/A _4782_/A vssd1 vssd1 vccd1 vccd1 _3639_/C sky130_fd_sc_hd__nand3b_4
XANTENNA__4766__A2_N _4720_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4102__B1 _5268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5850__A0 _6366_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5602__B1 _5362_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3953_ hold226/X hold91/X hold239/X hold161/X _5721_/C1 _4235_/S vssd1 vssd1 vccd1
+ vccd1 _5655_/A sky130_fd_sc_hd__mux4_1
XFILLER_0_18_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3884_ hold126/X hold75/X _3884_/S vssd1 vssd1 vccd1 vccd1 _3885_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_18_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4169__A0 _6289_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5623_ _5522_/D _5618_/X _5622_/X _5777_/A vssd1 vssd1 vccd1 vccd1 _5624_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_5_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5554_ _5554_/A vssd1 vssd1 vccd1 vccd1 _5554_/Y sky130_fd_sc_hd__inv_2
X_5485_ _5483_/X _5484_/X _5485_/S vssd1 vssd1 vccd1 vccd1 _5485_/X sky130_fd_sc_hd__mux2_1
X_4505_ _4435_/X hold203/X _4509_/S vssd1 vssd1 vccd1 vccd1 _6213_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_41_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4436_ hold118/X _4435_/X _4464_/S vssd1 vssd1 vccd1 vccd1 _4436_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_6_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4367_ _5769_/S _5078_/S1 _4802_/D _4366_/X vssd1 vssd1 vccd1 vccd1 _6129_/D sky130_fd_sc_hd__o22a_1
XFILLER_0_6_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3318_ _5387_/A _5314_/S vssd1 vssd1 vccd1 vccd1 _3396_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_67_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3695__A2 _5418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5570__S _5581_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6106_ hold594/X _6039_/A _6105_/X _6101_/A vssd1 vssd1 vccd1 vccd1 _6106_/X sky130_fd_sc_hd__o22a_1
X_4298_ _6310_/Q _4322_/B _4296_/X _4300_/B vssd1 vssd1 vccd1 vccd1 _4298_/X sky130_fd_sc_hd__a22o_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3249_ _3249_/A _3249_/B vssd1 vssd1 vccd1 vccd1 _4344_/A sky130_fd_sc_hd__nand2_4
X_6037_ _6070_/A _6037_/B vssd1 vssd1 vccd1 vccd1 _6037_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__5841__A0 _6365_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5745__S _6104_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold590 _6367_/Q vssd1 vssd1 vccd1 vccd1 hold590/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4635__B2 _4634_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4399__B1 _5384_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5270_ _5171_/A _5171_/B _5261_/X _5269_/X vssd1 vssd1 vccd1 vccd1 _5270_/X sky130_fd_sc_hd__o31a_1
XFILLER_0_2_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4221_ _3740_/B _3364_/Y _3761_/B _4220_/X vssd1 vssd1 vccd1 vccd1 _4221_/X sky130_fd_sc_hd__o211a_1
XANTENNA__4874__A1 _6364_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4152_ _6290_/Q _4152_/B vssd1 vssd1 vccd1 vccd1 _4153_/B sky130_fd_sc_hd__nor2_1
X_3103_ _6300_/Q _6299_/Q vssd1 vssd1 vccd1 vccd1 _3183_/A sky130_fd_sc_hd__or2_1
X_4083_ hold25/X _4462_/A2 _4463_/S vssd1 vssd1 vccd1 vccd1 _4083_/X sky130_fd_sc_hd__o21a_1
XANTENNA_clkbuf_leaf_20_wb_clk_i_A _6448_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4734__S _4770_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5051__A1 _6425_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4985_ _6422_/Q _6370_/Q _5105_/S vssd1 vssd1 vccd1 vccd1 _4985_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_92_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3936_ _4107_/B _4016_/A _6285_/Q vssd1 vssd1 vccd1 vccd1 _5170_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_73_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3867_ _3864_/Y _3866_/Y _3816_/B _3862_/X vssd1 vssd1 vccd1 vccd1 _3892_/B sky130_fd_sc_hd__a2bb2o_2
XANTENNA__6448__RESET_B fanout185/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5354__A2 _4150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5606_ _5777_/A _3278_/A _4326_/Y _4595_/B _5605_/X vssd1 vssd1 vccd1 vccd1 _5606_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_61_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3798_ _3714_/X _3717_/Y _3718_/X _3723_/Y vssd1 vssd1 vccd1 vccd1 _3818_/C sky130_fd_sc_hd__o211a_2
XFILLER_0_5_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5537_ hold391/X _5536_/X _5581_/S vssd1 vssd1 vccd1 vccd1 _5537_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_14_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5468_ _5468_/A _5468_/B vssd1 vssd1 vccd1 vccd1 _5470_/A sky130_fd_sc_hd__and2_1
X_5399_ _3527_/C _5398_/X hold315/X vssd1 vssd1 vccd1 vccd1 _6357_/D sky130_fd_sc_hd__a21oi_1
X_4419_ hold189/X _4408_/S _5731_/C1 _4418_/X vssd1 vssd1 vccd1 vccd1 _4419_/X sky130_fd_sc_hd__o211a_1
XANTENNA__4960__S1 _5100_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4617__A1 _6460_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4617__B2 _6311_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3840__A2 _3793_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5042__A1 _6313_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_24_wb_clk_i _6448_/CLK vssd1 vssd1 vccd1 vccd1 _6465_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_91_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3784__A _4675_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4608__A1 _6458_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4608__B2 _6309_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output37_A _6330_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4736__A1_N _6311_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3136__D_N _3168_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3292__B1 _3668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4554__S _4554_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4770_ _4227_/X _4769_/X _4770_/S vssd1 vssd1 vccd1 vccd1 _4770_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_70_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3721_ hold19/A _3700_/Y _4441_/S vssd1 vssd1 vccd1 vccd1 _3721_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_28_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3652_ _5522_/A _3652_/B _5388_/A _4595_/B vssd1 vssd1 vccd1 vccd1 _5770_/C sky130_fd_sc_hd__and4_1
XFILLER_0_70_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6440_ _6467_/CLK _6440_/D fanout177/X vssd1 vssd1 vccd1 vccd1 _6440_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__6070__A _6070_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3583_ _4313_/A _3581_/B _3643_/B _5218_/S vssd1 vssd1 vccd1 vccd1 _5367_/B sky130_fd_sc_hd__o31a_1
X_6371_ _6376_/CLK _6371_/D fanout172/X vssd1 vssd1 vccd1 vccd1 _6371_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_23_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5322_ _5322_/A _5322_/B vssd1 vssd1 vccd1 vccd1 _5322_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_11_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5253_ _5253_/A vssd1 vssd1 vccd1 vccd1 _5253_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4729__S _5232_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4204_ _5268_/A _6290_/Q vssd1 vssd1 vccd1 vccd1 _5194_/A sky130_fd_sc_hd__xor2_1
X_5184_ _5262_/C _5262_/D vssd1 vssd1 vccd1 vccd1 _5185_/B sky130_fd_sc_hd__xor2_1
X_4135_ _4438_/A _5304_/A _4123_/Y vssd1 vssd1 vccd1 vccd1 _4135_/X sky130_fd_sc_hd__a21o_1
X_4066_ _4064_/X _4065_/X _4156_/A vssd1 vssd1 vccd1 vccd1 _4066_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_78_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4464__S _4464_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4458__S0 _5731_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4968_ _4968_/A _4968_/B vssd1 vssd1 vccd1 vccd1 _4969_/B sky130_fd_sc_hd__and2_1
X_3919_ _3750_/A _3750_/B _3743_/B vssd1 vssd1 vccd1 vccd1 _3921_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_46_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4899_ hold99/A hold67/A _6454_/Q _6231_/Q _5100_/S0 _5100_/S1 vssd1 vssd1 vccd1
+ vccd1 _4899_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_34_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3338__A1 _3489_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout130 hold566/X vssd1 vssd1 vccd1 vccd1 _3489_/B sky130_fd_sc_hd__buf_6
Xfanout152 hold656/X vssd1 vssd1 vccd1 vccd1 _4675_/A sky130_fd_sc_hd__buf_4
Xfanout163 hold604/X vssd1 vssd1 vccd1 vccd1 _4324_/B sky130_fd_sc_hd__clkbuf_8
Xfanout174 fanout175/X vssd1 vssd1 vccd1 vccd1 fanout174/X sky130_fd_sc_hd__buf_4
Xfanout141 _4406_/B vssd1 vssd1 vccd1 vccd1 _5721_/A2 sky130_fd_sc_hd__buf_4
Xfanout185 input18/X vssd1 vssd1 vccd1 vccd1 fanout185/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_88_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4374__S _4376_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5015__A1 _5771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4549__S _4554_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5940_ _5964_/A _5939_/X _5041_/Y vssd1 vssd1 vccd1 vccd1 _5940_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_87_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5871_ _5872_/A _5872_/B _5870_/X vssd1 vssd1 vccd1 vccd1 _5884_/B sky130_fd_sc_hd__o21bai_1
XFILLER_0_34_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4822_ _4919_/S _4821_/X _4820_/Y vssd1 vssd1 vccd1 vccd1 _4822_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_28_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4753_ hold631/X _4752_/X _5232_/S vssd1 vssd1 vccd1 vccd1 _6313_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_50_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3704_ _5146_/A _3704_/B vssd1 vssd1 vccd1 vccd1 _4713_/A sky130_fd_sc_hd__or2_4
XANTENNA__4313__A _4313_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6004__S _6011_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4684_ _4713_/A _4683_/X _4714_/S vssd1 vssd1 vccd1 vccd1 _4684_/X sky130_fd_sc_hd__o21a_1
X_6423_ _6426_/CLK _6423_/D fanout171/X vssd1 vssd1 vccd1 vccd1 _6423_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_31_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3635_ _4800_/S _3636_/B vssd1 vssd1 vccd1 vccd1 _3635_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_3_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3566_ _5345_/A _5522_/D _3564_/X _3228_/C vssd1 vssd1 vccd1 vccd1 _3567_/C sky130_fd_sc_hd__o2bb2a_1
X_6354_ _6441_/CLK _6354_/D fanout184/X vssd1 vssd1 vccd1 vccd1 _6354_/Q sky130_fd_sc_hd__dfrtp_1
X_6285_ _6465_/CLK _6285_/D vssd1 vssd1 vccd1 vccd1 _6285_/Q sky130_fd_sc_hd__dfxtp_4
X_5305_ _3632_/C _5297_/X _5298_/Y _5304_/X vssd1 vssd1 vccd1 vccd1 _5305_/X sky130_fd_sc_hd__a22o_1
X_3497_ _3699_/A _3497_/B vssd1 vssd1 vccd1 vccd1 _5400_/A sky130_fd_sc_hd__and2_1
X_5236_ _6337_/Q _5202_/A _5235_/X _4223_/A vssd1 vssd1 vccd1 vccd1 _5236_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_52_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5493__A1 _5492_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5167_ _5166_/A _5166_/B _4060_/B vssd1 vssd1 vccd1 vccd1 _5167_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_98_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4118_ _4116_/A _3759_/Y _4117_/X _6383_/Q _4115_/X vssd1 vssd1 vccd1 vccd1 _4118_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4048__A2 _3799_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5098_ _5097_/X hold504/X _5098_/S vssd1 vssd1 vccd1 vccd1 _5098_/X sky130_fd_sc_hd__mux2_1
X_4049_ _6222_/Q _3804_/X _3807_/X _6138_/Q vssd1 vssd1 vccd1 vccd1 _4049_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_78_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4453__C1 _3701_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4207__B _6290_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6463__RESET_B fanout181/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5753__S _6104_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5705__C1 _5721_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5720__A2 _5721_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4369__S _4376_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5484__A1 _6366_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold8 hold8/A vssd1 vssd1 vccd1 vccd1 hold8/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5236__A1 _6337_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5928__S _5974_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6133__RESET_B fanout180/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4842__S0 _5404_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3972__A _6286_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold408 _5761_/X vssd1 vssd1 vccd1 vccd1 _6405_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3420_ _5316_/B vssd1 vssd1 vccd1 vccd1 _3420_/Y sky130_fd_sc_hd__inv_2
Xhold419 _6385_/Q vssd1 vssd1 vccd1 vccd1 hold419/X sky130_fd_sc_hd__buf_1
X_3351_ _4276_/A _4325_/A vssd1 vssd1 vccd1 vccd1 _4386_/B sky130_fd_sc_hd__nand2_2
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3282_ _3282_/A _3360_/B _4325_/C vssd1 vssd1 vccd1 vccd1 _3587_/B sky130_fd_sc_hd__or3_2
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6070_ _6070_/A _6070_/B vssd1 vssd1 vccd1 vccd1 _6070_/Y sky130_fd_sc_hd__nand2_1
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5021_ _5102_/A _5021_/B vssd1 vssd1 vccd1 vccd1 _5021_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_31_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5227__A1 _6381_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3212__A _5124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4986__A0 _4982_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5923_ _6423_/Q _5970_/A _5915_/A vssd1 vssd1 vccd1 vccd1 _5924_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_75_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6523__A _6529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5854_ _5872_/A _5854_/B vssd1 vssd1 vccd1 vccd1 _5854_/X sky130_fd_sc_hd__or2_1
X_4805_ _5345_/C _5523_/A vssd1 vssd1 vccd1 vccd1 _4806_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_75_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4202__A2 _5268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5785_ _6023_/A _5976_/S _5977_/S vssd1 vssd1 vccd1 vccd1 _5785_/Y sky130_fd_sc_hd__o21ai_4
X_4736_ _6311_/Q _4720_/X wire92/X hold462/X vssd1 vssd1 vccd1 vccd1 _4736_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_9_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4667_ hold615/X _4652_/X _4654_/Y _4666_/X vssd1 vssd1 vccd1 vccd1 _6299_/D sky130_fd_sc_hd__o22a_1
XFILLER_0_71_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3618_ _4253_/A _3618_/B vssd1 vssd1 vccd1 vccd1 _5372_/B sky130_fd_sc_hd__nand2_1
X_6406_ _6409_/CLK _6406_/D fanout171/X vssd1 vssd1 vccd1 vccd1 _6406_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6337_ _6340_/CLK _6337_/D fanout183/X vssd1 vssd1 vccd1 vccd1 _6337_/Q sky130_fd_sc_hd__dfstp_2
X_4598_ _3172_/A _4324_/B _4592_/X _4597_/X vssd1 vssd1 vccd1 vccd1 _4641_/B sky130_fd_sc_hd__a211oi_4
X_3549_ _5124_/A _5388_/A _4248_/C vssd1 vssd1 vccd1 vccd1 _3549_/X sky130_fd_sc_hd__and3_1
X_6268_ _6316_/CLK _6268_/D fanout174/X vssd1 vssd1 vccd1 vccd1 _6268_/Q sky130_fd_sc_hd__dfstp_1
X_5219_ _3994_/Y _5218_/X _5292_/S vssd1 vssd1 vccd1 vccd1 _5219_/X sky130_fd_sc_hd__mux2_1
X_6199_ _6265_/CLK _6199_/D vssd1 vssd1 vccd1 vccd1 _6199_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5748__S _6104_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4827__S _4948_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5570_ _5567_/A _5569_/X _5581_/S vssd1 vssd1 vccd1 vccd1 _5570_/X sky130_fd_sc_hd__mux2_1
X_4521_ _4416_/X hold292/X _4527_/S vssd1 vssd1 vccd1 vccd1 _4521_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_25_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold205 _4551_/X vssd1 vssd1 vccd1 vccd1 _6263_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4452_ _4459_/B _4452_/B vssd1 vssd1 vccd1 vccd1 _5301_/C sky130_fd_sc_hd__nor2_1
Xhold216 _4482_/X vssd1 vssd1 vccd1 vccd1 _6193_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3403_ _5617_/B _3619_/C vssd1 vssd1 vccd1 vccd1 _3404_/B sky130_fd_sc_hd__nor2_1
Xhold227 _4485_/X vssd1 vssd1 vccd1 vccd1 _6195_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold249 _6214_/Q vssd1 vssd1 vccd1 vccd1 hold249/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold238 _3912_/X vssd1 vssd1 vccd1 vccd1 _6111_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4383_ hold181/X _4138_/X _4385_/S vssd1 vssd1 vccd1 vccd1 _4383_/X sky130_fd_sc_hd__mux2_1
X_3334_ _5370_/C _3334_/B _3334_/C vssd1 vssd1 vccd1 vccd1 _3334_/X sky130_fd_sc_hd__and3b_1
X_6122_ _6417_/CLK _6122_/D fanout174/X vssd1 vssd1 vccd1 vccd1 _6122_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3265_ _4260_/B _3268_/B vssd1 vssd1 vccd1 vccd1 _3278_/B sky130_fd_sc_hd__nor2_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6053_ _6101_/B _4863_/X _5457_/X _6036_/X vssd1 vssd1 vccd1 vccd1 _6053_/X sky130_fd_sc_hd__o22a_1
XANTENNA__5422__A _6019_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5004_ _6485_/Q _5104_/A2 _5003_/X vssd1 vssd1 vccd1 vccd1 _5004_/X sky130_fd_sc_hd__a21o_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3196_ _4359_/C _3196_/B vssd1 vssd1 vccd1 vccd1 _3196_/Y sky130_fd_sc_hd__nand2_1
XANTENNA_fanout173_A fanout175/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5620__A1 _3168_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4472__S _4473_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5906_ _5964_/A _5905_/X _4982_/Y vssd1 vssd1 vccd1 vccd1 _5906_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_76_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5837_ _5855_/A _5837_/B vssd1 vssd1 vccd1 vccd1 _5837_/X sky130_fd_sc_hd__or2_1
XFILLER_0_36_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5768_ hold41/X _5767_/Y _5769_/S vssd1 vssd1 vccd1 vccd1 hold42/A sky130_fd_sc_hd__mux2_1
XANTENNA__5923__A2 _5970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4719_ _4719_/A vssd1 vssd1 vccd1 vccd1 _4719_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_44_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5699_ _6313_/Q _5630_/X _5653_/X _6487_/Q _5698_/X vssd1 vssd1 vccd1 vccd1 _5700_/C
+ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_49_wb_clk_i clkbuf_leaf_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6223_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_31_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3513__A2_N _4248_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4220__B _5374_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold552_A _6425_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4890__B _4930_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5611__A1 _5644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4382__S _4385_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5478__S _5478_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3622__B1 _4653_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3925__A1 _6383_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5941__S _5974_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4350__B2 _5605_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4102__A1 _6289_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_10_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_26_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5602__B2 _4595_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3952_ hold23/X _4462_/A2 _4463_/S vssd1 vssd1 vccd1 vccd1 _3952_/X sky130_fd_sc_hd__o21a_1
X_3883_ _3881_/X _3882_/X _3883_/S vssd1 vssd1 vccd1 vccd1 _3883_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4305__B _5783_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4169__A1 _5268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5622_ _5309_/A _5770_/B _5370_/D _5346_/A vssd1 vssd1 vccd1 vccd1 _5622_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_73_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5553_ _5553_/A _5553_/B vssd1 vssd1 vccd1 vccd1 _5554_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6012__S _6019_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4504_ _4428_/X hold224/X _4509_/S vssd1 vssd1 vccd1 vccd1 _4504_/X sky130_fd_sc_hd__mux2_1
X_5484_ _5605_/C _6366_/Q _5484_/S vssd1 vssd1 vccd1 vccd1 _5484_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_13_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4435_ _4432_/Y _4433_/X _4434_/X _4441_/S vssd1 vssd1 vccd1 vccd1 _4435_/X sky130_fd_sc_hd__a22o_2
XANTENNA__4341__A1 _5607_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4366_ _4366_/A _4366_/B vssd1 vssd1 vccd1 vccd1 _4366_/X sky130_fd_sc_hd__or2_1
XFILLER_0_1_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3317_ _3411_/A _5406_/B _4267_/B vssd1 vssd1 vccd1 vccd1 _3317_/X sky130_fd_sc_hd__and3_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4467__S _4473_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6105_ _6101_/B _5102_/B _5595_/Y _6036_/X vssd1 vssd1 vccd1 vccd1 _6105_/X sky130_fd_sc_hd__o22a_1
X_4297_ _4296_/A _4296_/B _4322_/B vssd1 vssd1 vccd1 vccd1 _4300_/B sky130_fd_sc_hd__a21oi_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6094__A1 _4366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3248_ _4557_/D _3627_/C vssd1 vssd1 vccd1 vccd1 _3307_/B sky130_fd_sc_hd__or2_2
X_6036_ _6036_/A _6036_/B vssd1 vssd1 vccd1 vccd1 _6036_/X sky130_fd_sc_hd__or2_4
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3179_ _3304_/B _3180_/B vssd1 vssd1 vccd1 vccd1 _3570_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_83_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4580__B2 _6159_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5761__S _5765_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold580 _5931_/X vssd1 vssd1 vccd1 vccd1 _6424_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold591 _5501_/X vssd1 vssd1 vccd1 vccd1 _6367_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5062__A _5064_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5832__B2 _5786_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5832__A1 _5976_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3843__B1 _3852_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5001__S _5101_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4571__A1 _6336_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4220_ _6385_/Q _5374_/C vssd1 vssd1 vccd1 vccd1 _4220_/X sky130_fd_sc_hd__or2_1
XANTENNA__4323__A1 _5581_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4323__B2 _6315_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5671__S _5734_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4151_ _6290_/Q _4152_/B vssd1 vssd1 vccd1 vccd1 _4157_/B sky130_fd_sc_hd__and2_1
XANTENNA__4287__S _5769_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3102_ _6300_/Q _6299_/Q vssd1 vssd1 vccd1 vccd1 _3322_/C sky130_fd_sc_hd__nor2_1
X_4082_ _4414_/A _4053_/Y _4081_/X vssd1 vssd1 vccd1 vccd1 _4082_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_37_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5823__A1 _5867_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3834__B1 _3801_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4984_ _6484_/Q _5104_/A2 _4983_/X vssd1 vssd1 vccd1 vccd1 _4984_/X sky130_fd_sc_hd__a21o_1
XANTENNA__6007__S _6011_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3935_ _6287_/Q _6337_/Q vssd1 vssd1 vccd1 vccd1 _4016_/A sky130_fd_sc_hd__or2_1
XFILLER_0_58_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4750__S _4768_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5605_ _5605_/A _5605_/B _5605_/C _5605_/D vssd1 vssd1 vccd1 vccd1 _5605_/X sky130_fd_sc_hd__and4_1
XANTENNA_fanout136_A _4313_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6000__A1 _4653_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3866_ _3885_/A _3865_/X _3852_/A vssd1 vssd1 vccd1 vccd1 _3866_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__5147__A _5292_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3797_ _6259_/Q _4546_/B _4501_/A _6194_/Q vssd1 vssd1 vccd1 vccd1 _3797_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_26_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4562__A1 _6311_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5536_ _6459_/Q _5535_/X _5598_/S vssd1 vssd1 vccd1 vccd1 _5536_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5467_ _5492_/A _5466_/B _5466_/C vssd1 vssd1 vccd1 vccd1 _5468_/B sky130_fd_sc_hd__a21o_1
XANTENNA__5581__S _5581_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4314__A1 _4313_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4418_ hold69/A _6355_/Q _4418_/C vssd1 vssd1 vccd1 vccd1 _4418_/X sky130_fd_sc_hd__or3_1
X_5398_ _5398_/A _5398_/B vssd1 vssd1 vccd1 vccd1 _5398_/X sky130_fd_sc_hd__or2_1
X_4349_ _5603_/A _4343_/X _4348_/X _5522_/A vssd1 vssd1 vccd1 vccd1 _4349_/X sky130_fd_sc_hd__o31a_1
X_6019_ _4668_/A hold628/X _6019_/S vssd1 vssd1 vccd1 vccd1 _6465_/D sky130_fd_sc_hd__mux2_1
XANTENNA__4925__S _5105_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5610__A _5645_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5509__A2_N _5520_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5042__A2 _4963_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5756__S _6104_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4002__B1 _6287_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5491__S _5593_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3720_ _3714_/X _3717_/Y _3718_/X vssd1 vssd1 vccd1 vccd1 _3816_/B sky130_fd_sc_hd__o21ai_4
XFILLER_0_23_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3651_ hold526/X hold1/X _3594_/B vssd1 vssd1 vccd1 vccd1 _6022_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_3_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3582_ _5146_/B _4386_/A _5146_/C _3619_/C _4338_/A vssd1 vssd1 vccd1 vccd1 _5218_/S
+ sky130_fd_sc_hd__a2111o_2
X_6370_ _6488_/CLK _6370_/D fanout172/X vssd1 vssd1 vccd1 vccd1 _6370_/Q sky130_fd_sc_hd__dfrtp_2
X_5321_ _3205_/B _5311_/X _5619_/A _4335_/B vssd1 vssd1 vccd1 vccd1 _5322_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_100_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5252_ _6097_/A _5251_/X _5292_/S vssd1 vssd1 vccd1 vccd1 _5253_/A sky130_fd_sc_hd__mux2_1
X_5183_ _5262_/A _5262_/B vssd1 vssd1 vccd1 vccd1 _5185_/A sky130_fd_sc_hd__xor2_1
X_4203_ _4203_/A _4203_/B vssd1 vssd1 vccd1 vccd1 _4206_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_48_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3215__A _5315_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4134_ _4134_/A _4134_/B vssd1 vssd1 vccd1 vccd1 _5304_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__6049__B2 _6036_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6049__A1 _6101_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4745__S _5289_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4065_ _4007_/A _4007_/B _4005_/A vssd1 vssd1 vccd1 vccd1 _4065_/X sky130_fd_sc_hd__a21o_1
XANTENNA__5272__A2 _5783_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6526__A _6529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4480__S _4482_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4967_ _4968_/A _4968_/B vssd1 vssd1 vccd1 vccd1 _4988_/B sky130_fd_sc_hd__nor2_1
XANTENNA__3885__A _3885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3918_ _3974_/A _3918_/B vssd1 vssd1 vccd1 vccd1 _3921_/A sky130_fd_sc_hd__and2_1
XFILLER_0_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4898_ _6239_/Q _6191_/Q _6175_/Q _6254_/Q _5100_/S0 _5100_/S1 vssd1 vssd1 vccd1
+ vccd1 _4898_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_73_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3849_ _6237_/Q _3884_/S _3848_/X _3883_/S vssd1 vssd1 vccd1 vccd1 _3852_/B sky130_fd_sc_hd__a211o_1
XFILLER_0_6_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3109__B _5605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5519_ _5519_/A _5519_/B vssd1 vssd1 vccd1 vccd1 _5519_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__5605__A _5605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout120 _3057_/Y vssd1 vssd1 vccd1 vccd1 _5605_/A sky130_fd_sc_hd__buf_4
Xfanout131 _4276_/A vssd1 vssd1 vccd1 vccd1 _4335_/B sky130_fd_sc_hd__clkbuf_8
Xfanout153 _4716_/A vssd1 vssd1 vccd1 vccd1 _4217_/A sky130_fd_sc_hd__buf_4
Xfanout164 _5600_/A vssd1 vssd1 vccd1 vccd1 _3699_/A sky130_fd_sc_hd__buf_4
Xfanout142 hold652/X vssd1 vssd1 vccd1 vccd1 _4406_/B sky130_fd_sc_hd__clkbuf_8
Xfanout175 fanout176/X vssd1 vssd1 vccd1 vccd1 fanout175/X sky130_fd_sc_hd__buf_4
XFILLER_0_69_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold632_A _6309_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4390__S _4397_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5971__A0 _6409_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4829__A2 _5108_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4137__S0 _5721_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5870_ _5870_/A _5870_/B vssd1 vssd1 vccd1 vccd1 _5870_/X sky130_fd_sc_hd__or2_1
X_4821_ _6203_/Q _6450_/Q _6211_/Q _6227_/Q _5078_/S1 _5404_/A0 vssd1 vssd1 vccd1
+ vccd1 _4821_/X sky130_fd_sc_hd__mux4_2
XFILLER_0_68_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4752_ _4080_/Y _4751_/X _4770_/S vssd1 vssd1 vccd1 vccd1 _4752_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5962__A0 _6408_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6081__A _6081_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3703_ _6345_/Q _6343_/Q _4150_/A vssd1 vssd1 vccd1 vccd1 _5247_/S sky130_fd_sc_hd__nand3_4
X_4683_ _6383_/Q _4682_/X _4712_/S vssd1 vssd1 vccd1 vccd1 _4683_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_50_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3634_ _5980_/A _3634_/B vssd1 vssd1 vccd1 vccd1 _3636_/C sky130_fd_sc_hd__nand2_1
X_6422_ _6422_/CLK _6422_/D fanout170/X vssd1 vssd1 vccd1 vccd1 _6422_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_70_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3565_ _4557_/C _3333_/C _3320_/Y _3563_/X _4338_/B vssd1 vssd1 vccd1 vccd1 _3567_/B
+ sky130_fd_sc_hd__o32a_1
XFILLER_0_59_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6353_ _6474_/CLK _6353_/D fanout179/X vssd1 vssd1 vccd1 vccd1 _6353_/Q sky130_fd_sc_hd__dfrtp_1
X_6284_ _6441_/CLK _6284_/D vssd1 vssd1 vccd1 vccd1 _6284_/Q sky130_fd_sc_hd__dfxtp_4
X_3496_ _5757_/A _5146_/A _5295_/A _4325_/A vssd1 vssd1 vccd1 vccd1 _3496_/X sky130_fd_sc_hd__a31o_1
X_5304_ _5304_/A _5304_/B _5304_/C _5304_/D vssd1 vssd1 vccd1 vccd1 _5304_/X sky130_fd_sc_hd__or4_2
X_5235_ _5260_/A _4056_/B _5234_/X _3774_/A vssd1 vssd1 vccd1 vccd1 _5235_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_11_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5166_ _5166_/A _5166_/B vssd1 vssd1 vccd1 vccd1 _5166_/Y sky130_fd_sc_hd__nor2_1
X_4117_ _4116_/A _4223_/A _4116_/Y _3759_/Y vssd1 vssd1 vccd1 vccd1 _4117_/X sky130_fd_sc_hd__a211o_1
XANTENNA__4475__S _4482_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5097_ _6408_/Q _5096_/Y _6070_/A vssd1 vssd1 vccd1 vccd1 _5097_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_78_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5245__A2 wire92/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4048_ _6155_/Q _3799_/X _3801_/X _6146_/Q _4047_/X vssd1 vssd1 vccd1 vccd1 _4051_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_91_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4205__A0 _5268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5999_ _3636_/C _3635_/Y hold479/X _3636_/B _5995_/C vssd1 vssd1 vccd1 vccd1 _5999_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_93_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5705__B1 _5721_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4692__A0 _6381_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3495__A1 _5478_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold9 hold9/A vssd1 vssd1 vccd1 vccd1 hold9/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4385__S _4385_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4842__S1 _5078_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5944__S _5977_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold409 _6332_/Q vssd1 vssd1 vccd1 vccd1 hold409/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3350_ _5145_/A _3786_/A vssd1 vssd1 vccd1 vccd1 _4251_/B sky130_fd_sc_hd__nor2_4
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3281_ _3281_/A _5398_/A _5360_/A vssd1 vssd1 vccd1 vccd1 _3281_/X sky130_fd_sc_hd__and3_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5020_ _5019_/X _5018_/X _5101_/S vssd1 vssd1 vccd1 vccd1 _5021_/B sky130_fd_sc_hd__mux2_4
XANTENNA__4683__A0 _6383_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6076__A _6076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4295__S _5232_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5227__A2 _5314_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3212__B _5315_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3789__A2 _3674_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5922_ _5922_/A _5970_/A vssd1 vssd1 vccd1 vccd1 _5924_/A sky130_fd_sc_hd__xnor2_1
X_5853_ _5867_/B _5852_/C _6418_/Q vssd1 vssd1 vccd1 vccd1 _5854_/B sky130_fd_sc_hd__a21oi_1
X_4804_ _5322_/A _5777_/B _4804_/C _4804_/D vssd1 vssd1 vccd1 vccd1 _4806_/C sky130_fd_sc_hd__and4bb_1
XFILLER_0_75_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6015__S _6019_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5935__B1 _5970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5784_ _6023_/A _5976_/S _5977_/S vssd1 vssd1 vccd1 vccd1 _5784_/X sky130_fd_sc_hd__o21a_2
XANTENNA__4202__A3 _6385_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4735_ hold630/X _4734_/X _5232_/S vssd1 vssd1 vccd1 vccd1 _6310_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_8_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4666_ input9/X _4668_/B vssd1 vssd1 vccd1 vccd1 _4666_/X sky130_fd_sc_hd__and2_1
XFILLER_0_43_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3617_ _3617_/A _3617_/B _5619_/A vssd1 vssd1 vccd1 vccd1 _3618_/B sky130_fd_sc_hd__and3_1
X_4597_ _4328_/A _4596_/X _5607_/B2 vssd1 vssd1 vccd1 vccd1 _4597_/X sky130_fd_sc_hd__o21a_1
X_6405_ _6409_/CLK _6405_/D fanout170/X vssd1 vssd1 vccd1 vccd1 _6405_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_0_101_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3548_ _3511_/A _3214_/Y _3547_/X _3213_/X vssd1 vssd1 vccd1 vccd1 _3548_/X sky130_fd_sc_hd__a31o_1
X_6336_ _6336_/CLK _6336_/D fanout183/X vssd1 vssd1 vccd1 vccd1 _6336_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_0_12_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3479_ _3493_/B _3472_/B _3481_/B _6433_/Q vssd1 vssd1 vccd1 vccd1 _3479_/X sky130_fd_sc_hd__a22o_1
X_6267_ _6312_/CLK _6267_/D fanout182/X vssd1 vssd1 vccd1 vccd1 _6267_/Q sky130_fd_sc_hd__dfstp_1
X_5218_ _3632_/C _5217_/X _5218_/S vssd1 vssd1 vccd1 vccd1 _5218_/X sky130_fd_sc_hd__mux2_1
X_6198_ _6263_/CLK _6198_/D vssd1 vssd1 vccd1 vccd1 _6198_/Q sky130_fd_sc_hd__dfxtp_1
X_5149_ _6334_/Q _5243_/S _5244_/S vssd1 vssd1 vccd1 vccd1 _5149_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_98_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3403__A _5617_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5764__S _5765_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3952__A2 _4462_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6486__SET_B fanout172/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5393__B2 _5362_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3943__A2 _3799_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4520_ _4404_/X hold149/X _4527_/S vssd1 vssd1 vccd1 vccd1 _4520_/X sky130_fd_sc_hd__mux2_1
Xhold206 _6252_/Q vssd1 vssd1 vccd1 vccd1 hold206/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold217 _6117_/Q vssd1 vssd1 vccd1 vccd1 hold217/X sky130_fd_sc_hd__dlygate4sd3_1
X_4451_ _4451_/A _4451_/B _4451_/C vssd1 vssd1 vccd1 vccd1 _4452_/B sky130_fd_sc_hd__nor3_1
X_3402_ _5145_/A _3489_/B vssd1 vssd1 vccd1 vccd1 _3619_/C sky130_fd_sc_hd__nand2_4
Xhold239 _6260_/Q vssd1 vssd1 vccd1 vccd1 hold239/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold228 _6232_/Q vssd1 vssd1 vccd1 vccd1 hold228/X sky130_fd_sc_hd__dlygate4sd3_1
X_6121_ _6316_/CLK _6121_/D fanout173/X vssd1 vssd1 vccd1 vccd1 _6121_/Q sky130_fd_sc_hd__dfrtp_1
X_4382_ hold103/X _4085_/X _4385_/S vssd1 vssd1 vccd1 vccd1 _4382_/X sky130_fd_sc_hd__mux2_1
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3333_ _4273_/A _4338_/A _3333_/C vssd1 vssd1 vccd1 vccd1 _3334_/B sky130_fd_sc_hd__or3_2
XFILLER_0_0_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3264_ _3057_/Y _3282_/A _3225_/X _3263_/X vssd1 vssd1 vccd1 vccd1 _3264_/X sky130_fd_sc_hd__o31a_1
XFILLER_0_56_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6052_ _4366_/A _6050_/X _6051_/Y hold493/X _6040_/Y vssd1 vssd1 vccd1 vccd1 _6052_/X
+ sky130_fd_sc_hd__o32a_1
XANTENNA__4319__A _5232_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5003_ _6311_/Q _4963_/B _5002_/B _4796_/Y vssd1 vssd1 vccd1 vccd1 _5003_/X sky130_fd_sc_hd__a22o_1
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3195_ _5605_/A _3304_/B _3311_/B vssd1 vssd1 vccd1 vccd1 _3196_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_56_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout166_A _6159_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4753__S _5232_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5905_ hold391/X _5848_/S _5972_/B1 _5904_/X vssd1 vssd1 vccd1 vccd1 _5905_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4054__A _6334_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5836_ _5867_/B _5835_/C _6417_/Q vssd1 vssd1 vccd1 vccd1 _5837_/B sky130_fd_sc_hd__a21oi_1
X_5767_ _5767_/A _5767_/B vssd1 vssd1 vccd1 vccd1 _5767_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_44_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4187__A2 _3804_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4592__C1 _5600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4718_ _4555_/Y _4717_/Y _5783_/A vssd1 vssd1 vccd1 vccd1 _4719_/A sky130_fd_sc_hd__a21o_2
XFILLER_0_44_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5698_ _6462_/Q _5645_/X _5697_/X _5632_/Y vssd1 vssd1 vccd1 vccd1 _5698_/X sky130_fd_sc_hd__a22o_1
X_4649_ _5567_/B _5418_/B vssd1 vssd1 vccd1 vccd1 _4668_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4895__B1 _6070_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3117__B _4557_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6319_ _6407_/CLK _6319_/D fanout170/X vssd1 vssd1 vccd1 vccd1 _6319_/Q sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_18_wb_clk_i _6448_/CLK vssd1 vssd1 vccd1 vccd1 _6308_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__3133__A _3205_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5759__S _5765_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5072__A0 _6407_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5375__A1 _4675_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5127__A1 _6333_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5678__A2 _4406_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4102__A2 _6290_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_6_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_26_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5602__A2 _3668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3697__B _5478_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3951_ _4438_/A _5302_/B _3942_/Y vssd1 vssd1 vccd1 vccd1 _3951_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_73_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3882_ hold87/A hold65/A _3884_/S vssd1 vssd1 vccd1 vccd1 _3882_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_45_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4305__C _5418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5621_ _4325_/A _4595_/B _3668_/A _5370_/B vssd1 vssd1 vccd1 vccd1 _5624_/C sky130_fd_sc_hd__o211a_1
XFILLER_0_45_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5552_ _5545_/A _5544_/Y _5543_/A vssd1 vssd1 vccd1 vccd1 _5553_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_81_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5417__B _5485_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4503_ _4416_/X hold159/X _4509_/S vssd1 vssd1 vccd1 vccd1 _4503_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5483_ _5483_/A _5483_/B vssd1 vssd1 vccd1 vccd1 _5483_/X sky130_fd_sc_hd__xor2_2
X_4434_ hold203/X hold81/X hold123/X hold151/X _5731_/C1 _4420_/S vssd1 vssd1 vccd1
+ vccd1 _4434_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_1_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4365_ _4919_/S _4364_/X _5769_/S vssd1 vssd1 vccd1 vccd1 _4365_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6529__A _6529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3316_ _3326_/B _3316_/B vssd1 vssd1 vccd1 vccd1 _4267_/B sky130_fd_sc_hd__or2_2
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6104_ hold597/X _6103_/X _6104_/S vssd1 vssd1 vccd1 vccd1 _6489_/D sky130_fd_sc_hd__mux2_1
X_4296_ _4296_/A _4296_/B vssd1 vssd1 vccd1 vccd1 _4296_/X sky130_fd_sc_hd__or2_1
X_6035_ _6036_/A _6036_/B vssd1 vssd1 vccd1 vccd1 _6037_/B sky130_fd_sc_hd__nor2_2
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3247_ _3247_/A _4260_/B vssd1 vssd1 vccd1 vccd1 _3307_/A sky130_fd_sc_hd__or2_2
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3178_ _4268_/A _3247_/A vssd1 vssd1 vccd1 vccd1 _3180_/B sky130_fd_sc_hd__or2_2
XFILLER_0_95_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5579__S _6070_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4801__A0 _5413_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5357__A1 _5600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5819_ _5976_/S _5814_/Y _5818_/X _5786_/Y vssd1 vssd1 vccd1 vccd1 _5819_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5109__A1 _5109_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3128__A _5124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5109__B2 _4924_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4231__B _4463_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold570 _6362_/Q vssd1 vssd1 vccd1 vccd1 hold570/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold581 _6361_/Q vssd1 vssd1 vccd1 vccd1 hold581/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3540__B1 _5384_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold592 _6368_/Q vssd1 vssd1 vccd1 vccd1 hold592/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4885__C _4924_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3843__A1 _3885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5489__S _5489_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5045__A0 _5041_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4393__S _4397_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4406__B _4406_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5596__B2 _5415_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4150_ _4150_/A _6384_/Q vssd1 vssd1 vccd1 vccd1 _4152_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_37_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5284__A0 _6340_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4081_ _4438_/A _6093_/A _4462_/A2 vssd1 vssd1 vccd1 vccd1 _4081_/X sky130_fd_sc_hd__o21a_1
XANTENNA__3204__C _3205_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4983_ _6310_/Q _4963_/B _4982_/B _4796_/Y vssd1 vssd1 vccd1 vccd1 _4983_/X sky130_fd_sc_hd__a22o_1
X_3934_ _6337_/Q _4105_/C vssd1 vssd1 vccd1 vccd1 _4107_/B sky130_fd_sc_hd__nor2_1
XANTENNA__3598__B1 _6529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5339__B2 _5605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3865_ _6172_/Q _6251_/Q _3865_/S vssd1 vssd1 vccd1 vccd1 _3865_/X sky130_fd_sc_hd__mux2_1
X_5604_ _4595_/B _5370_/B _4251_/B _5603_/X vssd1 vssd1 vccd1 vccd1 _5604_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_33_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3796_ _3852_/A _3883_/S _3884_/S vssd1 vssd1 vccd1 vccd1 _4501_/A sky130_fd_sc_hd__or3_1
XANTENNA__5147__B _5291_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5535_ hold391/X _5521_/B _5534_/Y _5417_/Y vssd1 vssd1 vccd1 vccd1 _5535_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_75_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5466_ _5492_/A _5466_/B _5466_/C vssd1 vssd1 vccd1 vccd1 _5468_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_78_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4478__S _4482_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4417_ hold63/X _4416_/X _4464_/S vssd1 vssd1 vccd1 vccd1 hold64/A sky130_fd_sc_hd__mux2_1
X_5397_ _6434_/Q _5600_/C _4354_/A vssd1 vssd1 vccd1 vccd1 _5397_/Y sky130_fd_sc_hd__a21oi_1
X_4348_ _3338_/X _4344_/Y _4346_/X _4347_/X _4333_/X vssd1 vssd1 vccd1 vccd1 _4348_/X
+ sky130_fd_sc_hd__a2111o_1
X_4279_ _3284_/B _4324_/B _5607_/B2 _4278_/X vssd1 vssd1 vccd1 vccd1 _4282_/A sky130_fd_sc_hd__a211o_1
X_6018_ input9/X hold627/X _6019_/S vssd1 vssd1 vccd1 vccd1 _6464_/D sky130_fd_sc_hd__mux2_1
XANTENNA__5610__B _5610_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5578__B2 _5415_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold508_A _6382_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4242__A _4276_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4388__S _5232_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_33_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6407_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_20_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5520__B _5520_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3321__A _5605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6108__S _6108_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5569__A1 _6462_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4152__A _6290_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3650_ _3650_/A _3650_/B _3650_/C vssd1 vssd1 vccd1 vccd1 _3650_/Y sky130_fd_sc_hd__nor3_1
X_3581_ _4338_/A _3581_/B vssd1 vssd1 vccd1 vccd1 _5323_/D sky130_fd_sc_hd__nor2_1
X_5320_ _5600_/A _5313_/X _5314_/X _5315_/Y _5319_/X vssd1 vssd1 vccd1 vccd1 _5320_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_51_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5251_ _5250_/X _5246_/X _5147_/C _3938_/Y vssd1 vssd1 vccd1 vccd1 _5251_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_2_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4202_ _5136_/A _5268_/A _6385_/Q _4060_/B _4201_/X vssd1 vssd1 vccd1 vccd1 _5160_/B
+ sky130_fd_sc_hd__o41a_2
XANTENNA__3913__A_N _6379_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5182_ _5182_/A _5264_/B vssd1 vssd1 vccd1 vccd1 _5186_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__3215__B _3281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4133_ _4190_/A _4052_/B _4053_/B _4053_/A vssd1 vssd1 vccd1 vccd1 _4134_/B sky130_fd_sc_hd__a22oi_2
XANTENNA__6049__A2 _4844_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4064_ _4068_/B _4064_/B vssd1 vssd1 vccd1 vccd1 _4064_/X sky130_fd_sc_hd__and2_1
XFILLER_0_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6018__S _6019_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4966_ _4962_/B _4965_/X _5106_/S vssd1 vssd1 vccd1 vccd1 _4966_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5158__A _5268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3917_ _6285_/Q _3917_/B _3917_/C vssd1 vssd1 vccd1 vccd1 _3918_/B sky130_fd_sc_hd__or3_1
X_4897_ _4896_/X hold371/X _5098_/S vssd1 vssd1 vccd1 vccd1 _4897_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_73_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3848_ _3712_/Y _3715_/Y _3725_/X _3728_/X hold81/A vssd1 vssd1 vccd1 vccd1 _3848_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_46_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3779_ _3979_/A _5162_/A _3763_/X _3778_/X _5294_/A vssd1 vssd1 vccd1 vccd1 _3779_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_61_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5518_ _5518_/A _5518_/B vssd1 vssd1 vccd1 vccd1 _5519_/B sky130_fd_sc_hd__nand2_1
XANTENNA__5605__B _5605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5449_ _6460_/Q _5448_/X _5512_/S vssd1 vssd1 vccd1 vccd1 _5449_/X sky130_fd_sc_hd__mux2_1
Xfanout110 _3183_/A vssd1 vssd1 vccd1 vccd1 _5387_/A sky130_fd_sc_hd__clkbuf_8
Xfanout121 _5478_/S vssd1 vssd1 vccd1 vccd1 _5593_/S sky130_fd_sc_hd__buf_6
XANTENNA__3125__B _3168_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout154 hold647/X vssd1 vssd1 vccd1 vccd1 _4716_/A sky130_fd_sc_hd__buf_4
Xfanout143 _6344_/Q vssd1 vssd1 vccd1 vccd1 _4150_/A sky130_fd_sc_hd__clkbuf_8
Xfanout165 _5600_/A vssd1 vssd1 vccd1 vccd1 _5522_/A sky130_fd_sc_hd__clkbuf_8
Xfanout132 _6430_/Q vssd1 vssd1 vccd1 vccd1 _4276_/A sky130_fd_sc_hd__clkbuf_8
Xfanout176 input18/X vssd1 vssd1 vccd1 vccd1 fanout176/X sky130_fd_sc_hd__buf_4
XANTENNA__3141__A _3497_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3795__B _3885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6308__RESET_B fanout185/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4846__S _4948_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4137__S1 _5721_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4820_ _4819_/X _4919_/S vssd1 vssd1 vccd1 vccd1 _4820_/Y sky130_fd_sc_hd__nand2b_1
X_4751_ _4749_/X _4750_/X _5289_/S vssd1 vssd1 vccd1 vccd1 _4751_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6081__B _6107_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3702_ _6343_/Q _4150_/A vssd1 vssd1 vccd1 vccd1 _3752_/B sky130_fd_sc_hd__nand2_1
X_4682_ _6379_/Q _6285_/Q _4711_/S vssd1 vssd1 vccd1 vccd1 _4682_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_43_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3633_ _3633_/A _4788_/B _3633_/C vssd1 vssd1 vccd1 vccd1 _3634_/B sky130_fd_sc_hd__or3_2
XANTENNA__5714__A1 _4300_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6421_ _6422_/CLK _6421_/D fanout171/X vssd1 vssd1 vccd1 vccd1 _6421_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_31_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3725__B1 _4463_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3564_ _3627_/C _4386_/B _5777_/B _3106_/A vssd1 vssd1 vccd1 vccd1 _3564_/X sky130_fd_sc_hd__o22a_1
X_6352_ _6475_/CLK _6352_/D fanout179/X vssd1 vssd1 vccd1 vccd1 _6352_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3495_ _5478_/S _3594_/A _6468_/Q _3665_/A vssd1 vssd1 vccd1 vccd1 _5499_/S sky130_fd_sc_hd__o31a_4
X_6283_ _6470_/CLK _6283_/D fanout179/X vssd1 vssd1 vccd1 vccd1 _6283_/Q sky130_fd_sc_hd__dfstp_4
X_5303_ _5303_/A _5303_/B _5303_/C _4053_/Y vssd1 vssd1 vccd1 vccd1 _5304_/D sky130_fd_sc_hd__or4b_1
X_5234_ _6345_/Q _3772_/B _4065_/X _5137_/Y _5233_/X vssd1 vssd1 vccd1 vccd1 _5234_/X
+ sky130_fd_sc_hd__a221o_1
X_5165_ _5165_/A _5165_/B vssd1 vssd1 vccd1 vccd1 _5166_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__4756__S _4768_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4116_ _4116_/A _4168_/B vssd1 vssd1 vccd1 vccd1 _4116_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_75_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5441__A _5492_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5096_ _5771_/A _5094_/X _5095_/Y vssd1 vssd1 vccd1 vccd1 _5096_/Y sky130_fd_sc_hd__o21ai_1
X_4047_ _6263_/Q _3793_/X _3795_/X _6198_/Q vssd1 vssd1 vccd1 vccd1 _4047_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4491__S _4491_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5998_ _5995_/C _5995_/B _5988_/X _3473_/X vssd1 vssd1 vccd1 vccd1 _5998_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_93_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4949_ _5064_/A _4949_/B vssd1 vssd1 vccd1 vccd1 _4949_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_74_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3716__B1 _4948_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4141__B1 _3801_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4692__A1 _6287_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3280_ _3639_/C _4325_/C vssd1 vssd1 vccd1 vccd1 _5405_/A sky130_fd_sc_hd__or2_2
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5261__A _6284_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5880__B1 _5867_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6076__B _6107_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5921_ _5977_/S _5920_/X _5784_/X hold586/X vssd1 vssd1 vccd1 vccd1 _5921_/X sky130_fd_sc_hd__o2bb2a_1
XANTENNA__4435__B2 _4441_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5852_ _5852_/A _5867_/B _5852_/C vssd1 vssd1 vccd1 vccd1 _5872_/A sky130_fd_sc_hd__and3_1
XANTENNA__4605__A _5767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4803_ _4803_/A _4803_/B vssd1 vssd1 vccd1 vccd1 _4806_/B sky130_fd_sc_hd__nor2_1
XANTENNA__4324__B _4324_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5783_ _5783_/A _5786_/B vssd1 vssd1 vccd1 vccd1 _5887_/S sky130_fd_sc_hd__or2_2
XANTENNA__5935__A1 _6421_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4734_ _3941_/Y _4733_/X _4770_/S vssd1 vssd1 vccd1 vccd1 _4734_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3946__B1 _3810_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4665_ _3986_/A _4652_/X _4654_/Y _4664_/X vssd1 vssd1 vccd1 vccd1 _6298_/D sky130_fd_sc_hd__o22a_1
X_3616_ _4557_/C _4784_/B _5774_/B _4803_/A vssd1 vssd1 vccd1 vccd1 _5373_/A sky130_fd_sc_hd__a211o_1
X_4596_ _4264_/X _4594_/Y _4595_/X _4593_/X _4276_/A vssd1 vssd1 vccd1 vccd1 _4596_/X
+ sky130_fd_sc_hd__a32o_1
X_6404_ _6407_/CLK _6404_/D fanout170/X vssd1 vssd1 vccd1 vccd1 _6404_/Q sky130_fd_sc_hd__dfrtp_2
X_3547_ _4782_/B _3547_/B _3547_/C vssd1 vssd1 vccd1 vccd1 _3547_/X sky130_fd_sc_hd__and3_1
X_6335_ _6383_/CLK _6335_/D fanout182/X vssd1 vssd1 vccd1 vccd1 _6335_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_0_3_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3478_ hold37/X _3472_/B _3477_/X vssd1 vssd1 vccd1 vccd1 hold38/A sky130_fd_sc_hd__a21o_1
X_6266_ _6488_/CLK _6266_/D vssd1 vssd1 vccd1 vccd1 _6266_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4123__B1 _4462_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5217_ _5291_/S _5215_/Y _5216_/X _5206_/X vssd1 vssd1 vccd1 vccd1 _5217_/X sky130_fd_sc_hd__a2bb2o_1
X_6197_ _6239_/CLK _6197_/D vssd1 vssd1 vccd1 vccd1 _6197_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4486__S _4491_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5148_ _3774_/A _6334_/Q _3773_/Y _5233_/B _5151_/B vssd1 vssd1 vccd1 vccd1 _5148_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA__3403__B _3619_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5079_ _6265_/Q _6200_/Q _6224_/Q _6117_/Q _5100_/S0 _5100_/S1 vssd1 vssd1 vccd1
+ vccd1 _5079_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_19_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4362__B1 _4363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5081__A _5102_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4396__S _4397_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5614__B1 _3489_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5090__A1 _5109_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5090__B2 _4924_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5020__S _5101_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4160__A _6290_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold207 _6261_/Q vssd1 vssd1 vccd1 vccd1 hold207/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4450_ _4451_/B _4451_/C _4451_/A vssd1 vssd1 vccd1 vccd1 _4459_/B sky130_fd_sc_hd__o21a_1
X_3401_ _5145_/A _3489_/B vssd1 vssd1 vccd1 vccd1 _5522_/D sky130_fd_sc_hd__and2_4
XFILLER_0_0_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4381_ hold173/X _4042_/X _4385_/S vssd1 vssd1 vccd1 vccd1 _6145_/D sky130_fd_sc_hd__mux2_1
Xhold218 _6219_/Q vssd1 vssd1 vccd1 vccd1 hold218/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold229 _4526_/X vssd1 vssd1 vccd1 vccd1 _6232_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3332_ _3332_/A _3379_/B vssd1 vssd1 vccd1 vccd1 _5370_/C sky130_fd_sc_hd__nand2_1
X_6120_ _6417_/CLK _6120_/D fanout173/X vssd1 vssd1 vccd1 vccd1 _6120_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3263_ _3326_/A _3547_/C _3268_/B _4273_/B vssd1 vssd1 vccd1 vccd1 _3263_/X sky130_fd_sc_hd__or4_1
X_6051_ _6085_/A _6071_/S vssd1 vssd1 vccd1 vccd1 _6051_/Y sky130_fd_sc_hd__nor2_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3194_ _3323_/A _3205_/B _3229_/A _3168_/B vssd1 vssd1 vccd1 vccd1 _3311_/B sky130_fd_sc_hd__or4bb_2
XANTENNA__3504__A _4325_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5002_ _5102_/A _5002_/B vssd1 vssd1 vccd1 vccd1 _5002_/Y sky130_fd_sc_hd__nand2_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4335__A _5605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5904_ _6403_/Q _6422_/Q _5971_/S vssd1 vssd1 vccd1 vccd1 _5904_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_76_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5908__A1 _5976_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5835_ _6417_/Q _5867_/B _5835_/C vssd1 vssd1 vccd1 vccd1 _5855_/A sky130_fd_sc_hd__and3_1
XFILLER_0_91_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4054__B _6337_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5908__B2 _5786_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5766_ _6316_/Q hold274/X _5766_/S vssd1 vssd1 vccd1 vccd1 _5766_/X sky130_fd_sc_hd__mux2_1
X_4717_ _6023_/A _5243_/S vssd1 vssd1 vccd1 vccd1 _4717_/Y sky130_fd_sc_hd__nand2_1
X_5697_ _4440_/X _5693_/X _4084_/X _5696_/X _5655_/B _5734_/S vssd1 vssd1 vccd1 vccd1
+ _5697_/X sky130_fd_sc_hd__mux4_2
X_4648_ _4653_/A hold365/X hold491/X _3373_/B vssd1 vssd1 vccd1 vccd1 _5418_/B sky130_fd_sc_hd__a211o_1
XFILLER_0_44_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4579_ _4289_/C _4576_/X _4578_/X _6159_/Q vssd1 vssd1 vccd1 vccd1 _5384_/B sky130_fd_sc_hd__a22oi_2
XANTENNA__4895__A1 _6365_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6318_ _6419_/CLK _6318_/D fanout173/X vssd1 vssd1 vccd1 vccd1 _6318_/Q sky130_fd_sc_hd__dfrtp_1
X_6249_ _6449_/CLK hold88/X vssd1 vssd1 vccd1 vccd1 hold87/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__5332__C _6431_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5105__S _5105_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4886__A1 _6365_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6088__B1 _6107_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3324__A _3674_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4638__B2 _6315_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4638__A1 _6464_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold90 hold90/A vssd1 vssd1 vccd1 vccd1 hold90/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3697__C _5344_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3950_ _4045_/A _3950_/B vssd1 vssd1 vccd1 vccd1 _5302_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_73_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6012__A0 _4650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3994__A _6085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3881_ hold55/A hold57/A _3884_/S vssd1 vssd1 vccd1 vccd1 _3881_/X sky130_fd_sc_hd__mux2_1
X_5620_ _3168_/B _3219_/A _4251_/B _5371_/B _5619_/Y vssd1 vssd1 vccd1 vccd1 _5624_/B
+ sky130_fd_sc_hd__a221o_1
X_5551_ _5594_/A _5551_/B vssd1 vssd1 vccd1 vccd1 _5553_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_26_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4502_ _4404_/X hold126/X _4509_/S vssd1 vssd1 vccd1 vccd1 _4502_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3218__B _4268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5482_ _5468_/B _5470_/B _5468_/A vssd1 vssd1 vccd1 vccd1 _5483_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_41_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4433_ hold33/X _3700_/Y _3698_/Y vssd1 vssd1 vccd1 vccd1 _4433_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_67_30 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4364_ _5601_/A _4362_/Y _4366_/B hold346/X vssd1 vssd1 vccd1 vccd1 _4364_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_6_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3315_ _3326_/B _3316_/B vssd1 vssd1 vccd1 vccd1 _3609_/C sky130_fd_sc_hd__nor2_1
X_4295_ _4303_/A _4294_/X _5232_/S vssd1 vssd1 vccd1 vccd1 _4295_/X sky130_fd_sc_hd__mux2_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6103_ _6067_/A _6107_/S _6100_/X _6102_/X vssd1 vssd1 vccd1 vccd1 _6103_/X sky130_fd_sc_hd__a2bb2o_1
X_3246_ _5605_/A _4268_/A vssd1 vssd1 vccd1 vccd1 _4273_/B sky130_fd_sc_hd__nand2_2
X_6034_ _3665_/A _6470_/Q _5418_/A vssd1 vssd1 vccd1 vccd1 _6036_/B sky130_fd_sc_hd__a21oi_2
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3177_ _3326_/A _3547_/C vssd1 vssd1 vccd1 vccd1 _3304_/B sky130_fd_sc_hd__nand2_4
XFILLER_0_83_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4764__S _4770_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5818_ _3094_/Y _5771_/A _4857_/Y _5817_/Y vssd1 vssd1 vccd1 vccd1 _5818_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3368__A1 _5757_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6245__RESET_B fanout180/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5749_ hold9/X _3814_/Y _6104_/S vssd1 vssd1 vccd1 vccd1 hold10/A sky130_fd_sc_hd__mux2_1
XFILLER_0_32_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3128__B _4273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4868__A1 _6364_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold571 _5438_/X vssd1 vssd1 vccd1 vccd1 _6362_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold560 _6426_/Q vssd1 vssd1 vccd1 vccd1 _5951_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold582 _5425_/X vssd1 vssd1 vccd1 vccd1 _6361_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold593 _5513_/X vssd1 vssd1 vccd1 vccd1 _6368_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3144__A _4782_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4406__C _4418_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5596__A2 _5520_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3531__A1 _4325_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3100_ _3100_/A vssd1 vssd1 vccd1 vccd1 _6448_/D sky130_fd_sc_hd__inv_2
XANTENNA__3054__A _5995_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4080_ _6093_/A vssd1 vssd1 vccd1 vccd1 _4080_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_37_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3834__A2 _3799_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3501__B _3501_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3598__A1 _4324_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4982_ _5102_/A _4982_/B vssd1 vssd1 vccd1 vccd1 _4982_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_92_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3933_ _6285_/Q _6286_/Q _6287_/Q vssd1 vssd1 vccd1 vccd1 _3933_/Y sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_3_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6237_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_73_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3864_ _3883_/S _3864_/B vssd1 vssd1 vccd1 vccd1 _3864_/Y sky130_fd_sc_hd__nor2_1
X_5603_ _5603_/A _5603_/B _5603_/C _5603_/D vssd1 vssd1 vccd1 vccd1 _5603_/X sky130_fd_sc_hd__or4_1
XFILLER_0_73_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4011__A2 _6287_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4332__B _4332_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3795_ _3816_/B _3885_/A _3865_/S vssd1 vssd1 vccd1 vccd1 _3795_/X sky130_fd_sc_hd__and3_4
XFILLER_0_26_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5534_ _5534_/A _5534_/B vssd1 vssd1 vccd1 vccd1 _5534_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__4759__S _5232_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5465_ _6479_/Q _4881_/X _5593_/S vssd1 vssd1 vccd1 vccd1 _5466_/C sky130_fd_sc_hd__mux2_1
XFILLER_0_68_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4416_ _4441_/S _4412_/X _4415_/X vssd1 vssd1 vccd1 vccd1 _4416_/X sky130_fd_sc_hd__a21o_2
XFILLER_0_78_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5396_ hold322/X _5645_/A _5513_/S vssd1 vssd1 vccd1 vccd1 _5396_/X sky130_fd_sc_hd__mux2_1
X_4347_ _3284_/B _3229_/C _5388_/A _4338_/X _4345_/X vssd1 vssd1 vccd1 vccd1 _4347_/X
+ sky130_fd_sc_hd__a41o_1
X_4278_ _4270_/X _4272_/X _4275_/X _4277_/X _5600_/A vssd1 vssd1 vccd1 vccd1 _4278_/X
+ sky130_fd_sc_hd__o311a_1
X_3229_ _3229_/A _3547_/B _3229_/C vssd1 vssd1 vccd1 vccd1 _3230_/A sky130_fd_sc_hd__and3_1
XFILLER_0_94_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6017_ input8/X hold620/X _6019_/S vssd1 vssd1 vccd1 vccd1 _6463_/D sky130_fd_sc_hd__mux2_1
XANTENNA__4494__S _4500_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5578__A2 _5520_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3139__A _5124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold390 _3492_/X vssd1 vssd1 vccd1 vccd1 _6438_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5266__A1 _5322_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3602__A _6529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3321__B _4276_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3580_ _5146_/C _3619_/C vssd1 vssd1 vccd1 vccd1 _3643_/B sky130_fd_sc_hd__or2_2
XFILLER_0_3_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5250_ _5290_/S _5249_/X _5147_/C vssd1 vssd1 vccd1 vccd1 _5250_/X sky130_fd_sc_hd__o21a_1
X_4201_ _4060_/B _4195_/X _4196_/Y _4200_/X vssd1 vssd1 vccd1 vccd1 _4201_/X sky130_fd_sc_hd__a31o_1
XANTENNA__6333__SET_B fanout183/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5181_ _5263_/A _5263_/B vssd1 vssd1 vccd1 vccd1 _5187_/A sky130_fd_sc_hd__xor2_1
X_4132_ _4132_/A _4132_/B vssd1 vssd1 vccd1 vccd1 _4134_/A sky130_fd_sc_hd__nor2_1
X_4063_ _6288_/Q _4063_/B _4063_/C vssd1 vssd1 vccd1 vccd1 _4064_/B sky130_fd_sc_hd__or3_1
XANTENNA__3512__A _4276_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3231__B _4268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5009__B2 _4924_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5009__A1 _5109_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4768__A0 hold572/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4965_ _6421_/Q _6369_/Q _5105_/S vssd1 vssd1 vccd1 vccd1 _4965_/X sky130_fd_sc_hd__mux2_1
X_3916_ _5136_/A _3974_/A vssd1 vssd1 vccd1 vccd1 _3916_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_86_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5439__A _5757_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout141_A _4406_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4896_ _6124_/Q _5783_/A _4894_/X _4895_/X vssd1 vssd1 vccd1 vccd1 _4896_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_34_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5717__C1 _3909_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3847_ _4052_/A _3847_/B vssd1 vssd1 vccd1 vccd1 _4437_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_34_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3778_ _4115_/A _5264_/A _3777_/X _3760_/Y _3775_/X vssd1 vssd1 vccd1 vccd1 _3778_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4489__S _4491_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5517_ _5594_/A _5517_/B vssd1 vssd1 vccd1 vccd1 _5518_/B sky130_fd_sc_hd__or2_1
XFILLER_0_100_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5605__C _5605_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5448_ _5446_/X _5447_/X _5499_/S vssd1 vssd1 vccd1 vccd1 _5448_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4918__S1 _6129_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout111 _4199_/A vssd1 vssd1 vccd1 vccd1 _5136_/A sky130_fd_sc_hd__buf_4
Xfanout122 _5410_/A vssd1 vssd1 vccd1 vccd1 _5478_/S sky130_fd_sc_hd__buf_8
X_5379_ _6033_/A _5378_/Y _5769_/S vssd1 vssd1 vccd1 vccd1 _5379_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_10_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout100 _5567_/B vssd1 vssd1 vccd1 vccd1 _6101_/A sky130_fd_sc_hd__buf_4
Xfanout155 _3284_/B vssd1 vssd1 vccd1 vccd1 _3229_/A sky130_fd_sc_hd__buf_4
Xfanout144 _4273_/A vssd1 vssd1 vccd1 vccd1 _3986_/A sky130_fd_sc_hd__clkbuf_8
Xfanout133 _5777_/A vssd1 vssd1 vccd1 vccd1 _3786_/A sky130_fd_sc_hd__buf_4
XANTENNA__5248__A1 _6383_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout166 _6159_/Q vssd1 vssd1 vccd1 vccd1 _5600_/A sky130_fd_sc_hd__clkbuf_8
Xfanout177 fanout180/X vssd1 vssd1 vccd1 vccd1 fanout177/X sky130_fd_sc_hd__clkbuf_8
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold618_A _6459_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5420__B2 _5567_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5708__C1 _5721_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3498__B1 _5567_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6348__RESET_B fanout185/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4462__A2 _4462_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4750_ hold359/X _4312_/B _4768_/S vssd1 vssd1 vccd1 vccd1 _4750_/X sky130_fd_sc_hd__mux2_1
X_4681_ _6081_/A _4714_/S vssd1 vssd1 vccd1 vccd1 _4681_/Y sky130_fd_sc_hd__nor2_1
X_3701_ _4418_/C _3701_/B vssd1 vssd1 vccd1 vccd1 _3717_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_16_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3632_ _4276_/A _6159_/Q _3632_/C _3632_/D vssd1 vssd1 vccd1 vccd1 _3633_/C sky130_fd_sc_hd__and4_1
X_6420_ _6422_/CLK _6420_/D fanout170/X vssd1 vssd1 vccd1 vccd1 _6420_/Q sky130_fd_sc_hd__dfrtp_4
X_6351_ _6377_/CLK _6351_/D fanout179/X vssd1 vssd1 vccd1 vccd1 _6351_/Q sky130_fd_sc_hd__dfrtp_1
X_3563_ _6431_/Q _3396_/B _4253_/A _5146_/D vssd1 vssd1 vccd1 vccd1 _3563_/X sky130_fd_sc_hd__o2bb2a_1
X_5302_ _5302_/A _5302_/B _5302_/C _5302_/D vssd1 vssd1 vccd1 vccd1 _5303_/C sky130_fd_sc_hd__or4_1
X_3494_ _3487_/B hold305/X _3493_/X _3472_/B vssd1 vssd1 vccd1 vccd1 _6439_/D sky130_fd_sc_hd__a22o_1
X_6282_ _6383_/CLK _6282_/D fanout182/X vssd1 vssd1 vccd1 vccd1 _6282_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA__5478__A1 _4901_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5233_ _4065_/X _5233_/B vssd1 vssd1 vccd1 vccd1 _5233_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_11_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5164_ _5164_/A _5164_/B vssd1 vssd1 vccd1 vccd1 _5165_/B sky130_fd_sc_hd__xnor2_1
X_4115_ _4115_/A _5262_/D vssd1 vssd1 vccd1 vccd1 _4115_/X sky130_fd_sc_hd__and2_1
X_5095_ _6464_/Q _5771_/A vssd1 vssd1 vccd1 vccd1 _5095_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__4989__B1 _5108_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4046_ _3902_/Y _4045_/X _4044_/X vssd1 vssd1 vccd1 vccd1 _4053_/A sky130_fd_sc_hd__o21bai_2
XFILLER_0_91_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5650__A1 _6458_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5997_ _3635_/Y _5996_/Y _4363_/A _3471_/B vssd1 vssd1 vccd1 vccd1 _6434_/D sky130_fd_sc_hd__o2bb2a_1
XANTENNA__5402__A1 _4595_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4948_ _4942_/B _4947_/X _4948_/S vssd1 vssd1 vccd1 vccd1 _4948_/X sky130_fd_sc_hd__mux2_1
X_4879_ hold85/A _6190_/Q _6174_/Q _6253_/Q _5100_/S0 _5100_/S1 vssd1 vssd1 vccd1
+ vccd1 _4879_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_34_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5705__A2 _5721_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5108__S _5108_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4947__S _5105_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold470_A _6287_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold568_A _6422_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4248__A _6430_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6441__RESET_B fanout185/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4682__S _4711_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5641__A1 _5734_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4904__A0 _4901_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5880__A1 _5866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3062__A _6159_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5920_ _5014_/Y _5786_/Y _5919_/X _5915_/X _5976_/S vssd1 vssd1 vccd1 vccd1 _5920_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_88_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5851_ _5866_/A _6463_/Q _5866_/C vssd1 vssd1 vccd1 vccd1 _5852_/C sky130_fd_sc_hd__or3_1
XANTENNA__4605__B _4605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5782_ _5778_/Y _5867_/B _5781_/X _5418_/A vssd1 vssd1 vccd1 vccd1 _5786_/B sky130_fd_sc_hd__o31a_1
X_4802_ _4802_/A _4802_/B _4802_/C _4802_/D vssd1 vssd1 vccd1 vccd1 _4924_/C sky130_fd_sc_hd__and4_4
XANTENNA__5935__A2 _6422_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4733_ _4731_/X _4732_/X _5289_/S vssd1 vssd1 vccd1 vccd1 _4733_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3936__S _6285_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4664_ input8/X _4668_/B vssd1 vssd1 vccd1 vccd1 _4664_/X sky130_fd_sc_hd__and2_1
XFILLER_0_43_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6403_ _6409_/CLK _6403_/D fanout170/X vssd1 vssd1 vccd1 vccd1 _6403_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__5699__A1 _6313_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3615_ _4784_/C _5307_/C _5310_/D _3615_/D vssd1 vssd1 vccd1 vccd1 _4803_/A sky130_fd_sc_hd__or4_1
XANTENNA__3237__A _4273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4595_ _6432_/Q _4595_/B vssd1 vssd1 vccd1 vccd1 _4595_/X sky130_fd_sc_hd__or2_1
X_3546_ _6432_/Q _3785_/B _3481_/B _3472_/B hold35/X vssd1 vssd1 vccd1 vccd1 hold36/A
+ sky130_fd_sc_hd__a32o_1
X_6334_ _6340_/CLK _6334_/D fanout183/X vssd1 vssd1 vccd1 vccd1 _6334_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA_fanout104_A _3390_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6265_ _6265_/CLK _6265_/D vssd1 vssd1 vccd1 vccd1 _6265_/Q sky130_fd_sc_hd__dfxtp_1
X_3477_ _3477_/A _3785_/B _5387_/C _3481_/B vssd1 vssd1 vccd1 vccd1 _3477_/X sky130_fd_sc_hd__and4_1
X_5216_ _5151_/B _5157_/X _5291_/S vssd1 vssd1 vccd1 vccd1 _5216_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_50_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6196_ _6376_/CLK _6196_/D vssd1 vssd1 vccd1 vccd1 _6196_/Q sky130_fd_sc_hd__dfxtp_1
X_5147_ _5292_/S _5291_/S _5147_/C vssd1 vssd1 vccd1 vccd1 _5147_/X sky130_fd_sc_hd__and3_1
XFILLER_0_79_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5078_ _6157_/Q _6148_/Q _6140_/Q _6184_/Q _5404_/A0 _5078_/S1 vssd1 vssd1 vccd1
+ vccd1 _5078_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_79_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5623__B2 _5777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4029_ _6089_/A vssd1 vssd1 vccd1 vccd1 _4029_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_39_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5139__B1 _6333_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5627__A _5734_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3147__A _5369_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4362__A1 _4948_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4677__S _4711_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4114__A1 _6290_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5362__A _5362_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4665__A2 _4652_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5081__B _6101_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4706__A _6067_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5378__B1 _6021_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4050__B1 _3810_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold208 _6264_/Q vssd1 vssd1 vccd1 vccd1 hold208/X sky130_fd_sc_hd__dlygate4sd3_1
X_3400_ _3308_/B _3399_/X _4325_/A vssd1 vssd1 vccd1 vccd1 _3400_/X sky130_fd_sc_hd__o21a_1
XANTENNA__4353__B2 _3284_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4380_ hold95/X _3998_/X _4385_/S vssd1 vssd1 vccd1 vccd1 hold96/A sky130_fd_sc_hd__mux2_1
Xhold219 _4512_/X vssd1 vssd1 vccd1 vccd1 _6219_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3331_ _4273_/A _5374_/B vssd1 vssd1 vccd1 vccd1 _3379_/B sky130_fd_sc_hd__nand2_1
XANTENNA__6363__RESET_B fanout175/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3262_ _3196_/B _3205_/X _4357_/C vssd1 vssd1 vccd1 vccd1 _3272_/B sky130_fd_sc_hd__o21ai_1
X_6050_ _5567_/B _6049_/X _6071_/S vssd1 vssd1 vccd1 vccd1 _6050_/X sky130_fd_sc_hd__o21a_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3193_ _3316_/B _3228_/C vssd1 vssd1 vccd1 vccd1 _3193_/X sky130_fd_sc_hd__and2_1
XANTENNA__3504__B _6019_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5001_ _5000_/X _4999_/X _5101_/S vssd1 vssd1 vccd1 vccd1 _5002_/B sky130_fd_sc_hd__mux2_2
XANTENNA__5853__A1 _5867_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4319__C _5783_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5903_ _5912_/B _5903_/B vssd1 vssd1 vccd1 vccd1 _5903_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_72_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5834_ _5866_/A _6462_/Q _5866_/C vssd1 vssd1 vccd1 vccd1 _5835_/C sky130_fd_sc_hd__or3_1
XFILLER_0_91_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5765_ _6316_/Q hold572/X _5765_/S vssd1 vssd1 vccd1 vccd1 _5765_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_29_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3395__A2 _5314_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4716_ _4716_/A _5124_/A _6159_/Q _5369_/B vssd1 vssd1 vccd1 vccd1 _5243_/S sky130_fd_sc_hd__and4_2
XFILLER_0_44_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5696_ _5696_/A _5696_/B vssd1 vssd1 vccd1 vccd1 _5696_/X sky130_fd_sc_hd__or2_1
X_4647_ hold298/X _4646_/X _3373_/B vssd1 vssd1 vccd1 vccd1 _4647_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_4_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4578_ _4276_/A _4595_/B _4267_/Y _4577_/X vssd1 vssd1 vccd1 vccd1 _4578_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_12_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4497__S _4500_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6317_ _6419_/CLK _6317_/D fanout173/X vssd1 vssd1 vccd1 vccd1 _6317_/Q sky130_fd_sc_hd__dfrtp_1
X_3529_ _4332_/B _4784_/D _3305_/B _5346_/A vssd1 vssd1 vccd1 vccd1 _3530_/B sky130_fd_sc_hd__a211o_1
X_6248_ _6248_/CLK _6248_/D fanout180/X vssd1 vssd1 vccd1 vccd1 _6248_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__4647__A2 _4646_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6179_ _6489_/CLK _6179_/D vssd1 vssd1 vccd1 vccd1 _6179_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5844__A1 _6365_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5910__A _6423_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6163__D _6163_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_27_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6384_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__4032__B1 _3801_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4583__A1 _5605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5780__B1 _5995_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold80 hold80/A vssd1 vssd1 vccd1 vccd1 hold80/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold91 hold91/A vssd1 vssd1 vccd1 vccd1 hold91/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6448__CLK _6448_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3880_ _3878_/X _3880_/B vssd1 vssd1 vccd1 vccd1 _5299_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_42_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4574__A1 _6339_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5550_ _6486_/Q _5021_/B _5593_/S vssd1 vssd1 vccd1 vccd1 _5551_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_26_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4501_ _4501_/A _6003_/B vssd1 vssd1 vccd1 vccd1 _4509_/S sky130_fd_sc_hd__or2_4
X_5481_ _5481_/A _5481_/B vssd1 vssd1 vccd1 vccd1 _5483_/A sky130_fd_sc_hd__nor2_1
XANTENNA__4326__A1 _3673_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4432_ _4414_/A _5300_/D _4030_/Y vssd1 vssd1 vccd1 vccd1 _4432_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_0_41_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4877__A2 _5783_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4363_ _4363_/A _4363_/B vssd1 vssd1 vccd1 vccd1 _4366_/B sky130_fd_sc_hd__or2_1
XFILLER_0_1_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6079__A1 _6101_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4110__S _6334_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3314_ _4784_/B _3314_/B vssd1 vssd1 vccd1 vccd1 _5346_/B sky130_fd_sc_hd__or2_1
XFILLER_0_67_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4294_ _4296_/B _4293_/Y _6309_/Q _4322_/B vssd1 vssd1 vccd1 vccd1 _4294_/X sky130_fd_sc_hd__a2bb2o_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6102_ hold597/X _6070_/A _6107_/S _6101_/X vssd1 vssd1 vccd1 vccd1 _6102_/X sky130_fd_sc_hd__o211a_1
XANTENNA__6079__B2 _6036_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3245_ _5315_/A _3183_/X _3333_/C _5398_/A vssd1 vssd1 vccd1 vccd1 _3253_/A sky130_fd_sc_hd__o22a_1
X_6033_ _6033_/A _6033_/B _6073_/B _4670_/C vssd1 vssd1 vccd1 vccd1 _6071_/S sky130_fd_sc_hd__or4b_4
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3837__B1 _3810_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3176_ _3229_/A _3229_/C vssd1 vssd1 vccd1 vccd1 _3176_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__3250__A _5315_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout171_A fanout172/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5817_ _5817_/A _5817_/B vssd1 vssd1 vccd1 vccd1 _5817_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__5762__A0 _6313_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4565__A1 _6314_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5748_ hold13/X _4641_/A _6104_/S vssd1 vssd1 vccd1 vccd1 hold14/A sky130_fd_sc_hd__mux2_1
XFILLER_0_17_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5679_ _6173_/Q _4406_/B _4420_/S _6252_/Q _5731_/C1 vssd1 vssd1 vccd1 vccd1 _5680_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_32_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold550 _6438_/Q vssd1 vssd1 vccd1 vccd1 _5988_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xhold561 _5956_/X vssd1 vssd1 vccd1 vccd1 _6426_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold572 _6409_/Q vssd1 vssd1 vccd1 vccd1 hold572/X sky130_fd_sc_hd__clkbuf_2
Xhold583 _6363_/Q vssd1 vssd1 vccd1 vccd1 hold583/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold594 _6490_/Q vssd1 vssd1 vccd1 vccd1 hold594/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3144__B _3172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout84_A _4408_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold648_A _6297_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5348__A3 _3304_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3319__B _5314_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4308__A1 _5581_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4403__S1 _5731_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4859__A2 _4957_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4748__A1_N _6313_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3070__A _4366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4981_ _4980_/X _4979_/X _5101_/S vssd1 vssd1 vccd1 vccd1 _4982_/B sky130_fd_sc_hd__mux2_2
X_3932_ _6285_/Q _6286_/Q _6287_/Q vssd1 vssd1 vccd1 vccd1 _4105_/C sky130_fd_sc_hd__o21a_1
XFILLER_0_73_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3863_ hold69/A _6188_/Q _3865_/S vssd1 vssd1 vccd1 vccd1 _3864_/B sky130_fd_sc_hd__mux2_1
X_5602_ _5346_/A _3668_/A _5362_/A _4595_/B _5362_/D vssd1 vssd1 vccd1 vccd1 _5603_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_73_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4011__A3 _6381_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5533_ _5519_/A _5519_/B _5518_/A vssd1 vssd1 vccd1 vccd1 _5534_/B sky130_fd_sc_hd__o21a_1
X_3794_ _3852_/A _3883_/S _3865_/S vssd1 vssd1 vccd1 vccd1 _4546_/B sky130_fd_sc_hd__or3_1
XFILLER_0_26_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5464_ _5757_/A _6462_/Q vssd1 vssd1 vccd1 vccd1 _5466_/B sky130_fd_sc_hd__or2_1
XFILLER_0_78_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5395_ _4406_/B _5394_/X _5769_/S vssd1 vssd1 vccd1 vccd1 _6355_/D sky130_fd_sc_hd__mux2_1
X_4415_ _6387_/Q _4462_/A2 _3942_/Y _4414_/Y _3698_/Y vssd1 vssd1 vccd1 vccd1 _4415_/X
+ sky130_fd_sc_hd__o221a_1
X_4346_ _5346_/A _3668_/A _5388_/B _3284_/B _4249_/B vssd1 vssd1 vccd1 vccd1 _4346_/X
+ sky130_fd_sc_hd__a221o_1
X_4277_ _4273_/X _4276_/X _4325_/C vssd1 vssd1 vccd1 vccd1 _4277_/X sky130_fd_sc_hd__a21o_1
X_3228_ _3627_/B _3316_/B _3228_/C vssd1 vssd1 vccd1 vccd1 _3228_/X sky130_fd_sc_hd__and3_1
X_6016_ input6/X hold621/X _6019_/S vssd1 vssd1 vccd1 vccd1 _6462_/D sky130_fd_sc_hd__mux2_1
X_3159_ _4360_/B _3527_/B vssd1 vssd1 vccd1 vccd1 _5345_/B sky130_fd_sc_hd__or2_1
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3139__B _5315_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold598_A _6338_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4710__A1 _4715_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold380 _5846_/X vssd1 vssd1 vccd1 vccd1 _6417_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold391 _6370_/Q vssd1 vssd1 vccd1 vccd1 hold391/X sky130_fd_sc_hd__buf_1
XANTENNA__3321__C _4595_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_42_wb_clk_i clkbuf_leaf_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6489_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_87_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4226__A0 _6465_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5974__A0 _6465_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4200_ _3753_/X _4197_/X _4199_/B _4199_/Y _5136_/B vssd1 vssd1 vccd1 vccd1 _4200_/X
+ sky130_fd_sc_hd__a32o_1
X_5180_ _5180_/A _5180_/B vssd1 vssd1 vccd1 vccd1 _5180_/Y sky130_fd_sc_hd__xnor2_1
X_4131_ _4190_/A _4131_/B vssd1 vssd1 vccd1 vccd1 _4132_/B sky130_fd_sc_hd__nor2_1
X_4062_ _4063_/B _4063_/C _6288_/Q vssd1 vssd1 vccd1 vccd1 _4068_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5965__B1 _5771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4964_ _6483_/Q _5104_/A2 _4796_/Y _4962_/B _4963_/X vssd1 vssd1 vccd1 vccd1 _4964_/X
+ sky130_fd_sc_hd__a221o_1
X_3915_ _3917_/B _3917_/C _6285_/Q vssd1 vssd1 vccd1 vccd1 _3974_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_80_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5439__B _6460_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4895_ _6365_/Q _5863_/S _6070_/A vssd1 vssd1 vccd1 vccd1 _4895_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_73_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout134_A _4313_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3846_ _3846_/A _3846_/B _3846_/C vssd1 vssd1 vccd1 vccd1 _3847_/B sky130_fd_sc_hd__or3_4
XFILLER_0_89_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3777_ _6378_/Q _4223_/A _3759_/Y vssd1 vssd1 vccd1 vccd1 _3777_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_80_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3728__C1 _4948_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5516_ _5594_/A _5517_/B vssd1 vssd1 vccd1 vccd1 _5518_/A sky130_fd_sc_hd__nand2_1
XANTENNA__4940__A1 _5101_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5447_ hold583/X _4658_/A _5510_/S vssd1 vssd1 vccd1 vccd1 _5447_/X sky130_fd_sc_hd__mux2_1
Xfanout101 _5499_/S vssd1 vssd1 vccd1 vccd1 _5567_/B sky130_fd_sc_hd__buf_6
X_5378_ _4641_/B _5377_/Y _6021_/S vssd1 vssd1 vccd1 vccd1 _5378_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_10_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout112 _6108_/S vssd1 vssd1 vccd1 vccd1 _6104_/S sky130_fd_sc_hd__buf_6
Xfanout156 _3284_/B vssd1 vssd1 vccd1 vccd1 _4782_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__3125__D _3205_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout145 _5605_/C vssd1 vssd1 vccd1 vccd1 _4273_/A sky130_fd_sc_hd__buf_4
Xfanout134 _4313_/A vssd1 vssd1 vccd1 vccd1 _5777_/A sky130_fd_sc_hd__buf_4
X_4329_ _3278_/A _3668_/A _4327_/X _5605_/B _4328_/X vssd1 vssd1 vccd1 vccd1 _4329_/X
+ sky130_fd_sc_hd__a221o_1
Xfanout123 _5384_/A vssd1 vssd1 vccd1 vccd1 _4366_/A sky130_fd_sc_hd__clkbuf_8
XANTENNA__5248__A2 _5314_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout178 fanout180/X vssd1 vssd1 vccd1 vccd1 fanout178/X sky130_fd_sc_hd__buf_4
Xfanout167 _5078_/S1 vssd1 vssd1 vccd1 vccd1 _5100_/S1 sky130_fd_sc_hd__clkbuf_8
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5708__B1 _5721_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3498__A1 _4363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3700_ _3700_/A _3700_/B vssd1 vssd1 vccd1 vccd1 _3700_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__5974__S _5974_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4680_ _4715_/B2 _4673_/Y _4679_/X hold310/X _4672_/Y vssd1 vssd1 vccd1 vccd1 _4680_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_0_16_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3631_ _4335_/B hold59/X hold328/X _6433_/Q _3630_/X vssd1 vssd1 vccd1 vccd1 _4788_/B
+ sky130_fd_sc_hd__a221o_2
X_3562_ _3786_/A _3619_/C vssd1 vssd1 vccd1 vccd1 _5146_/D sky130_fd_sc_hd__or2_4
XANTENNA__3725__A2 _3701_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6350_ _6377_/CLK _6350_/D fanout176/X vssd1 vssd1 vccd1 vccd1 _6350_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5275__A _6407_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5301_ _5301_/A _5301_/B _5301_/C _5300_/X vssd1 vssd1 vccd1 vccd1 _5302_/D sky130_fd_sc_hd__or4b_1
X_3493_ _3493_/A _3493_/B _3493_/C hold35/X vssd1 vssd1 vccd1 vccd1 _3493_/X sky130_fd_sc_hd__or4_1
X_6281_ _6383_/CLK _6281_/D fanout182/X vssd1 vssd1 vccd1 vccd1 _6281_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_0_11_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4686__A0 _6380_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5232_ hold603/X _5231_/X _5232_/S vssd1 vssd1 vccd1 vccd1 _6336_/D sky130_fd_sc_hd__mux2_1
X_5163_ _5163_/A _5256_/B vssd1 vssd1 vccd1 vccd1 _5164_/B sky130_fd_sc_hd__xnor2_1
X_4114_ _6288_/Q _6290_/Q _4716_/A vssd1 vssd1 vccd1 vccd1 _5262_/D sky130_fd_sc_hd__mux2_1
XANTENNA__3523__A _5322_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5094_ _5102_/A _5093_/Y _5081_/Y vssd1 vssd1 vccd1 vccd1 _5094_/X sky130_fd_sc_hd__o21a_1
XANTENNA__5635__C1 _5731_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4045_ _4045_/A _4045_/B _4038_/A vssd1 vssd1 vccd1 vccd1 _4045_/X sky130_fd_sc_hd__or3b_1
XANTENNA__3661__A1 _6283_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5996_ _3480_/B _5978_/Y _5995_/X vssd1 vssd1 vccd1 vccd1 _5996_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_19_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4947_ _6420_/Q _6368_/Q _5105_/S vssd1 vssd1 vccd1 vccd1 _4947_/X sky130_fd_sc_hd__mux2_1
X_4878_ _4877_/X hold355/X _5098_/S vssd1 vssd1 vccd1 vccd1 _4878_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6475__SET_B fanout175/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3829_ _6232_/Q _3731_/X _3804_/X _6455_/Q vssd1 vssd1 vccd1 vccd1 _3830_/C sky130_fd_sc_hd__a22o_1
XFILLER_0_42_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6479_ _6481_/CLK _6479_/D fanout176/X vssd1 vssd1 vccd1 vccd1 _6479_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA__4677__A0 _6378_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4141__A2 _3799_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3152__B _5605_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5154__A2_N _5292_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold630_A _6310_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4264__A _4675_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5095__A _6464_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5880__A2 _6465_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5850_ _6366_/Q _5849_/X _5974_/S vssd1 vssd1 vccd1 vccd1 _5850_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_68_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5781_ _4289_/C _4264_/B _5317_/B _5780_/X _6434_/Q vssd1 vssd1 vccd1 vccd1 _5781_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_0_61_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4801_ _5413_/B _4800_/X _4948_/S vssd1 vssd1 vccd1 vccd1 _4801_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5935__A3 _6423_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5396__A1 _5645_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4732_ hold456/X _4296_/A _4768_/S vssd1 vssd1 vccd1 vccd1 _4732_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_8_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3946__A2 _3731_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4663_ _3511_/A _4652_/X _4654_/Y _4662_/X vssd1 vssd1 vccd1 vccd1 _6297_/D sky130_fd_sc_hd__o22a_1
XFILLER_0_83_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3614_ _3614_/A _4260_/B vssd1 vssd1 vccd1 vccd1 _3615_/D sky130_fd_sc_hd__nor2_1
X_6402_ _6422_/CLK _6402_/D fanout170/X vssd1 vssd1 vccd1 vccd1 _6402_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4594_ _6432_/Q _4595_/B vssd1 vssd1 vccd1 vccd1 _4594_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_24_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6333_ _6340_/CLK _6333_/D fanout183/X vssd1 vssd1 vccd1 vccd1 _6333_/Q sky130_fd_sc_hd__dfstp_4
X_3545_ hold39/X _3472_/B _3492_/C vssd1 vssd1 vccd1 vccd1 hold40/A sky130_fd_sc_hd__a21o_1
XFILLER_0_10_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3476_ _3487_/B _3488_/A vssd1 vssd1 vccd1 vccd1 _3481_/B sky130_fd_sc_hd__and2_1
X_6264_ _6265_/CLK _6264_/D vssd1 vssd1 vccd1 vccd1 _6264_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5320__A1 _5600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5215_ _5215_/A _5215_/B vssd1 vssd1 vccd1 vccd1 _5215_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__4123__A2 _6097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6195_ _6490_/CLK _6195_/D vssd1 vssd1 vccd1 vccd1 _6195_/Q sky130_fd_sc_hd__dfxtp_1
X_5146_ _5146_/A _5146_/B _5146_/C _5146_/D vssd1 vssd1 vccd1 vccd1 _5147_/C sky130_fd_sc_hd__or4_4
XANTENNA__5879__S _6021_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5077_ _5076_/X hold427/X _5098_/S vssd1 vssd1 vccd1 vccd1 _5077_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5629__A_N _5644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4028_ _4227_/S _4026_/X _4027_/X vssd1 vssd1 vccd1 vccd1 _6089_/A sky130_fd_sc_hd__a21oi_4
XFILLER_0_79_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5979_ _6437_/Q _5988_/B vssd1 vssd1 vccd1 vccd1 _5979_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_47_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3428__A _4313_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3862__S _3883_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4693__S _4712_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5075__A0 _6463_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5614__A2 _4595_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4706__B _4714_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5378__A1 _4641_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4586__C1 _5388_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5029__S _5108_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold209 _6341_/Q vssd1 vssd1 vccd1 vccd1 _3632_/C sky130_fd_sc_hd__buf_1
XANTENNA__5550__A1 _5021_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4868__S _5105_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3330_ _3229_/A _4338_/A _3547_/C _3376_/B vssd1 vssd1 vccd1 vccd1 _3334_/C sky130_fd_sc_hd__a31o_1
XFILLER_0_21_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3261_ _3581_/B _3261_/B _3261_/C vssd1 vssd1 vccd1 vccd1 _5327_/B sky130_fd_sc_hd__and3_1
X_5000_ _6261_/Q _6196_/Q _6220_/Q _6113_/Q _5404_/A0 _5078_/S1 vssd1 vssd1 vccd1
+ vccd1 _5000_/X sky130_fd_sc_hd__mux4_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3192_ _3547_/C _3232_/C vssd1 vssd1 vccd1 vccd1 _3228_/C sky130_fd_sc_hd__nand2_1
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5066__A0 _6426_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3616__A1 _4557_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5902_ _6421_/Q _5970_/A _5912_/A vssd1 vssd1 vccd1 vccd1 _5903_/B sky130_fd_sc_hd__a21oi_1
X_5833_ _5977_/S _5832_/X _5784_/X hold375/X vssd1 vssd1 vccd1 vccd1 _5833_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_63_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5764_ _6315_/Q hold512/X _5765_/S vssd1 vssd1 vccd1 vccd1 _5764_/X sky130_fd_sc_hd__mux2_1
X_4715_ hold330/X _4672_/Y _4714_/X _4715_/B2 vssd1 vssd1 vccd1 vccd1 _4715_/X sky130_fd_sc_hd__o22a_1
X_5695_ _6138_/Q _5721_/A2 _4235_/S _6182_/Q _5721_/C1 vssd1 vssd1 vccd1 vccd1 _5696_/B
+ sky130_fd_sc_hd__o221a_1
X_4646_ _6445_/D _6445_/Q vssd1 vssd1 vccd1 vccd1 _4646_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_44_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4577_ _5774_/A _4595_/B _5317_/B vssd1 vssd1 vccd1 vccd1 _4577_/X sky130_fd_sc_hd__and3_1
XFILLER_0_71_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6316_ _6316_/CLK _6316_/D fanout174/X vssd1 vssd1 vccd1 vccd1 _6316_/Q sky130_fd_sc_hd__dfstp_2
X_3528_ hold347/X _5400_/B _3527_/X _5398_/A vssd1 vssd1 vccd1 vccd1 _3528_/X sky130_fd_sc_hd__a22o_1
X_6247_ _6248_/CLK hold48/X fanout180/X vssd1 vssd1 vccd1 vccd1 hold47/A sky130_fd_sc_hd__dfrtp_1
X_3459_ _5522_/A _3437_/Y _3456_/X _3458_/X _5995_/C vssd1 vssd1 vccd1 vccd1 _3464_/D
+ sky130_fd_sc_hd__a311oi_2
X_6178_ _6399_/CLK _6178_/D vssd1 vssd1 vccd1 vccd1 _6178_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5129_ _6021_/S _5783_/A vssd1 vssd1 vccd1 vccd1 _5132_/B sky130_fd_sc_hd__nor2_1
XANTENNA__5910__B _5970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4280__A1 _4276_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4280__B2 _5398_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4583__A2 _5605_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5780__A1 _4324_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4717__A _6023_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold81 hold81/A vssd1 vssd1 vccd1 vccd1 hold81/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5048__B1 _5108_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold92 hold92/A vssd1 vssd1 vccd1 vccd1 hold92/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold70 hold70/A vssd1 vssd1 vccd1 vccd1 hold70/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4500_ _4463_/X hold255/X _4500_/S vssd1 vssd1 vccd1 vccd1 _4500_/X sky130_fd_sc_hd__mux2_1
X_5480_ _5492_/A _5479_/B _5479_/C vssd1 vssd1 vccd1 vccd1 _5481_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_101_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_1 _3364_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4431_ _4431_/A _4431_/B vssd1 vssd1 vccd1 vccd1 _5300_/D sky130_fd_sc_hd__xnor2_1
X_4362_ _4948_/S _4363_/B _4363_/A vssd1 vssd1 vccd1 vccd1 _4362_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3313_ _3326_/B _4260_/B _3414_/B _3614_/A vssd1 vssd1 vccd1 vccd1 _5406_/B sky130_fd_sc_hd__o22a_1
XFILLER_0_67_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4293_ _4303_/A _3506_/B _4310_/S vssd1 vssd1 vccd1 vccd1 _4293_/Y sky130_fd_sc_hd__o21ai_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6101_ _6101_/A _6101_/B _6101_/C vssd1 vssd1 vccd1 vccd1 _6101_/X sky130_fd_sc_hd__or3_1
XANTENNA__6079__A2 _4982_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3244_ _5387_/A _3304_/B vssd1 vssd1 vccd1 vccd1 _3333_/C sky130_fd_sc_hd__or2_1
X_6032_ _6032_/A _6032_/B _6032_/C vssd1 vssd1 vccd1 vccd1 _6073_/B sky130_fd_sc_hd__or3_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3175_ _3240_/B _3174_/X _3106_/A vssd1 vssd1 vccd1 vccd1 _3186_/C sky130_fd_sc_hd__a21oi_1
XFILLER_0_76_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout164_A _5600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5816_ _5815_/X _6363_/Q _5816_/S vssd1 vssd1 vccd1 vccd1 _5817_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_17_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5747_ hold31/X _4636_/A _6104_/S vssd1 vssd1 vccd1 vccd1 hold32/A sky130_fd_sc_hd__mux2_1
XFILLER_0_32_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5678_ _6452_/Q _4406_/B _4420_/S _6229_/Q _3909_/Y vssd1 vssd1 vccd1 vccd1 _5680_/A
+ sky130_fd_sc_hd__o221a_1
X_4629_ _4602_/Y _4626_/X _4628_/X vssd1 vssd1 vccd1 vccd1 _4629_/X sky130_fd_sc_hd__a21o_1
Xhold551 _5979_/Y vssd1 vssd1 vccd1 vccd1 hold551/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold562 _6374_/Q vssd1 vssd1 vccd1 vccd1 hold562/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold540 _5599_/X vssd1 vssd1 vccd1 vccd1 _6376_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4301__S _4310_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold595 _6365_/Q vssd1 vssd1 vccd1 vccd1 hold595/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold584 _5450_/X vssd1 vssd1 vccd1 vccd1 _6363_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_49_wb_clk_i_A clkbuf_leaf_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold573 _5765_/X vssd1 vssd1 vccd1 vccd1 _6409_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3144__C _3284_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3828__A1 _3883_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3516__B1 _5322_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4939__S0 _5404_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3351__A _4276_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5977__S _5977_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4881__S _5101_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4980_ _6260_/Q _6195_/Q _6219_/Q _6112_/Q _5100_/S0 _5100_/S1 vssd1 vssd1 vccd1
+ vccd1 _4980_/X sky130_fd_sc_hd__mux4_1
X_3931_ _3770_/A _5267_/B _5264_/B _4115_/A _3930_/X vssd1 vssd1 vccd1 vccd1 _3938_/A
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5278__A _6461_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3862_ _3860_/X _3861_/X _3883_/S vssd1 vssd1 vccd1 vccd1 _3862_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_61_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5601_ _5601_/A _5601_/B vssd1 vssd1 vccd1 vccd1 _5601_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5532_ _5532_/A _5532_/B vssd1 vssd1 vccd1 vccd1 _5534_/A sky130_fd_sc_hd__nor2_1
X_3793_ _3816_/B _3885_/A _3884_/S vssd1 vssd1 vccd1 vccd1 _3793_/X sky130_fd_sc_hd__and3_4
XFILLER_0_14_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5463_ hold607/X _5462_/X _5513_/S vssd1 vssd1 vccd1 vccd1 _5463_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5394_ _3072_/Y _4948_/S _5645_/A _5644_/A vssd1 vssd1 vccd1 vccd1 _5394_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_1_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4414_ _4414_/A _4414_/B vssd1 vssd1 vccd1 vccd1 _4414_/Y sky130_fd_sc_hd__nor2_1
X_4345_ _4338_/A _4268_/Y _5370_/B _5605_/C vssd1 vssd1 vccd1 vccd1 _4345_/X sky130_fd_sc_hd__o211a_1
XANTENNA__4180__B1 _4463_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4276_ _4276_/A _5314_/S vssd1 vssd1 vccd1 vccd1 _4276_/X sky130_fd_sc_hd__or2_1
X_3227_ _3168_/B _3229_/A _3057_/Y _3205_/X vssd1 vssd1 vccd1 vccd1 _3227_/Y sky130_fd_sc_hd__a31oi_1
XANTENNA__3261__A _3581_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6015_ input7/X hold624/X _6019_/S vssd1 vssd1 vccd1 vccd1 _6461_/D sky130_fd_sc_hd__mux2_1
X_3158_ _4359_/C _3249_/B _3300_/B vssd1 vssd1 vccd1 vccd1 _3527_/B sky130_fd_sc_hd__a21o_1
XANTENNA__5887__S _5887_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3089_ _4670_/B vssd1 vssd1 vccd1 vccd1 _6033_/B sky130_fd_sc_hd__inv_2
XFILLER_0_92_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5983__A1 _5995_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_5_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold370 _5037_/X vssd1 vssd1 vccd1 vccd1 _6328_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold381 _6323_/Q vssd1 vssd1 vccd1 vccd1 hold381/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold392 _5537_/X vssd1 vssd1 vccd1 vccd1 _6370_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4267__A _4313_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_11_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6439_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_43_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4130_ _4130_/A vssd1 vssd1 vccd1 vccd1 _4132_/A sky130_fd_sc_hd__inv_2
X_4061_ _4199_/A _6382_/Q vssd1 vssd1 vccd1 vccd1 _4063_/C sky130_fd_sc_hd__and2_1
XANTENNA__4177__A _6067_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4905__A _6366_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4963_ _6309_/Q _4963_/B vssd1 vssd1 vccd1 vccd1 _4963_/X sky130_fd_sc_hd__and2_1
X_3914_ _4150_/A _6379_/Q vssd1 vssd1 vccd1 vccd1 _3917_/C sky130_fd_sc_hd__and2b_1
XFILLER_0_80_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4894_ _5817_/A _4893_/X _4882_/X vssd1 vssd1 vccd1 vccd1 _4894_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_6_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3955__S _4241_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3845_ _6230_/Q _3731_/X _3804_/X _6453_/Q vssd1 vssd1 vccd1 vccd1 _3846_/C sky130_fd_sc_hd__a22o_1
XFILLER_0_27_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3776_ _6345_/Q _6343_/Q _5136_/A _6346_/Q vssd1 vssd1 vccd1 vccd1 _4223_/A sky130_fd_sc_hd__and4b_4
XANTENNA_fanout127_A _4300_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5515_ _6483_/Q _4962_/B _5593_/S vssd1 vssd1 vccd1 vccd1 _5517_/B sky130_fd_sc_hd__mux2_1
XANTENNA__3256__A _3304_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5446_ hold583/X _5520_/B _5445_/X _5415_/X vssd1 vssd1 vccd1 vccd1 _5446_/X sky130_fd_sc_hd__a22o_1
Xfanout102 _5499_/S vssd1 vssd1 vccd1 vccd1 _5783_/A sky130_fd_sc_hd__buf_4
X_5377_ _5364_/A _5607_/B2 _5376_/X _3699_/A vssd1 vssd1 vccd1 vccd1 _5377_/Y sky130_fd_sc_hd__a22oi_4
Xfanout113 _6108_/S vssd1 vssd1 vccd1 vccd1 _5769_/S sky130_fd_sc_hd__clkbuf_8
Xfanout146 hold574/X vssd1 vssd1 vccd1 vccd1 _5605_/C sky130_fd_sc_hd__buf_4
Xfanout135 _4313_/A vssd1 vssd1 vccd1 vccd1 _4338_/A sky130_fd_sc_hd__buf_4
X_4328_ _4328_/A _4328_/B vssd1 vssd1 vccd1 vccd1 _4328_/X sky130_fd_sc_hd__or2_1
Xfanout124 hold526/X vssd1 vssd1 vccd1 vccd1 _5384_/A sky130_fd_sc_hd__buf_6
XFILLER_0_10_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout157 hold646/X vssd1 vssd1 vccd1 vccd1 _3284_/B sky130_fd_sc_hd__clkbuf_4
X_4259_ _4260_/B _5388_/A _4325_/A vssd1 vssd1 vccd1 vccd1 _4259_/X sky130_fd_sc_hd__and3b_1
Xfanout179 fanout180/X vssd1 vssd1 vccd1 vccd1 fanout179/X sky130_fd_sc_hd__clkbuf_8
Xfanout168 hold641/X vssd1 vssd1 vccd1 vccd1 _5078_/S1 sky130_fd_sc_hd__buf_6
XANTENNA__4456__B2 _4441_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4208__A1 _6290_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5956__B2 _5977_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold506_A _6289_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3195__A1 _5605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4695__A1 _4715_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3958__B1 _3795_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3422__A2 _3674_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3630_ _3489_/B hold192/X _6130_/Q _6432_/Q _3629_/Y vssd1 vssd1 vccd1 vccd1 _3630_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_50_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3561_ _5777_/A _3619_/C vssd1 vssd1 vccd1 vccd1 _3561_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_70_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5300_ _5299_/X _3891_/Y _5300_/C _5300_/D vssd1 vssd1 vccd1 vccd1 _5300_/X sky130_fd_sc_hd__and4bb_1
X_3492_ _3492_/A _3492_/B _3492_/C _3492_/D vssd1 vssd1 vccd1 vccd1 _3492_/X sky130_fd_sc_hd__or4_1
X_6280_ _6336_/CLK _6280_/D fanout182/X vssd1 vssd1 vccd1 vccd1 _6280_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_0_59_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4686__A1 _6286_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5231_ _4029_/Y _5230_/X _5292_/S vssd1 vssd1 vccd1 vccd1 _5231_/X sky130_fd_sc_hd__mux2_1
X_5162_ _5162_/A _5162_/B vssd1 vssd1 vccd1 vccd1 _5164_/A sky130_fd_sc_hd__xor2_1
XANTENNA__3523__B _5384_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4113_ _6289_/Q _3770_/A _3773_/Y _5174_/B vssd1 vssd1 vccd1 vccd1 _4113_/X sky130_fd_sc_hd__a22o_1
X_5093_ _6375_/Q _5848_/S _5972_/B1 _5092_/X vssd1 vssd1 vccd1 vccd1 _5093_/Y sky130_fd_sc_hd__a22oi_1
X_4044_ _3814_/Y _3948_/B _3962_/B _4036_/B _4190_/A vssd1 vssd1 vccd1 vccd1 _4044_/X
+ sky130_fd_sc_hd__o41a_1
XANTENNA__5938__A1 _6425_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5995_ _5988_/B _5995_/B _5995_/C _5995_/D vssd1 vssd1 vccd1 vccd1 _5995_/X sky130_fd_sc_hd__and4b_1
XFILLER_0_19_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4610__A1 _5757_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4946_ _6368_/Q _4922_/X _4968_/B _4808_/Y _4924_/C vssd1 vssd1 vccd1 vccd1 _4946_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA__5466__A _5492_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4877_ _4312_/A _5783_/A _4875_/X _4876_/X vssd1 vssd1 vccd1 vccd1 _4877_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_15_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3828_ _3883_/S _3825_/X _3827_/X vssd1 vssd1 vccd1 vccd1 _3830_/B sky130_fd_sc_hd__o21a_1
X_3759_ _6343_/Q _3928_/B vssd1 vssd1 vccd1 vccd1 _3759_/Y sky130_fd_sc_hd__nor2_4
XFILLER_0_42_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6478_ _6481_/CLK _6478_/D fanout176/X vssd1 vssd1 vccd1 vccd1 _6478_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA__4677__A1 _6284_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5429_ _5492_/A _5429_/B _5429_/C vssd1 vssd1 vccd1 vccd1 _5429_/X sky130_fd_sc_hd__and3_1
XANTENNA__4126__B1 _3807_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4248__C _4248_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5095__B _5771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4365__A0 _4919_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5880__A3 _5866_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output40_A _6332_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6481__SET_B fanout176/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4800_ _6361_/Q _6413_/Q _4800_/S vssd1 vssd1 vccd1 vccd1 _4800_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4605__D _4611_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5780_ _4324_/B _3530_/A _5995_/C vssd1 vssd1 vccd1 vccd1 _5780_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_8_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4731_ _6310_/Q _4719_/A _4730_/X _4957_/S vssd1 vssd1 vccd1 vccd1 _4731_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5935__A4 _6424_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4662_ input6/X _4668_/B vssd1 vssd1 vccd1 vccd1 _4662_/X sky130_fd_sc_hd__and2_1
XANTENNA__5148__A2 _6334_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3613_ _5346_/A _3364_/Y _3405_/A vssd1 vssd1 vccd1 vccd1 _5310_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_43_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6401_ _6483_/CLK hold12/X vssd1 vssd1 vccd1 vccd1 hold11/A sky130_fd_sc_hd__dfxtp_1
X_4593_ _4675_/A _4259_/X _3424_/B _3590_/A vssd1 vssd1 vccd1 vccd1 _4593_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3544_ _3419_/B _3525_/Y _3543_/X vssd1 vssd1 vccd1 vccd1 _3544_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_3_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6332_ _6419_/CLK _6332_/D fanout170/X vssd1 vssd1 vccd1 vccd1 _6332_/Q sky130_fd_sc_hd__dfrtp_2
X_3475_ _5995_/C _4363_/A vssd1 vssd1 vccd1 vccd1 _3488_/A sky130_fd_sc_hd__nor2_1
X_6263_ _6263_/CLK _6263_/D vssd1 vssd1 vccd1 vccd1 _6263_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5214_ _5214_/A _5214_/B vssd1 vssd1 vccd1 vccd1 _5215_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_86_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6194_ _6399_/CLK _6194_/D vssd1 vssd1 vccd1 vccd1 _6194_/Q sky130_fd_sc_hd__dfxtp_1
X_5145_ _5145_/A _5146_/C _6021_/S _5145_/D vssd1 vssd1 vccd1 vccd1 _5291_/S sky130_fd_sc_hd__or4_4
XFILLER_0_98_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5076_ _6407_/Q _5075_/X _6070_/A vssd1 vssd1 vccd1 vccd1 _5076_/X sky130_fd_sc_hd__mux2_1
X_4027_ _4027_/A _4087_/B vssd1 vssd1 vccd1 vccd1 _4027_/X sky130_fd_sc_hd__and2_1
XFILLER_0_79_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4831__B2 _4924_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4831__A1 _5109_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5978_ _5995_/C _5978_/B vssd1 vssd1 vccd1 vccd1 _5978_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_19_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4929_ _4929_/A _4929_/B _4929_/C vssd1 vssd1 vccd1 vccd1 _4929_/X sky130_fd_sc_hd__or3_1
XANTENNA__5139__A2 _4150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3444__A _4325_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4259__B _5388_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4822__A1 _4919_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4214__S _6334_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3619__A _5322_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4050__A2 _3731_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5834__A _5866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4889__A1 _6462_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4889__B2 _5109_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3260_ _3172_/A _3204_/X _3225_/X _3230_/Y _3219_/Y vssd1 vssd1 vccd1 vccd1 _3261_/C
+ sky130_fd_sc_hd__o32a_1
XANTENNA__3849__C1 _3883_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3191_ _3229_/A _3547_/B vssd1 vssd1 vccd1 vccd1 _3232_/C sky130_fd_sc_hd__nor2_1
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3801__B _3818_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4274__C1 _5388_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5901_ _5901_/A _5901_/B vssd1 vssd1 vccd1 vccd1 _5912_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_72_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6015__A0 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6372__RESET_B fanout172/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5832_ _5976_/S _5827_/Y _5831_/Y _5786_/Y vssd1 vssd1 vccd1 vccd1 _5832_/X sky130_fd_sc_hd__a22o_1
XANTENNA__6301__RESET_B fanout183/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5763_ _6314_/Q hold502/X _5765_/S vssd1 vssd1 vccd1 vccd1 _5763_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_29_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4714_ _4227_/X _4713_/X _4714_/S vssd1 vssd1 vccd1 vccd1 _4714_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6339__SET_B fanout185/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5694_ _6222_/Q _5721_/A2 _4235_/S _6115_/Q _5730_/C1 vssd1 vssd1 vccd1 vccd1 _5696_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_16_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4645_ _5393_/A1 _5268_/A _4582_/Y _4644_/X vssd1 vssd1 vccd1 vccd1 _4645_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_44_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4576_ _4595_/B _4264_/X _5364_/A vssd1 vssd1 vccd1 vccd1 _4576_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_4_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3552__A1 _3525_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3527_ _3699_/A _3527_/B _3527_/C vssd1 vssd1 vccd1 vccd1 _3527_/X sky130_fd_sc_hd__and3_1
X_6315_ _6316_/CLK _6315_/D fanout174/X vssd1 vssd1 vccd1 vccd1 _6315_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_0_4_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_39_wb_clk_i_A clkbuf_leaf_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_6246_ _6248_/CLK _6246_/D fanout180/X vssd1 vssd1 vccd1 vccd1 _6246_/Q sky130_fd_sc_hd__dfrtp_1
X_3458_ _5607_/B2 _3450_/B _3457_/X vssd1 vssd1 vccd1 vccd1 _3458_/X sky130_fd_sc_hd__a21bo_1
X_3389_ _6359_/Q _3390_/B vssd1 vssd1 vccd1 vccd1 _4354_/B sky130_fd_sc_hd__nor2_1
X_6177_ _6456_/CLK _6177_/D vssd1 vssd1 vccd1 vccd1 _6177_/Q sky130_fd_sc_hd__dfxtp_1
X_5128_ hold514/X _4555_/Y _5127_/X vssd1 vssd1 vccd1 vccd1 _5128_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_98_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3607__A2 _3281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5059_ _5058_/X _5101_/S vssd1 vssd1 vccd1 vccd1 _5059_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_79_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold419_A _6385_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4032__A2 _3799_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4583__A3 _3489_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5780__A2 _3530_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3791__A1 _5607_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3543__B2 _5384_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4099__A2 _6289_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_36_wb_clk_i clkbuf_leaf_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6376_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_30_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold60 hold60/A vssd1 vssd1 vccd1 vccd1 hold60/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 hold82/A vssd1 vssd1 vccd1 vccd1 hold82/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 hold71/A vssd1 vssd1 vccd1 vccd1 hold71/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold93 hold93/A vssd1 vssd1 vccd1 vccd1 hold93/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_2 _3387_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4430_ _4430_/A _4430_/B vssd1 vssd1 vccd1 vccd1 _4431_/B sky130_fd_sc_hd__nor2_1
X_4361_ _6100_/A _4361_/B vssd1 vssd1 vccd1 vccd1 _4363_/B sky130_fd_sc_hd__or2_1
XFILLER_0_6_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6100_ _6100_/A _6100_/B vssd1 vssd1 vccd1 vccd1 _6100_/X sky130_fd_sc_hd__or2_1
XANTENNA__5287__A1 _6340_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3312_ _5346_/A _5370_/B vssd1 vssd1 vccd1 vccd1 _3411_/A sky130_fd_sc_hd__nor2_1
X_4292_ _4313_/A _4303_/A _5418_/A vssd1 vssd1 vccd1 vccd1 _4296_/B sky130_fd_sc_hd__and3_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3243_ _5387_/A _3304_/B vssd1 vssd1 vccd1 vccd1 _5374_/B sky130_fd_sc_hd__nor2_1
XANTENNA__3298__B1 _5866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6031_ hold45/X _6026_/S _6023_/Y hold77/X vssd1 vssd1 vccd1 vccd1 hold78/A sky130_fd_sc_hd__a22o_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3837__A2 _3731_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3174_ _4557_/D _3174_/B vssd1 vssd1 vccd1 vccd1 _3174_/X sky130_fd_sc_hd__and2_1
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4798__B1 _4963_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5815_ _6415_/Q _5892_/S _4841_/X vssd1 vssd1 vccd1 vccd1 _5815_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_36_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3259__A _4557_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5746_ hold27/X _3839_/B _6104_/S vssd1 vssd1 vccd1 vccd1 hold28/A sky130_fd_sc_hd__mux2_1
XFILLER_0_17_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4970__A0 _6458_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5677_ _6336_/Q _5628_/X _5643_/X _6424_/Q vssd1 vssd1 vccd1 vccd1 _5687_/B sky130_fd_sc_hd__a22o_1
X_4628_ hold442/X _4604_/X _4605_/X _6487_/Q _4627_/X vssd1 vssd1 vccd1 vccd1 _4628_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5193__B _6289_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold530 _4620_/X vssd1 vssd1 vccd1 vccd1 _6286_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4559_ _5783_/A _4559_/B vssd1 vssd1 vccd1 vccd1 _5288_/S sky130_fd_sc_hd__nor2_2
Xhold541 _6371_/Q vssd1 vssd1 vccd1 vccd1 hold541/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold563 _5581_/X vssd1 vssd1 vccd1 vccd1 _6374_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold552 _6425_/Q vssd1 vssd1 vccd1 vccd1 _5933_/A sky130_fd_sc_hd__buf_1
XFILLER_0_40_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold574 _6298_/Q vssd1 vssd1 vccd1 vccd1 hold574/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold585 _6346_/Q vssd1 vssd1 vccd1 vccd1 hold585/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold596 _5476_/X vssd1 vssd1 vccd1 vccd1 _6365_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6229_ _6452_/CLK _6229_/D vssd1 vssd1 vccd1 vccd1 _6229_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4238__C1 _5655_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3367__B1_N _6339_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4410__C1 _5730_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5384__A _5384_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4939__S1 _5078_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput50 _3074_/Y vssd1 vssd1 vccd1 vccd1 io_out[32] sky130_fd_sc_hd__buf_12
XANTENNA__3632__A _4276_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3819__A2 _3793_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3351__B _4325_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3930_ _3927_/Y _3928_/Y _3929_/X _3759_/Y vssd1 vssd1 vccd1 vccd1 _3930_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_53_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3452__B1 _5777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5278__B _6460_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3079__A _6285_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3861_ _6451_/Q _6228_/Q _3861_/S vssd1 vssd1 vccd1 vccd1 _3861_/X sky130_fd_sc_hd__mux2_1
X_5600_ _5600_/A _5600_/B _5600_/C vssd1 vssd1 vccd1 vccd1 _5601_/B sky130_fd_sc_hd__and3_1
XFILLER_0_6_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3792_ _3892_/A vssd1 vssd1 vccd1 vccd1 _4052_/A sky130_fd_sc_hd__inv_2
X_5531_ _5531_/A _5531_/B vssd1 vssd1 vccd1 vccd1 _5532_/B sky130_fd_sc_hd__and2_1
XFILLER_0_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3807__A _3852_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4910__B _4930_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5462_ _6461_/Q _5461_/X _5512_/S vssd1 vssd1 vccd1 vccd1 _5462_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4704__B1 _4714_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5393_ _5393_/A1 hold405/X _3541_/C _5362_/A vssd1 vssd1 vccd1 vccd1 _5393_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_78_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4413_ _5299_/A _5299_/B vssd1 vssd1 vccd1 vccd1 _4414_/B sky130_fd_sc_hd__xnor2_1
X_4344_ _4344_/A _4344_/B vssd1 vssd1 vccd1 vccd1 _4344_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_1_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4275_ _5398_/A _5774_/A _5317_/B _4250_/X _4274_/X vssd1 vssd1 vccd1 vccd1 _4275_/X
+ sky130_fd_sc_hd__a311o_1
X_6014_ _4658_/A hold626/X _6019_/S vssd1 vssd1 vccd1 vccd1 _6460_/D sky130_fd_sc_hd__mux2_1
X_3226_ _3547_/B _3282_/A _3219_/Y _3225_/X vssd1 vssd1 vccd1 vccd1 _3226_/X sky130_fd_sc_hd__o31a_1
XFILLER_0_94_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3157_ _4268_/A _4248_/B _3249_/B vssd1 vssd1 vccd1 vccd1 _3300_/B sky130_fd_sc_hd__and3_1
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3088_ _3088_/A vssd1 vssd1 vccd1 vccd1 _6032_/C sky130_fd_sc_hd__inv_2
XFILLER_0_49_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5729_ _6316_/Q _5630_/X _5653_/X _6490_/Q vssd1 vssd1 vccd1 vccd1 _5737_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_45_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4820__B _4919_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4171__A1 _4332_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold371 _6321_/Q vssd1 vssd1 vccd1 vccd1 hold371/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold360 _5762_/X vssd1 vssd1 vccd1 vccd1 _6406_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold382 _4936_/X vssd1 vssd1 vccd1 vccd1 _6323_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold393 _6124_/Q vssd1 vssd1 vccd1 vccd1 _4312_/B sky130_fd_sc_hd__buf_1
XFILLER_0_99_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3682__B1 _5387_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4283__A _4605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4934__A0 _6367_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3627__A _5322_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5111__A0 _6409_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4060_ _6288_/Q _4060_/B _4063_/B vssd1 vssd1 vccd1 vccd1 _4070_/A sky130_fd_sc_hd__or3b_1
XFILLER_0_3_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5662__A1 _6310_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5414__A1 _5478_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4193__A _5268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4962_ _5102_/A _4962_/B vssd1 vssd1 vccd1 vccd1 _4962_/Y sky130_fd_sc_hd__nand2_1
X_3913_ _6379_/Q _4150_/A vssd1 vssd1 vccd1 vccd1 _3917_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_86_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4893_ _6365_/Q _5816_/S _5842_/B1 _4892_/X vssd1 vssd1 vccd1 vccd1 _4893_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_80_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3844_ _3883_/S _3841_/X _3843_/X vssd1 vssd1 vccd1 vccd1 _3846_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_61_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5717__A2 _6355_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3775_ _3770_/A _5267_/A _3773_/Y _6284_/Q vssd1 vssd1 vccd1 vccd1 _3775_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_42_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5514_ _5508_/A _5505_/Y _5507_/B vssd1 vssd1 vccd1 vccd1 _5519_/A sky130_fd_sc_hd__o21a_1
X_5445_ _5445_/A _5445_/B vssd1 vssd1 vccd1 vccd1 _5445_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_66_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5376_ _5375_/X _4335_/B _5376_/S vssd1 vssd1 vccd1 vccd1 _5376_/X sky130_fd_sc_hd__mux2_1
Xfanout103 _3390_/X vssd1 vssd1 vccd1 vccd1 _4948_/S sky130_fd_sc_hd__buf_6
XFILLER_0_10_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout147 hold648/X vssd1 vssd1 vccd1 vccd1 _5605_/B sky130_fd_sc_hd__buf_4
Xfanout125 _4715_/B2 vssd1 vssd1 vccd1 vccd1 _5757_/B sky130_fd_sc_hd__buf_4
X_4327_ _5315_/A _4326_/Y _5605_/D vssd1 vssd1 vccd1 vccd1 _4327_/X sky130_fd_sc_hd__a21o_1
Xfanout136 _4313_/A vssd1 vssd1 vccd1 vccd1 _3665_/A sky130_fd_sc_hd__buf_6
Xfanout114 _6108_/S vssd1 vssd1 vccd1 vccd1 _5513_/S sky130_fd_sc_hd__clkbuf_4
Xfanout158 _4782_/A vssd1 vssd1 vccd1 vccd1 _3323_/A sky130_fd_sc_hd__buf_4
XANTENNA__3703__C _4150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4258_ _4782_/A _4324_/B _4244_/Y _4257_/X _5607_/B2 vssd1 vssd1 vccd1 vccd1 _4258_/X
+ sky130_fd_sc_hd__a221o_1
Xfanout169 _6128_/Q vssd1 vssd1 vccd1 vccd1 _5101_/S sky130_fd_sc_hd__buf_8
X_3209_ _3304_/B _3514_/B vssd1 vssd1 vccd1 vccd1 _5317_/A sky130_fd_sc_hd__or2_2
XANTENNA__3664__B1 _4325_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4189_ _4189_/A _4189_/B vssd1 vssd1 vccd1 vccd1 _4190_/B sky130_fd_sc_hd__or2_1
XFILLER_0_96_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5956__A2 _5785_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5169__A0 _6335_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5708__A2 _5721_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3195__A2 _3304_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4977__S _5016_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3881__S _3884_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3498__A3 _3497_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5892__A1 _6421_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold190 _6199_/Q vssd1 vssd1 vccd1 vccd1 hold190/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3101__1 _6467_/CLK vssd1 vssd1 vccd1 vccd1 _6165_/CLK sky130_fd_sc_hd__inv_2
XANTENNA__4907__B1 _4924_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3560_ _3557_/X _3559_/X _3786_/A vssd1 vssd1 vccd1 vccd1 _3560_/X sky130_fd_sc_hd__a21o_1
XANTENNA__5580__A0 _6463_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5275__C _6408_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4887__S _4948_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3491_ _3493_/A hold47/X _3493_/C hold39/X _3472_/B vssd1 vssd1 vccd1 vccd1 _3492_/D
+ sky130_fd_sc_hd__o41a_1
X_5230_ _5147_/C _5225_/X _5229_/X _5221_/X vssd1 vssd1 vccd1 vccd1 _5230_/X sky130_fd_sc_hd__a31o_1
X_5161_ _5161_/A _5257_/B vssd1 vssd1 vccd1 vccd1 _5165_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__3092__A _6312_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3804__B _3883_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4112_ _5174_/B vssd1 vssd1 vccd1 vccd1 _5173_/B sky130_fd_sc_hd__inv_2
XFILLER_0_75_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5092_ _6408_/Q _5091_/X _5971_/S vssd1 vssd1 vccd1 vccd1 _5092_/X sky130_fd_sc_hd__mux2_1
X_4043_ _4042_/X hold285/X _4241_/S vssd1 vssd1 vccd1 vccd1 _6114_/D sky130_fd_sc_hd__mux2_1
XANTENNA__5511__S _5567_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5994_ _3480_/B _3636_/B _3635_/Y _5993_/X vssd1 vssd1 vccd1 vccd1 _6433_/D sky130_fd_sc_hd__a22o_1
XANTENNA__4354__C _5644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4945_ _4945_/A _4945_/B vssd1 vssd1 vccd1 vccd1 _4968_/B sky130_fd_sc_hd__nand2_1
XANTENNA__6060__A1 _4366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4876_ _6364_/Q _5863_/S _6070_/A vssd1 vssd1 vccd1 vccd1 _4876_/X sky130_fd_sc_hd__o21a_1
X_3827_ _3885_/A _3826_/X _3852_/A vssd1 vssd1 vccd1 vccd1 _3827_/X sky130_fd_sc_hd__o21a_1
X_3758_ _3774_/A _6345_/Q _5136_/A vssd1 vssd1 vccd1 vccd1 _3928_/B sky130_fd_sc_hd__or3_2
XFILLER_0_15_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3582__C1 _3619_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3689_ _3302_/X _3675_/X _3677_/X _3669_/Y vssd1 vssd1 vccd1 vccd1 _3689_/Y sky130_fd_sc_hd__a31oi_4
X_6477_ _6481_/CLK _6477_/D fanout176/X vssd1 vssd1 vccd1 vccd1 _6477_/Q sky130_fd_sc_hd__dfstp_1
X_5428_ _6476_/Q _4822_/X _5478_/S vssd1 vssd1 vccd1 vccd1 _5429_/C sky130_fd_sc_hd__mux2_1
XFILLER_0_100_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5359_ _3187_/X _3254_/Y _5350_/Y _4313_/A vssd1 vssd1 vccd1 vccd1 _5359_/X sky130_fd_sc_hd__o31a_1
XANTENNA__5626__B2 _6435_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_hold616_A _6458_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3573__C1 _5322_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5314__A0 _5360_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4500__S _4500_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3624__B _5757_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3340__A2 _3673_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6042__A1 _5567_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4730_ _6310_/Q _4720_/X _5224_/A2 hold436/X vssd1 vssd1 vccd1 vccd1 _4730_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_16_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4661_ _4217_/A _4652_/X _4654_/Y _4660_/X vssd1 vssd1 vccd1 vccd1 _6296_/D sky130_fd_sc_hd__o22a_1
XFILLER_0_43_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3612_ _3205_/B _4357_/C _3281_/A _3434_/B vssd1 vssd1 vccd1 vccd1 _5307_/C sky130_fd_sc_hd__a31o_1
XFILLER_0_9_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6400_ _6400_/CLK hold8/X vssd1 vssd1 vccd1 vccd1 hold7/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4592_ _4250_/X _4586_/X _4590_/X _4591_/X _5600_/A vssd1 vssd1 vccd1 vccd1 _4592_/X
+ sky130_fd_sc_hd__o311a_2
X_6331_ _6426_/CLK _6331_/D fanout171/X vssd1 vssd1 vccd1 vccd1 _6331_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_101_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3543_ _3110_/A _3176_/Y _3541_/C hold599/X _5384_/A vssd1 vssd1 vccd1 vccd1 _3543_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA_clkbuf_leaf_29_wb_clk_i_A clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_24_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3474_ _3493_/A _3472_/B _3487_/B _3473_/X vssd1 vssd1 vccd1 vccd1 _3474_/X sky130_fd_sc_hd__a22o_1
X_6262_ _6265_/CLK _6262_/D vssd1 vssd1 vccd1 vccd1 _6262_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4659__A2 _4652_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5213_ _5213_/A _5213_/B vssd1 vssd1 vccd1 vccd1 _5214_/B sky130_fd_sc_hd__xnor2_1
XANTENNA_clkbuf_2_2__f_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6193_ _6456_/CLK _6193_/D vssd1 vssd1 vccd1 vccd1 _6193_/Q sky130_fd_sc_hd__dfxtp_1
X_5144_ hold643/X _5143_/X _5232_/S vssd1 vssd1 vccd1 vccd1 _6333_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_19_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3550__A _5605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5075_ _6463_/Q _5074_/X _5974_/S vssd1 vssd1 vccd1 vccd1 _5075_/X sky130_fd_sc_hd__mux2_1
X_4026_ _6461_/Q _5221_/B _6347_/Q vssd1 vssd1 vccd1 vccd1 _4026_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_29_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5977_ _5969_/A _5976_/X _5977_/S vssd1 vssd1 vccd1 vccd1 _5977_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5477__A _5757_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4928_ _6464_/Q _4963_/B _4926_/X _5109_/A1 vssd1 vssd1 vccd1 vccd1 _4929_/C sky130_fd_sc_hd__a22o_1
XFILLER_0_47_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4347__A1 _3284_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4859_ _3091_/Y _4957_/S _4858_/X vssd1 vssd1 vccd1 vccd1 _4859_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__6248__RESET_B fanout180/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6529_ _6529_/A vssd1 vssd1 vccd1 vccd1 _6529_/X sky130_fd_sc_hd__buf_1
XFILLER_0_15_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3444__B _5777_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold399_A _6384_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4259__C _4325_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold566_A _6431_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3953__S0 _5721_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4556__A _6159_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4291__A _5605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4889__A2 _4963_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5834__B _6462_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3635__A _4800_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3190_ _3627_/B _3414_/B _3376_/B _4557_/C vssd1 vssd1 vccd1 vccd1 _3190_/X sky130_fd_sc_hd__a211o_1
XANTENNA__5697__S0 _5655_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4274__B1 _5362_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5900_ hold588/X _5899_/X _5977_/S vssd1 vssd1 vccd1 vccd1 _5900_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_76_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4026__A0 _6461_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5831_ _6364_/Q _5974_/S _5830_/X vssd1 vssd1 vccd1 vccd1 _5831_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__4405__S _4464_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5762_ _6313_/Q hold359/X _5765_/S vssd1 vssd1 vccd1 vccd1 _5762_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_29_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4713_ _4713_/A _4713_/B vssd1 vssd1 vccd1 vccd1 _4713_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_6_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6377_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_8_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5693_ _5693_/A _5693_/B vssd1 vssd1 vccd1 vccd1 _5693_/X sky130_fd_sc_hd__or2_1
XANTENNA__4329__B2 _5605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4644_ hold578/X _4604_/X _4605_/X hold594/X _4643_/X vssd1 vssd1 vccd1 vccd1 _4644_/X
+ sky130_fd_sc_hd__a221o_1
X_4575_ hold446/X _6340_/Q _4575_/S vssd1 vssd1 vccd1 vccd1 _4575_/X sky130_fd_sc_hd__mux2_1
X_3526_ _5384_/A hold328/X _4264_/B _3525_/Y _3524_/X vssd1 vssd1 vccd1 vccd1 _3526_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout102_A _5499_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6314_ _6336_/CLK _6314_/D fanout182/X vssd1 vssd1 vccd1 vccd1 _6314_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_0_24_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6245_ _6248_/CLK hold38/X fanout180/X vssd1 vssd1 vccd1 vccd1 hold37/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5829__A1 _6364_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3457_ _5315_/B _3457_/B vssd1 vssd1 vccd1 vccd1 _3457_/X sky130_fd_sc_hd__or2_1
X_3388_ _3530_/A _3497_/B _3665_/A vssd1 vssd1 vccd1 vccd1 _3388_/X sky130_fd_sc_hd__o21a_1
X_6176_ _6452_/CLK hold98/X vssd1 vssd1 vccd1 vccd1 hold97/A sky130_fd_sc_hd__dfxtp_1
X_5127_ _6333_/Q _5244_/S _5126_/Y _5123_/A vssd1 vssd1 vccd1 vccd1 _5127_/X sky130_fd_sc_hd__a211o_1
X_5058_ _6156_/Q _6147_/Q _6139_/Q _6183_/Q _5100_/S0 _5100_/S1 vssd1 vssd1 vccd1
+ vccd1 _5058_/X sky130_fd_sc_hd__mux4_1
X_4009_ _5136_/B _4003_/X _4007_/A _3753_/X vssd1 vssd1 vccd1 vccd1 _4009_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_79_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4568__A1 _6333_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5765__A0 _6316_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4099__A3 _6383_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4985__S _5105_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold50 hold50/A vssd1 vssd1 vccd1 vccd1 hold50/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 hold83/A vssd1 vssd1 vccd1 vccd1 hold83/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold72 hold72/A vssd1 vssd1 vccd1 vccd1 hold72/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold61 hold61/A vssd1 vssd1 vccd1 vccd1 hold61/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 hold94/A vssd1 vssd1 vccd1 vccd1 hold94/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_85_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_3 _6067_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4360_ _5600_/A _4360_/B vssd1 vssd1 vccd1 vccd1 _4360_/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_6_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5056__S _6070_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4731__A1 _6310_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3311_ _3326_/B _3311_/B vssd1 vssd1 vccd1 vccd1 _5370_/B sky130_fd_sc_hd__nor2_4
XFILLER_0_1_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4731__B2 _4957_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4291_ _5605_/B _5757_/A _4768_/S vssd1 vssd1 vccd1 vccd1 _4310_/S sky130_fd_sc_hd__or3b_4
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3242_ _3180_/B _3240_/X _3241_/X vssd1 vssd1 vccd1 vccd1 _3273_/A sky130_fd_sc_hd__o21a_1
XANTENNA__3298__A1 _4313_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6030_ hold77/X _6026_/S _6023_/Y _3700_/A vssd1 vssd1 vccd1 vccd1 _6030_/X sky130_fd_sc_hd__a22o_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3173_ _4782_/A _3172_/Y _3326_/A vssd1 vssd1 vccd1 vccd1 _3174_/B sky130_fd_sc_hd__mux2_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5692__C1 _5721_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4798__A1 _5413_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4798__B2 _6458_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5814_ _5826_/B _5814_/B vssd1 vssd1 vccd1 vccd1 _5814_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_8_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3222__A1 _3168_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5745_ hold3/X _3847_/B _6104_/S vssd1 vssd1 vccd1 vccd1 hold4/A sky130_fd_sc_hd__mux2_1
XFILLER_0_29_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5676_ _6478_/Q _5629_/X _5646_/X hold375/X vssd1 vssd1 vccd1 vccd1 _5687_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_4_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4627_ _6462_/Q _4606_/X _4607_/X _6313_/Q vssd1 vssd1 vccd1 vccd1 _4627_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4722__A1 _6309_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold520 _6484_/Q vssd1 vssd1 vccd1 vccd1 hold520/X sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA__4722__B2 _5783_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4558_ wire92/X vssd1 vssd1 vccd1 vccd1 _4559_/B sky130_fd_sc_hd__inv_2
Xhold542 _5549_/X vssd1 vssd1 vccd1 vccd1 _6371_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold531 _6375_/Q vssd1 vssd1 vccd1 vccd1 hold531/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold553 _5944_/X vssd1 vssd1 vccd1 vccd1 _6425_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold564 _6285_/Q vssd1 vssd1 vccd1 vccd1 hold564/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold575 _3360_/B vssd1 vssd1 vccd1 vccd1 hold575/X sky130_fd_sc_hd__dlygate4sd3_1
X_3509_ _4324_/B hold347/X _3554_/A _5398_/B _3527_/C vssd1 vssd1 vccd1 vccd1 _3509_/X
+ sky130_fd_sc_hd__o41a_1
Xhold586 _6423_/Q vssd1 vssd1 vccd1 vccd1 hold586/X sky130_fd_sc_hd__dlygate4sd3_1
X_4489_ _4138_/X hold190/X _4491_/S vssd1 vssd1 vccd1 vccd1 _4489_/X sky130_fd_sc_hd__mux2_1
Xhold597 _6489_/Q vssd1 vssd1 vccd1 vccd1 hold597/X sky130_fd_sc_hd__buf_1
XANTENNA__5490__A _5757_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6228_ _6456_/CLK _6228_/D vssd1 vssd1 vccd1 vccd1 _6228_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6159_ _6474_/CLK _6159_/D fanout179/X vssd1 vssd1 vccd1 vccd1 _6159_/Q sky130_fd_sc_hd__dfstp_4
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5921__A1_N _5977_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold431_A _6435_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold529_A _6286_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3169__B _4557_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3884__S _3884_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput51 _3662_/X vssd1 vssd1 vccd1 vccd1 io_out[33] sky130_fd_sc_hd__buf_12
Xoutput40 _6332_/Q vssd1 vssd1 vccd1 vccd1 io_out[21] sky130_fd_sc_hd__buf_12
XFILLER_0_31_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3632__B _6159_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5426__C1 _5478_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5278__C _6465_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3860_ _6204_/Q _6212_/Q _3861_/S vssd1 vssd1 vccd1 vccd1 _3860_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_66_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3791_ _5607_/B2 _3789_/X _3790_/X _3788_/Y vssd1 vssd1 vccd1 vccd1 _3791_/X sky130_fd_sc_hd__a31o_1
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5530_ _5594_/A _5531_/B vssd1 vssd1 vccd1 vccd1 _5532_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_26_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5461_ _5459_/X _5460_/X _5567_/B vssd1 vssd1 vccd1 vccd1 _5461_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3807__B _3883_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4412_ _5732_/A _4409_/X _4410_/X _4411_/X vssd1 vssd1 vccd1 vccd1 _4412_/X sky130_fd_sc_hd__o31a_1
XANTENNA__4704__A1 _4713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5392_ _5513_/S _6023_/A _5391_/X _5386_/Y vssd1 vssd1 vccd1 vccd1 _5392_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_1_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4343_ _5398_/A _5362_/A _5603_/C _4271_/X _5624_/A vssd1 vssd1 vccd1 vccd1 _4343_/X
+ sky130_fd_sc_hd__a2111o_1
XANTENNA__4180__A2 _4462_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4274_ _4276_/A _3396_/B _4273_/X _5362_/A _5388_/A vssd1 vssd1 vccd1 vccd1 _4274_/X
+ sky130_fd_sc_hd__a311o_1
X_3225_ _3511_/A _3268_/B vssd1 vssd1 vccd1 vccd1 _3225_/X sky130_fd_sc_hd__or2_1
X_6013_ _4656_/A hold618/X _6019_/S vssd1 vssd1 vccd1 vccd1 _6459_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_94_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3156_ _3323_/A _3168_/B _3229_/A _3205_/B vssd1 vssd1 vccd1 vccd1 _3249_/B sky130_fd_sc_hd__and4b_2
X_3087_ _6349_/Q vssd1 vssd1 vccd1 vccd1 _5117_/A sky130_fd_sc_hd__inv_2
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5196__B2 _6380_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5196__A1 _6379_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3989_ _3773_/Y _5260_/B _3988_/X _6380_/Q vssd1 vssd1 vccd1 vccd1 _3989_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_9_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5728_ _6340_/Q _5628_/X _5629_/X _6482_/Q vssd1 vssd1 vccd1 vccd1 _5737_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_72_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5659_ _4412_/X _5658_/X _5734_/S vssd1 vssd1 vccd1 vccd1 _5659_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_60_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5932__B _5970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold361 _6402_/Q vssd1 vssd1 vccd1 vccd1 hold361/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold350 _4817_/X vssd1 vssd1 vccd1 vccd1 _6317_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold383 _6324_/Q vssd1 vssd1 vccd1 vccd1 hold383/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold372 _4897_/X vssd1 vssd1 vccd1 vccd1 _6321_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold394 _4311_/X vssd1 vssd1 vccd1 vccd1 _6124_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5656__C1 _5730_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout82_A _4408_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3682__A1 _3352_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4503__S _4509_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4698__A0 _6284_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_20_wb_clk_i _6448_/CLK vssd1 vssd1 vccd1 vccd1 _6307_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_3_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3122__B1 _6434_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4961_ _4960_/X _4959_/X _5101_/S vssd1 vssd1 vccd1 vccd1 _4962_/B sky130_fd_sc_hd__mux2_2
X_3912_ _3911_/X hold237/X _4241_/S vssd1 vssd1 vccd1 vccd1 _3912_/X sky130_fd_sc_hd__mux2_1
X_4892_ _6365_/Q _4891_/X _5892_/S vssd1 vssd1 vccd1 vccd1 _4892_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_80_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3843_ _3885_/A _3842_/X _3852_/A vssd1 vssd1 vccd1 vccd1 _3843_/X sky130_fd_sc_hd__o21a_1
XANTENNA__4925__A1 _6367_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3774_ _3774_/A _3774_/B vssd1 vssd1 vccd1 vccd1 _5260_/A sky130_fd_sc_hd__or2_1
XANTENNA__3537__B _5388_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5513_ hold592/X _5512_/X _5513_/S vssd1 vssd1 vccd1 vccd1 _5513_/X sky130_fd_sc_hd__mux2_1
X_5444_ _5432_/A _5431_/B _5429_/X vssd1 vssd1 vccd1 vccd1 _5445_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_100_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4689__B1 _4714_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5375_ _4675_/A _4335_/C _5522_/D _5374_/X vssd1 vssd1 vccd1 vccd1 _5375_/X sky130_fd_sc_hd__a31o_1
XANTENNA__4649__A _5567_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout104 _3390_/X vssd1 vssd1 vccd1 vccd1 _5106_/S sky130_fd_sc_hd__clkbuf_4
Xfanout137 hold638/X vssd1 vssd1 vccd1 vccd1 _4313_/A sky130_fd_sc_hd__clkbuf_8
Xfanout126 _4715_/B2 vssd1 vssd1 vccd1 vccd1 _5393_/A1 sky130_fd_sc_hd__buf_2
X_4326_ _3673_/B _3575_/Y _3590_/Y vssd1 vssd1 vccd1 vccd1 _4326_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_10_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout115 _5489_/S vssd1 vssd1 vccd1 vccd1 _5232_/S sky130_fd_sc_hd__clkbuf_8
Xfanout159 hold611/X vssd1 vssd1 vccd1 vccd1 _4782_/A sky130_fd_sc_hd__buf_4
Xfanout148 _4268_/A vssd1 vssd1 vccd1 vccd1 _3511_/A sky130_fd_sc_hd__buf_4
X_4257_ _5774_/A _3219_/B _5317_/B _4250_/X _4256_/X vssd1 vssd1 vccd1 vccd1 _4257_/X
+ sky130_fd_sc_hd__a311o_1
X_3208_ _3304_/B _4325_/C vssd1 vssd1 vccd1 vccd1 _3590_/A sky130_fd_sc_hd__nor2_2
X_4188_ _6118_/Q _3731_/X _3810_/X _6185_/Q _4187_/X vssd1 vssd1 vccd1 vccd1 _4189_/B
+ sky130_fd_sc_hd__a221o_1
X_3139_ _5124_/A _5315_/A _3326_/B vssd1 vssd1 vccd1 vccd1 _3639_/D sky130_fd_sc_hd__or3_2
XANTENNA__3664__A1 _5757_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5646__C _5734_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3447__B _3619_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold180 _3479_/X vssd1 vssd1 vccd1 vccd1 _6246_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4559__A _5783_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold191 _4489_/X vssd1 vssd1 vccd1 vccd1 _6199_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3407__A1 _5777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3958__A2 _3793_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4907__A1 _6366_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3357__B _4268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_19_wb_clk_i_A _6448_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3490_ _3530_/A _3489_/Y _3471_/B _4800_/S vssd1 vssd1 vccd1 vccd1 _3492_/C sky130_fd_sc_hd__o211a_1
XFILLER_0_59_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3373__A _6442_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5160_ _5160_/A _5160_/B vssd1 vssd1 vccd1 vccd1 _5166_/A sky130_fd_sc_hd__xor2_1
XANTENNA__3804__C _3884_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4111_ _4203_/A _4111_/B vssd1 vssd1 vccd1 vccd1 _5174_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__6366__RESET_B fanout181/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5091_ _6427_/Q _4793_/Y _5083_/X _5090_/X vssd1 vssd1 vccd1 vccd1 _5091_/X sky130_fd_sc_hd__a211o_1
XANTENNA__5635__A2 _5721_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4042_ _4039_/X _4040_/X _4041_/X _4441_/S vssd1 vssd1 vccd1 vccd1 _4042_/X sky130_fd_sc_hd__a22o_2
XANTENNA__4408__S _4408_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5993_ _5995_/C _5995_/B hold551/X _5978_/Y hold472/X vssd1 vssd1 vccd1 vccd1 _5993_/X
+ sky130_fd_sc_hd__a32o_1
X_4944_ _6361_/Q _6362_/Q _6363_/Q _6364_/Q vssd1 vssd1 vccd1 vccd1 _4945_/B sky130_fd_sc_hd__and4_1
XFILLER_0_86_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4875_ _5817_/A _4874_/X _4864_/X vssd1 vssd1 vccd1 vccd1 _4875_/X sky130_fd_sc_hd__a21o_1
XANTENNA_fanout132_A _6430_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3826_ hold97/A hold71/A _3865_/S vssd1 vssd1 vccd1 vccd1 _3826_/X sky130_fd_sc_hd__mux2_1
X_3757_ _6345_/Q _4150_/A _6346_/Q vssd1 vssd1 vccd1 vccd1 _3761_/B sky130_fd_sc_hd__and3b_1
XFILLER_0_40_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3688_ _5296_/A _5296_/B vssd1 vssd1 vccd1 vccd1 _6036_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_30_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6476_ _6481_/CLK _6476_/D fanout176/X vssd1 vssd1 vccd1 vccd1 _6476_/Q sky130_fd_sc_hd__dfstp_1
X_5427_ _6469_/Q _5427_/B vssd1 vssd1 vccd1 vccd1 _5429_/B sky130_fd_sc_hd__nand2_1
XANTENNA__4126__A2 _3804_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5358_ _4281_/B _5368_/S _5357_/X hold585/X _5757_/B vssd1 vssd1 vccd1 vccd1 _6346_/D
+ sky130_fd_sc_hd__a32o_1
X_4309_ _4312_/B _4309_/B vssd1 vssd1 vccd1 vccd1 _4309_/Y sky130_fd_sc_hd__nor2_1
X_5289_ _5288_/X hold572/X _5289_/S vssd1 vssd1 vccd1 vccd1 _5289_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3637__A1 _6457_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3270__C1 _3685_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5566__A2_N _5520_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5314__A1 _4325_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4289__A _4716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3876__A1 _3883_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5865__A2 _6023_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3640__B _6446_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4825__B1 _4963_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4760__A2_N _4720_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output26_A _6529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5567__B _5567_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4660_ input7/X _4668_/B vssd1 vssd1 vccd1 vccd1 _4660_/X sky130_fd_sc_hd__and2_1
XFILLER_0_83_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3611_ _4806_/A _4804_/C _3611_/C vssd1 vssd1 vccd1 vccd1 _4786_/B sky130_fd_sc_hd__nand3_1
XANTENNA__3564__B1 _5777_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4591_ _4675_/A _4276_/X _3514_/B vssd1 vssd1 vccd1 vccd1 _4591_/X sky130_fd_sc_hd__a21o_1
X_6330_ _6407_/CLK _6330_/D fanout170/X vssd1 vssd1 vccd1 vccd1 _6330_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_0_101_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3542_ _5384_/A hold192/X _3540_/Y _3541_/X vssd1 vssd1 vccd1 vccd1 _3542_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_101_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3473_ _5980_/A _4363_/A vssd1 vssd1 vccd1 vccd1 _3473_/X sky130_fd_sc_hd__and2_1
XANTENNA__5305__B2 _5304_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6261_ _6376_/CLK _6261_/D vssd1 vssd1 vccd1 vccd1 _6261_/Q sky130_fd_sc_hd__dfxtp_1
X_5212_ _6461_/Q _6460_/Q vssd1 vssd1 vccd1 vccd1 _5213_/B sky130_fd_sc_hd__xor2_1
X_6192_ _6452_/CLK hold54/X vssd1 vssd1 vccd1 vccd1 hold53/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5143_ _5292_/S _5134_/Y _5142_/X _5119_/Y vssd1 vssd1 vccd1 vccd1 _5143_/X sky130_fd_sc_hd__a31o_1
XANTENNA__5069__A0 _6463_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5074_ _5964_/A _5073_/X _5063_/Y vssd1 vssd1 vccd1 vccd1 _5074_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_79_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4025_ _3979_/A _5256_/B _4023_/X _4024_/X vssd1 vssd1 vccd1 vccd1 _5221_/B sky130_fd_sc_hd__a211o_1
XFILLER_0_79_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4662__A input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5976_ _5975_/X _5970_/Y _5976_/S vssd1 vssd1 vccd1 vccd1 _5976_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_59_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5477__B _6463_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4927_ _6481_/Q _5104_/A2 _4796_/Y _4920_/B _4793_/Y vssd1 vssd1 vccd1 vccd1 _4929_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_51_80 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4858_ _3094_/Y _5771_/A _4856_/Y _4857_/Y _5783_/A vssd1 vssd1 vccd1 vccd1 _4858_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_74_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3809_ _6218_/Q _6003_/A _4400_/A _6134_/Q vssd1 vssd1 vccd1 vccd1 _3809_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_7_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4789_ _5861_/S _4789_/B vssd1 vssd1 vccd1 vccd1 _4789_/Y sky130_fd_sc_hd__nor2_1
X_6528_ _6529_/A vssd1 vssd1 vccd1 vccd1 _6528_/X sky130_fd_sc_hd__buf_1
X_6459_ _6465_/CLK _6459_/D fanout181/X vssd1 vssd1 vccd1 vccd1 _6459_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6101__B _6101_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3741__A _4150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4556__B _5489_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4291__B _5757_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3619__C _3619_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4511__S _4518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5834__C _5866_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5697__S1 _5734_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4274__A1 _4276_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5471__A0 _5605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5223__A0 _6312_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5830_ _5817_/A _5829_/X _4864_/X vssd1 vssd1 vccd1 vccd1 _5830_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_91_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5761_ _6312_/Q hold407/X _5765_/S vssd1 vssd1 vccd1 vccd1 _5761_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_29_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4712_ _6287_/Q _4711_/X _4712_/S vssd1 vssd1 vccd1 vccd1 _4713_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_56_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5692_ _6174_/Q _5721_/A2 _5721_/B1 _6253_/Q _5721_/C1 vssd1 vssd1 vccd1 vccd1 _5693_/B
+ sky130_fd_sc_hd__o221a_1
XANTENNA__4329__A2 _3668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4643_ hold628/X _4606_/X _4607_/X hold629/X _4642_/X vssd1 vssd1 vccd1 vccd1 _4643_/X
+ sky130_fd_sc_hd__a221o_1
X_4574_ hold481/X _6339_/Q _4575_/S vssd1 vssd1 vccd1 vccd1 _4574_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_4_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3525_ _5384_/A _5146_/C vssd1 vssd1 vccd1 vccd1 _3525_/Y sky130_fd_sc_hd__nor2_2
X_6313_ _6417_/CLK _6313_/D fanout174/X vssd1 vssd1 vccd1 vccd1 _6313_/Q sky130_fd_sc_hd__dfstp_4
X_6244_ _6439_/CLK _6244_/D fanout178/X vssd1 vssd1 vccd1 vccd1 _6244_/Q sky130_fd_sc_hd__dfrtp_1
X_3456_ _5371_/B _3456_/B _3456_/C _3456_/D vssd1 vssd1 vccd1 vccd1 _3456_/X sky130_fd_sc_hd__or4_1
XANTENNA__3561__A _5777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5252__S _5292_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3387_ _4802_/A _4802_/B _3386_/Y vssd1 vssd1 vccd1 vccd1 _3387_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_41_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6175_ _6454_/CLK _6175_/D vssd1 vssd1 vccd1 vccd1 _6175_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5126_ _4716_/A _6333_/Q _5244_/S vssd1 vssd1 vccd1 vccd1 _5126_/Y sky130_fd_sc_hd__a21oi_1
X_5057_ _5056_/X hold411/X _5098_/S vssd1 vssd1 vccd1 vccd1 _5057_/X sky130_fd_sc_hd__mux2_1
X_4008_ _4007_/A _4007_/B _4156_/A vssd1 vssd1 vccd1 vccd1 _4008_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__4265__A1 _5605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5462__A0 _6461_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4017__A1 _6334_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5959_ _5959_/A _5959_/B vssd1 vssd1 vccd1 vccd1 _5961_/A sky130_fd_sc_hd__or2_1
XANTENNA__5765__A1 hold572/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3736__A _5600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3471__A _4800_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold40 hold40/A vssd1 vssd1 vccd1 vccd1 hold40/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 hold73/A vssd1 vssd1 vccd1 vccd1 hold73/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 hold62/A vssd1 vssd1 vccd1 vccd1 hold62/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 hold51/A vssd1 vssd1 vccd1 vccd1 hold51/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4256__A1 _5388_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold84 hold84/A vssd1 vssd1 vccd1 vccd1 hold84/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 hold95/A vssd1 vssd1 vccd1 vccd1 hold95/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5398__A _5398_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_45_wb_clk_i clkbuf_leaf_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6400_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__4506__S _4509_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4730__A1_N _6310_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3519__B1 _5384_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4241__S _4241_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_4 _5697_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3310_ _3310_/A _3608_/A _4785_/A _3394_/A vssd1 vssd1 vccd1 vccd1 _3310_/Y sky130_fd_sc_hd__nor4_1
XFILLER_0_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4290_ _5124_/A _5478_/S _4768_/S vssd1 vssd1 vccd1 vccd1 _4322_/B sky130_fd_sc_hd__and3_2
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3241_ _3240_/B _3174_/B _3986_/A _5387_/A vssd1 vssd1 vccd1 vccd1 _3241_/X sky130_fd_sc_hd__a211o_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3172_ _3172_/A _3547_/B vssd1 vssd1 vccd1 vccd1 _3172_/Y sky130_fd_sc_hd__nand2_1
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5692__B1 _5721_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5813_ _5813_/A _5813_/B _5811_/X vssd1 vssd1 vccd1 vccd1 _5814_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_57_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5744_ hold33/X _3859_/B _5769_/S vssd1 vssd1 vccd1 vccd1 hold34/A sky130_fd_sc_hd__mux2_1
X_5675_ _5757_/B hold554/X _5611_/Y _5674_/X vssd1 vssd1 vccd1 vccd1 _5675_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_32_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4626_ _3847_/B _4052_/B _4641_/B vssd1 vssd1 vccd1 vccd1 _4626_/X sky130_fd_sc_hd__mux2_1
Xhold510 _6278_/Q vssd1 vssd1 vccd1 vccd1 hold510/X sky130_fd_sc_hd__dlygate4sd3_1
X_4557_ _5322_/A _5387_/A _4557_/C _4557_/D vssd1 vssd1 vccd1 vccd1 wire92/A sky130_fd_sc_hd__nor4_1
Xhold543 _6473_/Q vssd1 vssd1 vccd1 vccd1 _3640_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold554 _6380_/Q vssd1 vssd1 vccd1 vccd1 hold554/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5771__A _5771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold532 _5591_/X vssd1 vssd1 vccd1 vccd1 _6375_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold521 _6082_/X vssd1 vssd1 vccd1 vccd1 _6484_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold565 _4615_/X vssd1 vssd1 vccd1 vccd1 _6285_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3508_ _5400_/A _3638_/B vssd1 vssd1 vccd1 vccd1 _5398_/B sky130_fd_sc_hd__nor2_1
Xhold576 _3510_/X vssd1 vssd1 vccd1 vccd1 _6159_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold587 _5921_/X vssd1 vssd1 vccd1 vccd1 _6423_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4488_ _4085_/X hold213/X _4491_/S vssd1 vssd1 vccd1 vccd1 _6198_/D sky130_fd_sc_hd__mux2_1
X_3439_ _5309_/A _3406_/Y _3415_/X _3456_/B vssd1 vssd1 vccd1 vccd1 _3440_/C sky130_fd_sc_hd__a211o_1
Xhold598 _6338_/Q vssd1 vssd1 vccd1 vccd1 hold598/X sky130_fd_sc_hd__dlygate4sd3_1
X_6227_ _6452_/CLK _6227_/D vssd1 vssd1 vccd1 vccd1 _6227_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5490__B _6464_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6158_ _6488_/CLK _6158_/D vssd1 vssd1 vccd1 vccd1 _6158_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5109_ _5109_/A1 _5106_/X _5108_/X _4924_/C vssd1 vssd1 vccd1 vccd1 _5109_/X sky130_fd_sc_hd__a22o_1
X_6089_ _6089_/A _6107_/S vssd1 vssd1 vccd1 vccd1 _6089_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__4238__A1 _5730_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5986__A1 _5995_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5738__A1 _5757_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4946__C1 _4924_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5157__S _5289_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3466__A _6021_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4996__S _5974_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput52 _3659_/X vssd1 vssd1 vccd1 vccd1 io_out[34] sky130_fd_sc_hd__buf_12
Xoutput41 _6305_/Q vssd1 vssd1 vccd1 vccd1 io_out[22] sky130_fd_sc_hd__buf_12
Xoutput30 _6323_/Q vssd1 vssd1 vccd1 vccd1 io_out[12] sky130_fd_sc_hd__buf_12
XANTENNA__3913__B _4150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5278__D _6464_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5729__A1 _6316_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3790_ _4675_/A _5317_/B _3665_/A vssd1 vssd1 vccd1 vccd1 _3790_/X sky130_fd_sc_hd__a21o_1
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5460_ hold607/X input7/X _5510_/S vssd1 vssd1 vccd1 vccd1 _5460_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_54_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3807__C _3884_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4411_ _5730_/C1 _4408_/X _4407_/X _5655_/B vssd1 vssd1 vccd1 vccd1 _4411_/X sky130_fd_sc_hd__a211o_1
X_5391_ _5391_/A _5391_/B _5391_/C _5377_/Y vssd1 vssd1 vccd1 vccd1 _5391_/X sky130_fd_sc_hd__or4b_1
XFILLER_0_22_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4342_ _4324_/A _4341_/Y _4324_/X _4782_/A vssd1 vssd1 vccd1 vccd1 _5644_/A sky130_fd_sc_hd__a2bb2o_4
XANTENNA__6487__SET_B fanout176/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4273_ _4273_/A _4273_/B vssd1 vssd1 vccd1 vccd1 _4273_/X sky130_fd_sc_hd__and2_1
X_3224_ _6299_/Q _6300_/Q _3986_/A vssd1 vssd1 vccd1 vccd1 _3268_/B sky130_fd_sc_hd__nand3b_4
X_6012_ _4650_/A hold616/X _6019_/S vssd1 vssd1 vccd1 vccd1 _6458_/D sky130_fd_sc_hd__mux2_1
.ends

