magic
tech sky130B
magscale 1 2
timestamp 1717329487
<< obsli1 >>
rect 1104 2159 43884 42449
<< obsm1 >>
rect 934 2128 43884 42480
<< metal2 >>
rect 1490 44200 1546 45000
rect 2686 44200 2742 45000
rect 3882 44200 3938 45000
rect 5078 44200 5134 45000
rect 6274 44200 6330 45000
rect 7470 44200 7526 45000
rect 8666 44200 8722 45000
rect 9862 44200 9918 45000
rect 11058 44200 11114 45000
rect 12254 44200 12310 45000
rect 13450 44200 13506 45000
rect 14646 44200 14702 45000
rect 15842 44200 15898 45000
rect 17038 44200 17094 45000
rect 18234 44200 18290 45000
rect 19430 44200 19486 45000
rect 20626 44200 20682 45000
rect 21822 44200 21878 45000
rect 23018 44200 23074 45000
rect 24214 44200 24270 45000
rect 25410 44200 25466 45000
rect 26606 44200 26662 45000
rect 27802 44200 27858 45000
rect 28998 44200 29054 45000
rect 30194 44200 30250 45000
rect 31390 44200 31446 45000
rect 32586 44200 32642 45000
rect 33782 44200 33838 45000
rect 34978 44200 35034 45000
rect 36174 44200 36230 45000
rect 37370 44200 37426 45000
rect 38566 44200 38622 45000
rect 39762 44200 39818 45000
rect 40958 44200 41014 45000
rect 42154 44200 42210 45000
rect 43350 44200 43406 45000
rect 22466 0 22522 800
<< obsm2 >>
rect 938 44144 1434 44200
rect 1602 44144 2630 44200
rect 2798 44144 3826 44200
rect 3994 44144 5022 44200
rect 5190 44144 6218 44200
rect 6386 44144 7414 44200
rect 7582 44144 8610 44200
rect 8778 44144 9806 44200
rect 9974 44144 11002 44200
rect 11170 44144 12198 44200
rect 12366 44144 13394 44200
rect 13562 44144 14590 44200
rect 14758 44144 15786 44200
rect 15954 44144 16982 44200
rect 17150 44144 18178 44200
rect 18346 44144 19374 44200
rect 19542 44144 20570 44200
rect 20738 44144 21766 44200
rect 21934 44144 22962 44200
rect 23130 44144 24158 44200
rect 24326 44144 25354 44200
rect 25522 44144 26550 44200
rect 26718 44144 27746 44200
rect 27914 44144 28942 44200
rect 29110 44144 30138 44200
rect 30306 44144 31334 44200
rect 31502 44144 32530 44200
rect 32698 44144 33726 44200
rect 33894 44144 34922 44200
rect 35090 44144 36118 44200
rect 36286 44144 37314 44200
rect 37482 44144 38510 44200
rect 38678 44144 39706 44200
rect 39874 44144 40902 44200
rect 41070 44144 42098 44200
rect 42266 44144 43294 44200
rect 43462 44144 43866 44200
rect 938 856 43866 44144
rect 938 800 22410 856
rect 22578 800 43866 856
<< metal3 >>
rect 0 41352 800 41472
rect 0 40264 800 40384
rect 0 39176 800 39296
rect 44200 39176 45000 39296
rect 0 38088 800 38208
rect 0 37000 800 37120
rect 0 35912 800 36032
rect 0 34824 800 34944
rect 0 33736 800 33856
rect 0 32648 800 32768
rect 0 31560 800 31680
rect 0 30472 800 30592
rect 0 29384 800 29504
rect 0 28296 800 28416
rect 44200 28024 45000 28144
rect 0 27208 800 27328
rect 0 26120 800 26240
rect 0 25032 800 25152
rect 0 23944 800 24064
rect 0 22856 800 22976
rect 0 21768 800 21888
rect 0 20680 800 20800
rect 0 19592 800 19712
rect 0 18504 800 18624
rect 0 17416 800 17536
rect 44200 16872 45000 16992
rect 0 16328 800 16448
rect 0 15240 800 15360
rect 0 14152 800 14272
rect 0 13064 800 13184
rect 0 11976 800 12096
rect 0 10888 800 11008
rect 0 9800 800 9920
rect 0 8712 800 8832
rect 0 7624 800 7744
rect 0 6536 800 6656
rect 44200 5720 45000 5840
rect 0 5448 800 5568
rect 0 4360 800 4480
rect 0 3272 800 3392
<< obsm3 >>
rect 800 41552 44200 42465
rect 880 41272 44200 41552
rect 800 40464 44200 41272
rect 880 40184 44200 40464
rect 800 39376 44200 40184
rect 880 39096 44120 39376
rect 800 38288 44200 39096
rect 880 38008 44200 38288
rect 800 37200 44200 38008
rect 880 36920 44200 37200
rect 800 36112 44200 36920
rect 880 35832 44200 36112
rect 800 35024 44200 35832
rect 880 34744 44200 35024
rect 800 33936 44200 34744
rect 880 33656 44200 33936
rect 800 32848 44200 33656
rect 880 32568 44200 32848
rect 800 31760 44200 32568
rect 880 31480 44200 31760
rect 800 30672 44200 31480
rect 880 30392 44200 30672
rect 800 29584 44200 30392
rect 880 29304 44200 29584
rect 800 28496 44200 29304
rect 880 28224 44200 28496
rect 880 28216 44120 28224
rect 800 27944 44120 28216
rect 800 27408 44200 27944
rect 880 27128 44200 27408
rect 800 26320 44200 27128
rect 880 26040 44200 26320
rect 800 25232 44200 26040
rect 880 24952 44200 25232
rect 800 24144 44200 24952
rect 880 23864 44200 24144
rect 800 23056 44200 23864
rect 880 22776 44200 23056
rect 800 21968 44200 22776
rect 880 21688 44200 21968
rect 800 20880 44200 21688
rect 880 20600 44200 20880
rect 800 19792 44200 20600
rect 880 19512 44200 19792
rect 800 18704 44200 19512
rect 880 18424 44200 18704
rect 800 17616 44200 18424
rect 880 17336 44200 17616
rect 800 17072 44200 17336
rect 800 16792 44120 17072
rect 800 16528 44200 16792
rect 880 16248 44200 16528
rect 800 15440 44200 16248
rect 880 15160 44200 15440
rect 800 14352 44200 15160
rect 880 14072 44200 14352
rect 800 13264 44200 14072
rect 880 12984 44200 13264
rect 800 12176 44200 12984
rect 880 11896 44200 12176
rect 800 11088 44200 11896
rect 880 10808 44200 11088
rect 800 10000 44200 10808
rect 880 9720 44200 10000
rect 800 8912 44200 9720
rect 880 8632 44200 8912
rect 800 7824 44200 8632
rect 880 7544 44200 7824
rect 800 6736 44200 7544
rect 880 6456 44200 6736
rect 800 5920 44200 6456
rect 800 5648 44120 5920
rect 880 5640 44120 5648
rect 880 5368 44200 5640
rect 800 4560 44200 5368
rect 880 4280 44200 4560
rect 800 3472 44200 4280
rect 880 3192 44200 3472
rect 800 2143 44200 3192
<< metal4 >>
rect 4208 2128 4528 42480
rect 19568 2128 19888 42480
rect 34928 2128 35248 42480
<< obsm4 >>
rect 3187 2619 4128 38453
rect 4608 2619 19488 38453
rect 19968 2619 28645 38453
<< labels >>
rlabel metal3 s 44200 28024 45000 28144 6 custom_settings[0]
port 1 nsew signal input
rlabel metal3 s 44200 39176 45000 39296 6 custom_settings[1]
port 2 nsew signal input
rlabel metal2 s 1490 44200 1546 45000 6 io_in[0]
port 3 nsew signal input
rlabel metal2 s 13450 44200 13506 45000 6 io_in[10]
port 4 nsew signal input
rlabel metal2 s 14646 44200 14702 45000 6 io_in[11]
port 5 nsew signal input
rlabel metal2 s 15842 44200 15898 45000 6 io_in[12]
port 6 nsew signal input
rlabel metal2 s 17038 44200 17094 45000 6 io_in[13]
port 7 nsew signal input
rlabel metal2 s 18234 44200 18290 45000 6 io_in[14]
port 8 nsew signal input
rlabel metal2 s 19430 44200 19486 45000 6 io_in[15]
port 9 nsew signal input
rlabel metal2 s 20626 44200 20682 45000 6 io_in[16]
port 10 nsew signal input
rlabel metal2 s 21822 44200 21878 45000 6 io_in[17]
port 11 nsew signal input
rlabel metal2 s 23018 44200 23074 45000 6 io_in[18]
port 12 nsew signal input
rlabel metal2 s 24214 44200 24270 45000 6 io_in[19]
port 13 nsew signal input
rlabel metal2 s 2686 44200 2742 45000 6 io_in[1]
port 14 nsew signal input
rlabel metal2 s 25410 44200 25466 45000 6 io_in[20]
port 15 nsew signal input
rlabel metal2 s 26606 44200 26662 45000 6 io_in[21]
port 16 nsew signal input
rlabel metal2 s 27802 44200 27858 45000 6 io_in[22]
port 17 nsew signal input
rlabel metal2 s 28998 44200 29054 45000 6 io_in[23]
port 18 nsew signal input
rlabel metal2 s 30194 44200 30250 45000 6 io_in[24]
port 19 nsew signal input
rlabel metal2 s 31390 44200 31446 45000 6 io_in[25]
port 20 nsew signal input
rlabel metal2 s 32586 44200 32642 45000 6 io_in[26]
port 21 nsew signal input
rlabel metal2 s 33782 44200 33838 45000 6 io_in[27]
port 22 nsew signal input
rlabel metal2 s 34978 44200 35034 45000 6 io_in[28]
port 23 nsew signal input
rlabel metal2 s 36174 44200 36230 45000 6 io_in[29]
port 24 nsew signal input
rlabel metal2 s 3882 44200 3938 45000 6 io_in[2]
port 25 nsew signal input
rlabel metal2 s 37370 44200 37426 45000 6 io_in[30]
port 26 nsew signal input
rlabel metal2 s 38566 44200 38622 45000 6 io_in[31]
port 27 nsew signal input
rlabel metal2 s 39762 44200 39818 45000 6 io_in[32]
port 28 nsew signal input
rlabel metal2 s 40958 44200 41014 45000 6 io_in[33]
port 29 nsew signal input
rlabel metal2 s 42154 44200 42210 45000 6 io_in[34]
port 30 nsew signal input
rlabel metal2 s 43350 44200 43406 45000 6 io_in[35]
port 31 nsew signal input
rlabel metal2 s 5078 44200 5134 45000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 6274 44200 6330 45000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 7470 44200 7526 45000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 8666 44200 8722 45000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 9862 44200 9918 45000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 11058 44200 11114 45000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 12254 44200 12310 45000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 22466 0 22522 800 6 io_oeb
port 39 nsew signal output
rlabel metal3 s 0 3272 800 3392 6 io_out[0]
port 40 nsew signal output
rlabel metal3 s 0 14152 800 14272 6 io_out[10]
port 41 nsew signal output
rlabel metal3 s 0 15240 800 15360 6 io_out[11]
port 42 nsew signal output
rlabel metal3 s 0 16328 800 16448 6 io_out[12]
port 43 nsew signal output
rlabel metal3 s 0 17416 800 17536 6 io_out[13]
port 44 nsew signal output
rlabel metal3 s 0 18504 800 18624 6 io_out[14]
port 45 nsew signal output
rlabel metal3 s 0 19592 800 19712 6 io_out[15]
port 46 nsew signal output
rlabel metal3 s 0 20680 800 20800 6 io_out[16]
port 47 nsew signal output
rlabel metal3 s 0 21768 800 21888 6 io_out[17]
port 48 nsew signal output
rlabel metal3 s 0 22856 800 22976 6 io_out[18]
port 49 nsew signal output
rlabel metal3 s 0 23944 800 24064 6 io_out[19]
port 50 nsew signal output
rlabel metal3 s 0 4360 800 4480 6 io_out[1]
port 51 nsew signal output
rlabel metal3 s 0 25032 800 25152 6 io_out[20]
port 52 nsew signal output
rlabel metal3 s 0 26120 800 26240 6 io_out[21]
port 53 nsew signal output
rlabel metal3 s 0 27208 800 27328 6 io_out[22]
port 54 nsew signal output
rlabel metal3 s 0 28296 800 28416 6 io_out[23]
port 55 nsew signal output
rlabel metal3 s 0 29384 800 29504 6 io_out[24]
port 56 nsew signal output
rlabel metal3 s 0 30472 800 30592 6 io_out[25]
port 57 nsew signal output
rlabel metal3 s 0 31560 800 31680 6 io_out[26]
port 58 nsew signal output
rlabel metal3 s 0 32648 800 32768 6 io_out[27]
port 59 nsew signal output
rlabel metal3 s 0 33736 800 33856 6 io_out[28]
port 60 nsew signal output
rlabel metal3 s 0 34824 800 34944 6 io_out[29]
port 61 nsew signal output
rlabel metal3 s 0 5448 800 5568 6 io_out[2]
port 62 nsew signal output
rlabel metal3 s 0 35912 800 36032 6 io_out[30]
port 63 nsew signal output
rlabel metal3 s 0 37000 800 37120 6 io_out[31]
port 64 nsew signal output
rlabel metal3 s 0 38088 800 38208 6 io_out[32]
port 65 nsew signal output
rlabel metal3 s 0 39176 800 39296 6 io_out[33]
port 66 nsew signal output
rlabel metal3 s 0 40264 800 40384 6 io_out[34]
port 67 nsew signal output
rlabel metal3 s 0 41352 800 41472 6 io_out[35]
port 68 nsew signal output
rlabel metal3 s 0 6536 800 6656 6 io_out[3]
port 69 nsew signal output
rlabel metal3 s 0 7624 800 7744 6 io_out[4]
port 70 nsew signal output
rlabel metal3 s 0 8712 800 8832 6 io_out[5]
port 71 nsew signal output
rlabel metal3 s 0 9800 800 9920 6 io_out[6]
port 72 nsew signal output
rlabel metal3 s 0 10888 800 11008 6 io_out[7]
port 73 nsew signal output
rlabel metal3 s 0 11976 800 12096 6 io_out[8]
port 74 nsew signal output
rlabel metal3 s 0 13064 800 13184 6 io_out[9]
port 75 nsew signal output
rlabel metal3 s 44200 16872 45000 16992 6 rst_n
port 76 nsew signal input
rlabel metal4 s 4208 2128 4528 42480 6 vccd1
port 77 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 42480 6 vccd1
port 77 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 42480 6 vssd1
port 78 nsew ground bidirectional
rlabel metal3 s 44200 5720 45000 5840 6 wb_clk_i
port 79 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 45000 45000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 5535944
string GDS_FILE /home/tholin/Desktop/ci2406-rej-pommedeterrible-tholin/openlane/MOS6502/runs/24_06_02_13_45/results/signoff/wrapped_6502.magic.gds
string GDS_START 922100
<< end >>

