* NGSPICE file created from execution_unit.ext - technology: sky130B

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_4 abstract view
.subckt sky130_fd_sc_hd__o41a_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_4 abstract view
.subckt sky130_fd_sc_hd__o311a_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_2 abstract view
.subckt sky130_fd_sc_hd__a2111oi_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_2 abstract view
.subckt sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_4 abstract view
.subckt sky130_fd_sc_hd__o311ai_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_4 abstract view
.subckt sky130_fd_sc_hd__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_2 abstract view
.subckt sky130_fd_sc_hd__o2111a_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_4 abstract view
.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_4 abstract view
.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_4 abstract view
.subckt sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_4 abstract view
.subckt sky130_fd_sc_hd__a311o_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_4 abstract view
.subckt sky130_fd_sc_hd__a21bo_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

.subckt execution_unit busy curr_PC[0] curr_PC[10] curr_PC[11] curr_PC[12] curr_PC[13]
+ curr_PC[14] curr_PC[15] curr_PC[16] curr_PC[17] curr_PC[18] curr_PC[19] curr_PC[1]
+ curr_PC[20] curr_PC[21] curr_PC[22] curr_PC[23] curr_PC[24] curr_PC[25] curr_PC[26]
+ curr_PC[27] curr_PC[2] curr_PC[3] curr_PC[4] curr_PC[5] curr_PC[6] curr_PC[7] curr_PC[8]
+ curr_PC[9] dest_idx[0] dest_idx[1] dest_idx[2] dest_idx[3] dest_idx[4] dest_mask[0]
+ dest_mask[1] dest_pred[0] dest_pred[1] dest_pred[2] dest_pred_val dest_val[0] dest_val[10]
+ dest_val[11] dest_val[12] dest_val[13] dest_val[14] dest_val[15] dest_val[16] dest_val[17]
+ dest_val[18] dest_val[19] dest_val[1] dest_val[20] dest_val[21] dest_val[22] dest_val[23]
+ dest_val[24] dest_val[25] dest_val[26] dest_val[27] dest_val[28] dest_val[29] dest_val[2]
+ dest_val[30] dest_val[31] dest_val[3] dest_val[4] dest_val[5] dest_val[6] dest_val[7]
+ dest_val[8] dest_val[9] instruction[0] instruction[10] instruction[11] instruction[12]
+ instruction[13] instruction[14] instruction[15] instruction[16] instruction[17]
+ instruction[18] instruction[19] instruction[1] instruction[20] instruction[21] instruction[22]
+ instruction[23] instruction[24] instruction[25] instruction[26] instruction[27]
+ instruction[28] instruction[29] instruction[2] instruction[30] instruction[31] instruction[32]
+ instruction[33] instruction[34] instruction[35] instruction[36] instruction[37]
+ instruction[38] instruction[39] instruction[3] instruction[40] instruction[41] instruction[4]
+ instruction[5] instruction[6] instruction[7] instruction[8] instruction[9] is_load
+ is_store loadstore_address[0] loadstore_address[10] loadstore_address[11] loadstore_address[12]
+ loadstore_address[13] loadstore_address[14] loadstore_address[15] loadstore_address[16]
+ loadstore_address[17] loadstore_address[18] loadstore_address[19] loadstore_address[1]
+ loadstore_address[20] loadstore_address[21] loadstore_address[22] loadstore_address[23]
+ loadstore_address[24] loadstore_address[25] loadstore_address[26] loadstore_address[27]
+ loadstore_address[28] loadstore_address[29] loadstore_address[2] loadstore_address[30]
+ loadstore_address[31] loadstore_address[3] loadstore_address[4] loadstore_address[5]
+ loadstore_address[6] loadstore_address[7] loadstore_address[8] loadstore_address[9]
+ loadstore_dest[0] loadstore_dest[1] loadstore_dest[2] loadstore_dest[3] loadstore_dest[4]
+ loadstore_size[0] loadstore_size[1] new_PC[0] new_PC[10] new_PC[11] new_PC[12] new_PC[13]
+ new_PC[14] new_PC[15] new_PC[16] new_PC[17] new_PC[18] new_PC[19] new_PC[1] new_PC[20]
+ new_PC[21] new_PC[22] new_PC[23] new_PC[24] new_PC[25] new_PC[26] new_PC[27] new_PC[2]
+ new_PC[3] new_PC[4] new_PC[5] new_PC[6] new_PC[7] new_PC[8] new_PC[9] pred_idx[0]
+ pred_idx[1] pred_idx[2] pred_val reg1_idx[0] reg1_idx[1] reg1_idx[2] reg1_idx[3]
+ reg1_idx[4] reg1_val[0] reg1_val[10] reg1_val[11] reg1_val[12] reg1_val[13] reg1_val[14]
+ reg1_val[15] reg1_val[16] reg1_val[17] reg1_val[18] reg1_val[19] reg1_val[1] reg1_val[20]
+ reg1_val[21] reg1_val[22] reg1_val[23] reg1_val[24] reg1_val[25] reg1_val[26] reg1_val[27]
+ reg1_val[28] reg1_val[29] reg1_val[2] reg1_val[30] reg1_val[31] reg1_val[3] reg1_val[4]
+ reg1_val[5] reg1_val[6] reg1_val[7] reg1_val[8] reg1_val[9] reg2_idx[0] reg2_idx[1]
+ reg2_idx[2] reg2_idx[3] reg2_idx[4] reg2_val[0] reg2_val[10] reg2_val[11] reg2_val[12]
+ reg2_val[13] reg2_val[14] reg2_val[15] reg2_val[16] reg2_val[17] reg2_val[18] reg2_val[19]
+ reg2_val[1] reg2_val[20] reg2_val[21] reg2_val[22] reg2_val[23] reg2_val[24] reg2_val[25]
+ reg2_val[26] reg2_val[27] reg2_val[28] reg2_val[29] reg2_val[2] reg2_val[30] reg2_val[31]
+ reg2_val[3] reg2_val[4] reg2_val[5] reg2_val[6] reg2_val[7] reg2_val[8] reg2_val[9]
+ rst sign_extend take_branch vccd1 vssd1 wb_clk_i
XFILLER_0_94_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06883_ instruction[1] instruction[2] instruction[0] pred_val vssd1 vssd1 vccd1 vccd1
+ _06921_/B sky130_fd_sc_hd__and4b_4
X_09671_ _09668_/X _09670_/X _11010_/S vssd1 vssd1 vccd1 vccd1 _09671_/X sky130_fd_sc_hd__mux2_1
X_08622_ _08621_/A _08622_/B vssd1 vssd1 vccd1 vccd1 _08625_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_27_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12815__C1 _13128_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08553_ _08681_/A _08553_/B vssd1 vssd1 vccd1 vccd1 _08558_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_76_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08484_ _08493_/A _08493_/B vssd1 vssd1 vccd1 vccd1 _08485_/B sky130_fd_sc_hd__nand2b_1
X_07504_ instruction[7] _07503_/X reg1_val[31] vssd1 vssd1 vccd1 vccd1 _07504_/Y sky130_fd_sc_hd__a21boi_4
XFILLER_0_49_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07435_ _12838_/A _10167_/A1 _10022_/B1 _12840_/A vssd1 vssd1 vccd1 vccd1 _07436_/B
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_64_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_339 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07366_ _09548_/A _07508_/B vssd1 vssd1 vccd1 vccd1 _07366_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_45_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09105_ _09103_/X _09104_/X _09330_/S vssd1 vssd1 vccd1 vccd1 _09105_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_60_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07297_ _11472_/A _10167_/A1 _10022_/B1 _11558_/A vssd1 vssd1 vccd1 vccd1 _07298_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_33_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08798__B1 _08752_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09036_ _09036_/A _09036_/B vssd1 vssd1 vccd1 vccd1 _09036_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_60_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09938_ _09939_/A _09939_/B vssd1 vssd1 vccd1 vccd1 _09938_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__07773__A1 _07955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07773__B2 _07896_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09869_ _09869_/A _09869_/B _09869_/C vssd1 vssd1 vccd1 vccd1 _09870_/B sky130_fd_sc_hd__or3_1
X_12880_ hold277/X hold47/X vssd1 vssd1 vccd1 vccd1 _13174_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__08619__A _08733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11900_ _12290_/A _11872_/X _11873_/Y _11876_/Y _11899_/X vssd1 vssd1 vccd1 vccd1
+ _11900_/X sky130_fd_sc_hd__o311a_1
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09278__A1 _09351_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11831_ _11830_/B _11831_/B vssd1 vssd1 vccd1 vccd1 _11832_/B sky130_fd_sc_hd__and2b_1
XTAP_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12821__A2 _12818_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07828__A2 _07087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11762_ _11761_/B _11762_/B vssd1 vssd1 vccd1 vccd1 _11763_/B sky130_fd_sc_hd__and2b_1
XTAP_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10713_ _10554_/Y _10557_/B _10562_/A vssd1 vssd1 vccd1 vccd1 _10714_/B sky130_fd_sc_hd__a21o_1
X_11693_ _11693_/A _11693_/B _11693_/C vssd1 vssd1 vccd1 vccd1 _11694_/B sky130_fd_sc_hd__nand3_1
X_10644_ _09527_/B _09354_/B _10644_/S vssd1 vssd1 vccd1 vccd1 _10644_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_70_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13363_ _13384_/CLK _13363_/D vssd1 vssd1 vccd1 vccd1 hold292/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10575_ _10575_/A _10575_/B vssd1 vssd1 vccd1 vccd1 _10576_/C sky130_fd_sc_hd__or2_1
XANTENNA__07461__B1 _10571_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12314_ fanout9/X fanout8/X fanout4/X fanout12/X vssd1 vssd1 vccd1 vccd1 _12315_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13294_ _13307_/CLK _13294_/D vssd1 vssd1 vccd1 vccd1 hold189/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12245_ hold281/A _12245_/B vssd1 vssd1 vccd1 vccd1 _12301_/B sky130_fd_sc_hd__or2_1
XANTENNA__10899__A1 _07074_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12176_ _12176_/A _12176_/B vssd1 vssd1 vccd1 vccd1 _12176_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__09753__A2 _11558_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11127_ hold212/A _11127_/B vssd1 vssd1 vccd1 vccd1 _11236_/B sky130_fd_sc_hd__or2_1
XANTENNA__06959__D _09351_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11058_ _11261_/A _11058_/B vssd1 vssd1 vccd1 vccd1 _11059_/B sky130_fd_sc_hd__xnor2_1
X_10009_ _10448_/A _10009_/B vssd1 vssd1 vccd1 vccd1 _10010_/A sky130_fd_sc_hd__xor2_1
XANTENNA__09124__S _09142_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13065__A2 _13087_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07220_ _07220_/A _07220_/B _07220_/C vssd1 vssd1 vccd1 vccd1 _08038_/C sky130_fd_sc_hd__and3_2
XFILLER_0_73_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08264__A _08731_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07151_ _07343_/B _07151_/B vssd1 vssd1 vccd1 vccd1 _12264_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_42_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11379__A2 _11989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09992__A2 _09172_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07082_ reg1_val[18] _07254_/B _06997_/C _07364_/B1 vssd1 vssd1 vccd1 vccd1 _07083_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_30_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10051__A2 _10574_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09807__B _09808_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09744__A2 _07099_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07608__A _11261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout138 _12812_/A vssd1 vssd1 vccd1 vccd1 _08739_/A1 sky130_fd_sc_hd__buf_6
Xfanout127 _10022_/B1 vssd1 vssd1 vccd1 vccd1 _08564_/B sky130_fd_sc_hd__clkbuf_8
Xfanout116 _06986_/Y vssd1 vssd1 vccd1 vccd1 _08304_/B sky130_fd_sc_hd__buf_8
Xfanout105 _11987_/A vssd1 vssd1 vccd1 vccd1 _11180_/A sky130_fd_sc_hd__buf_8
X_07984_ _07984_/A _07984_/B vssd1 vssd1 vccd1 vccd1 _07986_/C sky130_fd_sc_hd__and2_1
XFILLER_0_38_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10034__A _12810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout149 _08724_/A vssd1 vssd1 vccd1 vccd1 _11163_/A sky130_fd_sc_hd__clkbuf_16
X_06935_ _12455_/S _06935_/B vssd1 vssd1 vccd1 vccd1 dest_mask[1] sky130_fd_sc_hd__nand2_8
X_09723_ _09564_/A _09564_/B _09565_/X vssd1 vssd1 vccd1 vccd1 _09724_/B sky130_fd_sc_hd__a21oi_2
XANTENNA__07046__C _11987_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06866_ _06866_/A _06866_/B _11437_/A vssd1 vssd1 vccd1 vccd1 _06873_/B sky130_fd_sc_hd__or3b_1
X_09654_ _09653_/A _09853_/A _09853_/B vssd1 vssd1 vccd1 vccd1 _09655_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_97_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08439__A _08681_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08605_ _08606_/A _08605_/B _08605_/C vssd1 vssd1 vccd1 vccd1 _08615_/A sky130_fd_sc_hd__nand3_1
XANTENNA__08180__B2 _12820_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08180__A1 _12818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06797_ reg1_val[2] _10250_/S vssd1 vssd1 vccd1 vccd1 _06798_/B sky130_fd_sc_hd__nand2_1
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09585_ fanout75/X _11751_/A _11766_/A _08304_/B vssd1 vssd1 vccd1 vccd1 _09586_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12803__A2 _12818_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08536_ _08745_/A _08536_/B vssd1 vssd1 vccd1 vccd1 _08573_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_65_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08467_ _08467_/A _08467_/B vssd1 vssd1 vccd1 vccd1 _08495_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_65_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07418_ _06612_/B _07142_/Y _07343_/Y instruction[7] vssd1 vssd1 vccd1 vccd1 _07420_/B
+ sky130_fd_sc_hd__o31a_1
X_08398_ _08394_/X _08398_/B vssd1 vssd1 vccd1 vccd1 _08447_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_52_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07349_ _07349_/A _07349_/B vssd1 vssd1 vccd1 vccd1 _07350_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_80_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08174__A _08728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09432__A1 _12848_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09432__B2 _10941_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10360_ _10360_/A _10360_/B vssd1 vssd1 vccd1 vccd1 _10361_/B sky130_fd_sc_hd__xor2_4
X_09019_ _09014_/Y _09018_/Y _08491_/B vssd1 vssd1 vccd1 vccd1 _09021_/B sky130_fd_sc_hd__a21o_1
X_10291_ _10292_/A _10292_/B _10292_/C vssd1 vssd1 vccd1 vccd1 _10293_/A sky130_fd_sc_hd__o21ai_1
Xhold170 hold170/A vssd1 vssd1 vccd1 vccd1 hold170/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09196__B1 _12812_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12030_ _12170_/A _12030_/B _12030_/C vssd1 vssd1 vccd1 vccd1 _12030_/Y sky130_fd_sc_hd__nand3_1
Xhold192 hold192/A vssd1 vssd1 vccd1 vccd1 hold192/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold181 hold181/A vssd1 vssd1 vccd1 vccd1 hold181/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11542__A2 _11343_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12932_ _13159_/B _13160_/A _12885_/X vssd1 vssd1 vccd1 vccd1 _13165_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_88_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12863_ hold140/X hold256/X vssd1 vssd1 vccd1 vccd1 _12863_/X sky130_fd_sc_hd__and2b_1
XANTENNA__13047__A2 _13087_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12794_ _12794_/A _12798_/B vssd1 vssd1 vccd1 vccd1 _12794_/Y sky130_fd_sc_hd__nand2_1
X_11814_ _09111_/S _10638_/X _11813_/X vssd1 vssd1 vccd1 vccd1 _11814_/Y sky130_fd_sc_hd__a21boi_1
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10805__B2 _10574_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10805__A1 _10575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11745_ _11745_/A _11745_/B vssd1 vssd1 vccd1 vccd1 _11746_/B sky130_fd_sc_hd__or2_1
XFILLER_0_28_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10281__A2 _10574_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11676_ _11768_/B _11676_/B vssd1 vssd1 vccd1 vccd1 _11677_/B sky130_fd_sc_hd__or2_1
XFILLER_0_113_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10627_ _06750_/A _10505_/X _06749_/Y vssd1 vssd1 vccd1 vccd1 _10627_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__09423__A1 _12802_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09423__B2 _09423_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13346_ _13380_/CLK hold71/X vssd1 vssd1 vccd1 vccd1 hold301/A sky130_fd_sc_hd__dfxtp_1
X_10558_ _11146_/A fanout30/X _07688_/B _11294_/A vssd1 vssd1 vccd1 vccd1 _10559_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_3_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13277_ _13378_/CLK hold30/X vssd1 vssd1 vccd1 vccd1 hold29/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09119__S _09142_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09759__A2_N fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09187__A0 _08673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12228_ _12228_/A _12332_/A vssd1 vssd1 vccd1 vccd1 _12228_/Y sky130_fd_sc_hd__nand2_1
X_10489_ _10489_/A _10489_/B vssd1 vssd1 vccd1 vccd1 _10490_/B sky130_fd_sc_hd__xnor2_4
X_12159_ _12159_/A _12159_/B _12159_/C vssd1 vssd1 vccd1 vccd1 _12160_/B sky130_fd_sc_hd__and3_1
XFILLER_0_75_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06720_ reg2_val[13] _06720_/B vssd1 vssd1 vccd1 vccd1 _06720_/X sky130_fd_sc_hd__and2_1
XANTENNA__06986__B _06986_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07163__A _09897_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06651_ _06695_/A _12664_/B vssd1 vssd1 vccd1 vccd1 _06651_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_79_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11836__A3 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08259__A _08724_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13038__A2 _12788_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06582_ instruction[0] pred_val instruction[1] vssd1 vssd1 vccd1 vccd1 _06897_/A
+ sky130_fd_sc_hd__and3b_1
X_09370_ _09163_/X _09364_/Y _12394_/B _09142_/S vssd1 vssd1 vccd1 vccd1 _09371_/C
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_59_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12797__A1 _09251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08465__A2 _08741_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08321_ _08740_/A _08321_/B vssd1 vssd1 vccd1 vccd1 _08322_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_74_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08252_ _08252_/A _08252_/B vssd1 vssd1 vccd1 vccd1 _08295_/A sky130_fd_sc_hd__xor2_1
X_07203_ _10449_/A _07203_/B vssd1 vssd1 vccd1 vccd1 _07208_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_55_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout125_A _10537_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08183_ _08745_/A _08183_/B vssd1 vssd1 vccd1 vccd1 _08187_/B sky130_fd_sc_hd__xnor2_1
X_07134_ _07223_/A _07135_/D vssd1 vssd1 vccd1 vccd1 _07134_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_70_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08722__A _08722_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07065_ _07100_/B _07066_/B _06963_/A vssd1 vssd1 vccd1 vccd1 _07067_/A sky130_fd_sc_hd__o21bai_2
XFILLER_0_71_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07967_ _07854_/A _07854_/B _07854_/C vssd1 vssd1 vccd1 vccd1 _07969_/B sky130_fd_sc_hd__a21oi_1
X_06918_ instruction[20] _06884_/Y _06917_/X _06694_/B vssd1 vssd1 vccd1 vccd1 reg2_idx[2]
+ sky130_fd_sc_hd__o211a_4
X_09706_ _09706_/A _09953_/A _09953_/B _10232_/A vssd1 vssd1 vccd1 vccd1 _09706_/X
+ sky130_fd_sc_hd__or4_1
XANTENNA__06896__B _06896_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07898_ _07897_/B _07897_/C _11564_/A vssd1 vssd1 vccd1 vccd1 _07911_/B sky130_fd_sc_hd__a21o_1
XANTENNA__08153__A1 _07885_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08153__B2 _08721_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06849_ _06838_/Y _06848_/Y _12389_/A vssd1 vssd1 vccd1 vccd1 _06849_/X sky130_fd_sc_hd__o21ba_1
X_09637_ _09637_/A _09637_/B vssd1 vssd1 vccd1 vccd1 _09639_/A sky130_fd_sc_hd__xnor2_4
X_09568_ _09568_/A _09568_/B vssd1 vssd1 vccd1 vccd1 _09570_/C sky130_fd_sc_hd__or2_1
X_08519_ _08519_/A _08519_/B vssd1 vssd1 vccd1 vccd1 _08540_/B sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout38_A _12836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11530_ reg1_val[18] curr_PC[18] vssd1 vssd1 vccd1 vccd1 _11532_/B sky130_fd_sc_hd__nand2_1
X_09499_ _09094_/X _09112_/X _09666_/S vssd1 vssd1 vccd1 vccd1 _09499_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_93_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11460__A1 _07819_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout4_A fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11460__B2 fanout24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11461_ _12073_/A _11461_/B vssd1 vssd1 vccd1 vccd1 _11465_/A sky130_fd_sc_hd__xnor2_1
X_13200_ hold265/X _13213_/A2 _13199_/X _13213_/B2 vssd1 vssd1 vccd1 vccd1 _13201_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_116_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08632__A _08632_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10412_ _10412_/A _10412_/B vssd1 vssd1 vccd1 vccd1 _10490_/A sky130_fd_sc_hd__and2_2
X_11392_ _11392_/A _11392_/B vssd1 vssd1 vccd1 vccd1 _11393_/B sky130_fd_sc_hd__nand2_1
X_13131_ hold273/X _13130_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13131_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_104_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10343_ _10344_/A _10344_/B vssd1 vssd1 vccd1 vccd1 _10345_/A sky130_fd_sc_hd__and2_1
X_13062_ hold92/X _12791_/A _13080_/B1 hold99/X _13128_/A vssd1 vssd1 vccd1 vccd1
+ hold100/A sky130_fd_sc_hd__o221a_1
X_10274_ _09811_/A _09811_/B _09957_/A _09957_/B _09853_/B vssd1 vssd1 vccd1 vccd1
+ _10275_/D sky130_fd_sc_hd__a221oi_2
X_12013_ _12013_/A _12089_/B _12013_/C vssd1 vssd1 vccd1 vccd1 _12093_/A sky130_fd_sc_hd__nand3_2
XANTENNA__07195__A2 _12838_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12915_ hold132/X hold260/A vssd1 vssd1 vccd1 vccd1 _12915_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_88_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12846_ _12846_/A _12848_/B vssd1 vssd1 vccd1 vccd1 _12846_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_0_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12777_ _12777_/A _12777_/B vssd1 vssd1 vccd1 vccd1 _12779_/A sky130_fd_sc_hd__nand2_2
X_11728_ _11727_/A _09527_/B _11727_/Y _12307_/B1 vssd1 vssd1 vccd1 vccd1 _11728_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_83_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11659_ _11847_/A fanout9/X fanout4/X _11766_/A vssd1 vssd1 vccd1 vccd1 _11661_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_126_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13329_ _13340_/CLK _13329_/D vssd1 vssd1 vccd1 vccd1 hold121/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07958__A1 _08798_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07958__B2 _07821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08870_ _08865_/A _08865_/B _08862_/X vssd1 vssd1 vccd1 vccd1 _08885_/A sky130_fd_sc_hd__a21o_1
X_07821_ _07821_/A _09614_/A vssd1 vssd1 vccd1 vccd1 _07822_/C sky130_fd_sc_hd__or2_1
X_07752_ _09614_/A _07752_/B vssd1 vssd1 vccd1 vccd1 _07753_/C sky130_fd_sc_hd__or2_1
X_06703_ reg2_val[16] _06720_/B _06703_/B1 _06702_/Y vssd1 vssd1 vccd1 vccd1 _11343_/A
+ sky130_fd_sc_hd__o2bb2a_4
X_07683_ _07685_/A _07685_/B vssd1 vssd1 vccd1 vccd1 _07683_/X sky130_fd_sc_hd__or2_1
X_06634_ instruction[36] _06634_/B vssd1 vssd1 vccd1 vccd1 _12680_/B sky130_fd_sc_hd__and2_4
X_09422_ _09237_/Y _09244_/X _09245_/A vssd1 vssd1 vccd1 vccd1 _09427_/A sky130_fd_sc_hd__a21o_1
XANTENNA__09312__S _09351_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09353_ _09350_/Y _09351_/Y _09352_/Y vssd1 vssd1 vccd1 vccd1 _09361_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_19_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08436__B _08436_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08304_ _08752_/A _08304_/B vssd1 vssd1 vccd1 vccd1 _08305_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_117_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09284_ _09282_/Y _09284_/B vssd1 vssd1 vccd1 vccd1 _09285_/B sky130_fd_sc_hd__and2b_1
XANTENNA__07110__A2 _09768_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08235_ _08235_/A _08235_/B vssd1 vssd1 vccd1 vccd1 _08287_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__09548__A _09548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09399__B1 _10664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08166_ _08162_/Y _08166_/B vssd1 vssd1 vccd1 vccd1 _08167_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_70_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07117_ _07117_/A vssd1 vssd1 vccd1 vccd1 _07270_/A sky130_fd_sc_hd__inv_2
XFILLER_0_42_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08097_ _08098_/A _08098_/B vssd1 vssd1 vccd1 vccd1 _08097_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_30_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07048_ _07048_/A _07048_/B vssd1 vssd1 vccd1 vccd1 _07048_/X sky130_fd_sc_hd__and2_1
XFILLER_0_100_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09571__B1 _08507_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08999_ _08699_/A _09004_/B _08997_/Y _08623_/Y vssd1 vssd1 vccd1 vccd1 _09000_/B
+ sky130_fd_sc_hd__a211oi_1
XANTENNA__10181__A1 _10445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10181__B2 _10706_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11130__A0 _09527_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10961_ _10961_/A _10961_/B _10961_/C vssd1 vssd1 vccd1 vccd1 _10962_/B sky130_fd_sc_hd__or3_1
XFILLER_0_97_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12700_ _12701_/A _12701_/B _12701_/C vssd1 vssd1 vccd1 vccd1 _12705_/B sky130_fd_sc_hd__a21o_1
X_10892_ _13295_/Q _11633_/B _11014_/B _11968_/B1 vssd1 vssd1 vccd1 vccd1 _10892_/Y
+ sky130_fd_sc_hd__a31oi_1
XFILLER_0_38_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12631_ _12631_/A _12631_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[1] sky130_fd_sc_hd__xor2_4
XFILLER_0_108_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11053__A _11180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12562_ reg1_val[18] curr_PC[18] _12586_/S vssd1 vssd1 vccd1 vccd1 _12564_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_19_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12493_ _12502_/A _12493_/B vssd1 vssd1 vccd1 vccd1 _12495_/C sky130_fd_sc_hd__nand2_1
X_11513_ _11317_/Y _11512_/Y _11510_/X vssd1 vssd1 vccd1 vccd1 _11513_/X sky130_fd_sc_hd__a21bo_1
X_11444_ _12394_/A _11442_/X _11443_/X _09172_/B vssd1 vssd1 vccd1 vccd1 _11444_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__08362__A _09445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11375_ _11908_/A _11375_/B vssd1 vssd1 vccd1 vccd1 _11377_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__08062__B1 _08739_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10944__B1 _11470_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13114_ _12903_/X _13114_/B vssd1 vssd1 vccd1 vccd1 _13115_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_0_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10326_ _10326_/A _10326_/B vssd1 vssd1 vccd1 vccd1 _10328_/B sky130_fd_sc_hd__xnor2_1
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10257_ _09835_/B _10522_/C hold294/A vssd1 vssd1 vccd1 vccd1 _10257_/Y sky130_fd_sc_hd__a21oi_2
X_13045_ _07203_/B _12830_/B hold151/X vssd1 vssd1 vccd1 vccd1 _13325_/D sky130_fd_sc_hd__a21boi_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06610__A _06612_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_59 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10188_ fanout74/X _10571_/B fanout51/X _10948_/B2 vssd1 vssd1 vccd1 vccd1 _10189_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_72_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09865__A1 fanout23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09865__B2 _11171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11672__A1 fanout27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09132__S _09142_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07441__A _09548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06983__C _06986_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11672__B2 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12829_ hold25/X _12830_/B _12828_/Y _13245_/A vssd1 vssd1 vccd1 vccd1 hold26/A sky130_fd_sc_hd__o211a_1
XANTENNA__12059__A _12455_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11975__A2 _11343_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13177__B2 _12790_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08020_ _08021_/A _08021_/B vssd1 vssd1 vccd1 vccd1 _08020_/X sky130_fd_sc_hd__and2_1
XFILLER_0_25_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08272__A _08740_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout7 fanout8/X vssd1 vssd1 vccd1 vccd1 fanout7/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_4_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10307__A _10959_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08053__B1 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09971_ _10248_/S _09320_/X _09970_/X vssd1 vssd1 vccd1 vccd1 _09972_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_40_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08922_ _08922_/A _08922_/B vssd1 vssd1 vccd1 vccd1 _08923_/B sky130_fd_sc_hd__or2_1
XANTENNA__10026__B _10027_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08356__B2 _08739_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08356__A1 _12810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07616__A _10710_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08853_ _08853_/A _08853_/B vssd1 vssd1 vccd1 vccd1 _08857_/A sky130_fd_sc_hd__or2_1
X_07804_ _08722_/A _07804_/B vssd1 vssd1 vccd1 vccd1 _07806_/B sky130_fd_sc_hd__xor2_1
X_08784_ _08252_/A _08252_/B _08212_/Y vssd1 vssd1 vccd1 vccd1 _08787_/B sky130_fd_sc_hd__a21oi_1
X_07735_ _07738_/A _07738_/B vssd1 vssd1 vccd1 vccd1 _07741_/B sky130_fd_sc_hd__or2_1
XANTENNA__10466__A2 _10571_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09405_ _09403_/X _09405_/B vssd1 vssd1 vccd1 vccd1 _09408_/A sky130_fd_sc_hd__and2b_1
X_07666_ _07666_/A _07666_/B vssd1 vssd1 vccd1 vccd1 _08916_/B sky130_fd_sc_hd__xnor2_1
X_06617_ reg1_val[29] _06838_/B vssd1 vssd1 vccd1 vccd1 _06621_/A sky130_fd_sc_hd__nand2_1
X_07597_ _07597_/A _07597_/B vssd1 vssd1 vccd1 vccd1 _07598_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_47_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09336_ _09139_/X _09141_/X _09336_/S vssd1 vssd1 vccd1 vccd1 _09336_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_75_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07619__B1 _11146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09267_ _09266_/B _09266_/C _09746_/A vssd1 vssd1 vccd1 vccd1 _09273_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_90_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08218_ fanout99/X _08732_/A2 _08656_/B _12818_/A vssd1 vssd1 vccd1 vccd1 _08219_/B
+ sky130_fd_sc_hd__o22a_1
X_09198_ _09199_/A _09199_/B vssd1 vssd1 vccd1 vccd1 _09200_/A sky130_fd_sc_hd__or2_1
XFILLER_0_50_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11179__B1 _12067_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08149_ _08147_/Y _08149_/B vssd1 vssd1 vccd1 vccd1 _08150_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_120_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08595__A1 _08730_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08595__B2 _12804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11160_ _11160_/A _11160_/B vssd1 vssd1 vccd1 vccd1 _11188_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_30_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10111_ _11010_/S _09338_/X _09179_/B vssd1 vssd1 vccd1 vccd1 _10111_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11091_ _11092_/A _11092_/B vssd1 vssd1 vccd1 vccd1 _11210_/A sky130_fd_sc_hd__or2_1
X_10042_ _10042_/A _10042_/B _10042_/C vssd1 vssd1 vccd1 vccd1 _10192_/B sky130_fd_sc_hd__or3_1
Xhold30 hold30/A vssd1 vssd1 vccd1 vccd1 hold30/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 hold41/A vssd1 vssd1 vccd1 vccd1 hold41/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11351__B1 _11345_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold63 hold63/A vssd1 vssd1 vccd1 vccd1 hold63/X sky130_fd_sc_hd__clkbuf_2
Xhold74 hold74/A vssd1 vssd1 vccd1 vccd1 hold74/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 hold52/A vssd1 vssd1 vccd1 vccd1 hold52/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold96 hold96/A vssd1 vssd1 vccd1 vccd1 hold96/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 hold85/A vssd1 vssd1 vccd1 vccd1 hold85/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12300__C1 _06924_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11993_ _11993_/A _11993_/B vssd1 vssd1 vccd1 vccd1 _12013_/A sky130_fd_sc_hd__and2_1
XFILLER_0_85_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08357__A _09441_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10944_ _10943_/B _10943_/C _11470_/A vssd1 vssd1 vccd1 vccd1 _10947_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_85_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10875_ _12031_/A _09007_/X _09009_/D _11876_/A vssd1 vssd1 vccd1 vccd1 _10875_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_128_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12614_ _12614_/A _12614_/B vssd1 vssd1 vccd1 vccd1 new_PC[25] sky130_fd_sc_hd__xnor2_4
X_12545_ _12551_/B _12545_/B vssd1 vssd1 vccd1 vccd1 new_PC[14] sky130_fd_sc_hd__and2_4
XANTENNA__07086__A1 _11269_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12476_ reg1_val[5] curr_PC[5] _12622_/S vssd1 vssd1 vccd1 vccd1 _12478_/B sky130_fd_sc_hd__mux2_1
XANTENNA__08092__A _08742_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11427_ _11606_/A _11427_/B vssd1 vssd1 vccd1 vccd1 _11649_/B sky130_fd_sc_hd__xor2_4
XANTENNA_5 instruction[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10917__B1 fanout59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11358_ curr_PC[16] _11357_/C curr_PC[17] vssd1 vssd1 vccd1 vccd1 _11358_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10309_ _10928_/A _10309_/B vssd1 vssd1 vccd1 vccd1 _10312_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__09535__B1 _09354_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09127__S _09127_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12342__A _12423_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11289_ _09745_/B fanout9/X fanout4/X _10418_/A vssd1 vssd1 vccd1 vccd1 _11290_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11342__B1 _12307_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13028_ hold104/X _12788_/A _13236_/B hold296/A _13109_/A vssd1 vssd1 vccd1 vccd1
+ hold105/A sky130_fd_sc_hd__o221a_1
XANTENNA__07436__A _10449_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12437__A3 _11973_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07520_ _07520_/A _07520_/B vssd1 vssd1 vccd1 vccd1 _07558_/A sky130_fd_sc_hd__nand2_1
XANTENNA__10797__A _11065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07171__A _09441_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08510__A1 _08740_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11645__B2 _11876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07451_ _07453_/B _07453_/A vssd1 vssd1 vccd1 vccd1 _07456_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_57_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07382_ _11653_/A _10413_/A _10567_/A fanout66/X vssd1 vssd1 vccd1 vccd1 _07383_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_45_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09121_ _09119_/X _09120_/X _09330_/S vssd1 vssd1 vccd1 vccd1 _09121_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_44_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07077__A1 _10664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12070__A1 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07077__B2 fanout94/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12070__B2 _12316_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09052_ _12106_/A _12031_/B _12031_/C vssd1 vssd1 vccd1 vccd1 _09059_/A sky130_fd_sc_hd__nand3b_2
XFILLER_0_44_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08003_ _08004_/B _08004_/A vssd1 vssd1 vccd1 vccd1 _08003_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_40_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09526__B1 _11624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09954_ _09307_/A _09307_/B _09953_/X vssd1 vssd1 vccd1 vccd1 _09956_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_0_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09885_ _09885_/A _09885_/B vssd1 vssd1 vccd1 vccd1 _09931_/A sky130_fd_sc_hd__xor2_4
X_08905_ _08897_/X _08903_/B _08901_/X vssd1 vssd1 vccd1 vccd1 _08905_/X sky130_fd_sc_hd__a21o_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08836_ _08838_/A _08838_/B vssd1 vssd1 vccd1 vccd1 _08836_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__09829__A1 _12394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08767_ _08767_/A _08767_/B vssd1 vssd1 vccd1 vccd1 _08780_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_94_101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08698_ _08995_/A _08995_/B _09004_/B _08624_/X vssd1 vssd1 vccd1 vccd1 _08699_/B
+ sky130_fd_sc_hd__o211ai_2
X_07718_ _07718_/A _07718_/B vssd1 vssd1 vccd1 vccd1 _07719_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_95_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07649_ _08733_/A _07649_/B vssd1 vssd1 vccd1 vccd1 _07656_/A sky130_fd_sc_hd__xnor2_1
X_10660_ _12031_/A _10782_/A vssd1 vssd1 vccd1 vccd1 _10660_/X sky130_fd_sc_hd__or2_1
XFILLER_0_48_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09319_ _09101_/X _09103_/X _09330_/S vssd1 vssd1 vccd1 vccd1 _09319_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout20_A _09609_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07607__A3 _07087_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10591_ _10700_/A _10592_/A vssd1 vssd1 vccd1 vccd1 _10722_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_50_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12330_ _12330_/A _12330_/B vssd1 vssd1 vccd1 vccd1 _12413_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_23_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12261_ _12261_/A _12261_/B vssd1 vssd1 vccd1 vccd1 _12263_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_105_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11212_ _10988_/A _11098_/A _11098_/B vssd1 vssd1 vccd1 vccd1 _11212_/Y sky130_fd_sc_hd__a21boi_1
X_12192_ _12434_/B1 _12248_/B hold223/A vssd1 vssd1 vccd1 vccd1 _12194_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_101_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11143_ _10783_/B _10871_/Y _10996_/Y _11650_/B _11792_/A vssd1 vssd1 vccd1 vccd1
+ _11218_/A sky130_fd_sc_hd__a41o_1
XANTENNA__10127__A1 _07036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11324__B1 _11649_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11074_ _10926_/A _10926_/B _10923_/A vssd1 vssd1 vccd1 vccd1 _11078_/A sky130_fd_sc_hd__a21o_1
XANTENNA__07791__A2 _08741_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10025_ _07187_/Y fanout7/X _10024_/Y _09433_/A vssd1 vssd1 vccd1 vccd1 _10027_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10678__A2 _10571_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11976_ _10113_/A _10387_/Y _10398_/Y _12254_/A1 _11975_/X vssd1 vssd1 vccd1 vccd1
+ _11976_/X sky130_fd_sc_hd__o221a_1
XANTENNA__08087__A _08742_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10927_ _10927_/A1 _07262_/A _07262_/B fanout36/X _11367_/A vssd1 vssd1 vccd1 vccd1
+ _10928_/B sky130_fd_sc_hd__o32a_1
XFILLER_0_128_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10858_ _10858_/A _10858_/B _10859_/A vssd1 vssd1 vccd1 vccd1 _10858_/X sky130_fd_sc_hd__and3_1
XANTENNA__12052__A1 _09111_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08256__B1 _07752_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10789_ _10789_/A _10789_/B vssd1 vssd1 vccd1 vccd1 _10793_/A sky130_fd_sc_hd__xor2_1
X_12528_ _12537_/A _12528_/B vssd1 vssd1 vccd1 vccd1 _12530_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_81_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12459_ _12460_/A _12460_/B _12460_/C vssd1 vssd1 vccd1 vccd1 _12467_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_112_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09756__B1 _09568_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout309 _12341_/A vssd1 vssd1 vccd1 vccd1 _12423_/A sky130_fd_sc_hd__buf_6
XANTENNA__12072__A _12073_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07166__A _07166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06951_ reg1_val[12] _06951_/B vssd1 vssd1 vccd1 vccd1 _06954_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_118_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09670_ _09176_/A _09669_/X _09974_/A vssd1 vssd1 vccd1 vccd1 _09670_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_118_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06882_ instruction[2] _06897_/A vssd1 vssd1 vccd1 vccd1 _06882_/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_94_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08621_ _08621_/A _08621_/B _08621_/C vssd1 vssd1 vccd1 vccd1 _08622_/B sky130_fd_sc_hd__or3_1
XANTENNA__09381__A _09548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13107__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08552_ _08730_/A1 _12810_/A _08038_/A _12808_/A vssd1 vssd1 vccd1 vccd1 _08553_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_77_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08483_ _08483_/A _08483_/B vssd1 vssd1 vccd1 vccd1 _08493_/B sky130_fd_sc_hd__xnor2_1
X_07503_ reg1_val[29] reg1_val[30] _07503_/C vssd1 vssd1 vccd1 vccd1 _07503_/X sky130_fd_sc_hd__or3_2
XFILLER_0_92_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07434_ _07434_/A _07434_/B vssd1 vssd1 vccd1 vccd1 _07437_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_76_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07365_ reg1_val[30] _07365_/B vssd1 vssd1 vccd1 vccd1 _07508_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_18_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09104_ reg1_val[12] reg1_val[19] _09108_/S vssd1 vssd1 vccd1 vccd1 _09104_/X sky130_fd_sc_hd__mux2_1
XANTENNA__11251__C1 _11250_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07296_ _10165_/A _07296_/B vssd1 vssd1 vccd1 vccd1 _07999_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_33_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08798__B2 _08798_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08798__A1 _08752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09035_ _08719_/B _08786_/Y _08788_/B vssd1 vssd1 vccd1 vccd1 _09043_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_32_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11554__B1 fanout4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09937_ _09787_/A _09787_/B _09785_/Y vssd1 vssd1 vccd1 vccd1 _09939_/B sky130_fd_sc_hd__a21boi_4
XANTENNA__07773__A2 _11653_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07076__A _11164_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09868_ _09869_/A _09869_/B _09869_/C vssd1 vssd1 vccd1 vccd1 _09870_/A sky130_fd_sc_hd__o21ai_2
XANTENNA_fanout68_A fanout69/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06733__B1 _06732_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09799_ _09799_/A _09799_/B vssd1 vssd1 vccd1 vccd1 _09800_/B sky130_fd_sc_hd__xor2_2
XANTENNA__07804__A _08722_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08819_ _08819_/A _08819_/B vssd1 vssd1 vccd1 vccd1 _08834_/A sky130_fd_sc_hd__nor2_1
XANTENNA__09278__A2 _12264_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10230__A _10231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11326__A _11707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11830_ _11831_/B _11830_/B vssd1 vssd1 vccd1 vccd1 _11918_/A sky130_fd_sc_hd__and2b_1
XTAP_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11761_ _11762_/B _11761_/B vssd1 vssd1 vccd1 vccd1 _11763_/A sky130_fd_sc_hd__and2b_1
XTAP_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07828__A3 _07087_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10712_ _10712_/A _10712_/B vssd1 vssd1 vccd1 vccd1 _10714_/A sky130_fd_sc_hd__xnor2_2
XTAP_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08635__A _09442_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11692_ _11693_/A _11693_/B _11693_/C vssd1 vssd1 vccd1 vccd1 _11782_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_119_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10643_ hold203/A _11633_/B _10764_/B _11968_/B1 vssd1 vssd1 vccd1 vccd1 _10643_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_48_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13362_ _13384_/CLK _13362_/D vssd1 vssd1 vccd1 vccd1 hold271/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10574_ _10574_/A _10574_/B vssd1 vssd1 vccd1 vccd1 _10576_/B sky130_fd_sc_hd__or2_1
XFILLER_0_106_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12313_ _07343_/B _12404_/A _12290_/X _12312_/Y _06881_/X vssd1 vssd1 vccd1 vccd1
+ dest_val[28] sky130_fd_sc_hd__a221oi_4
XANTENNA__07461__A1 _10818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11996__A _12317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13293_ _13299_/CLK _13293_/D vssd1 vssd1 vccd1 vccd1 hold203/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09738__B1 _10022_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07461__B2 _10963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12244_ _09821_/X _12243_/Y _12244_/S vssd1 vssd1 vccd1 vccd1 _12244_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10899__A2 _12404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12175_ _12176_/A _12175_/B vssd1 vssd1 vccd1 vccd1 _12175_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__08410__B1 _08564_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11126_ _11126_/A _11126_/B vssd1 vssd1 vccd1 vccd1 _11126_/X sky130_fd_sc_hd__or2_2
XFILLER_0_64_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11057_ fanout66/X _12150_/A _12067_/A _07087_/X vssd1 vssd1 vccd1 vccd1 _11058_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11848__A1 _11847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10008_ _06971_/Y _12214_/A fanout51/X _10445_/A vssd1 vssd1 vccd1 vccd1 _10009_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_98_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12273__A1 fanout59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11959_ _11959_/A _11959_/B vssd1 vssd1 vccd1 vccd1 _11959_/X sky130_fd_sc_hd__or2_1
XFILLER_0_80_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08477__B1 _08673_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_54 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12067__A _12067_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07150_ _07343_/B _07151_/B vssd1 vssd1 vccd1 vccd1 _07150_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_124_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07081_ _07254_/B _06997_/C _07364_/B1 vssd1 vssd1 vccd1 vccd1 _07096_/B sky130_fd_sc_hd__o21ai_2
XFILLER_0_124_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout128 _07222_/Y vssd1 vssd1 vccd1 vccd1 _10022_/B1 sky130_fd_sc_hd__buf_8
Xfanout117 _08741_/B2 vssd1 vssd1 vccd1 vccd1 _11065_/A sky130_fd_sc_hd__buf_6
XFILLER_0_10_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout106 _11987_/A vssd1 vssd1 vccd1 vccd1 _11908_/A sky130_fd_sc_hd__buf_8
Xfanout139 _12810_/A vssd1 vssd1 vccd1 vccd1 _08721_/B1 sky130_fd_sc_hd__buf_6
X_09722_ _09722_/A _09722_/B vssd1 vssd1 vccd1 vccd1 _09724_/A sky130_fd_sc_hd__xnor2_4
X_07983_ _07983_/A _07983_/B vssd1 vssd1 vccd1 vccd1 _07984_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_10_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10034__B _10797_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06934_ _12341_/A is_load _06635_/A _06931_/X vssd1 vssd1 vccd1 vccd1 _06935_/B sky130_fd_sc_hd__a22o_2
X_06865_ _12626_/A _09351_/B vssd1 vssd1 vccd1 vccd1 _06865_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__06715__B1 _06714_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09653_ _09653_/A _09853_/A _09853_/B vssd1 vssd1 vccd1 vccd1 _09655_/B sky130_fd_sc_hd__nand3_1
XANTENNA__09901__B1 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07343__B _07343_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08604_ _08627_/A _08627_/B _08601_/C vssd1 vssd1 vccd1 vccd1 _08605_/C sky130_fd_sc_hd__a21o_1
X_09584_ _09584_/A _09584_/B vssd1 vssd1 vccd1 vccd1 _09588_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__11146__A _11146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10050__A _11470_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08180__A2 _08732_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06796_ reg1_val[2] _10250_/S vssd1 vssd1 vccd1 vccd1 _09684_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_89_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08535_ _08673_/A _08744_/A2 _08564_/B _08798_/B2 vssd1 vssd1 vccd1 vccd1 _08536_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08466_ _08742_/A _08466_/B vssd1 vssd1 vccd1 vccd1 _08495_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_65_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07417_ _07427_/A vssd1 vssd1 vccd1 vccd1 _07417_/Y sky130_fd_sc_hd__inv_2
X_08397_ _08394_/B _08394_/C _08394_/A vssd1 vssd1 vccd1 vccd1 _08398_/B sky130_fd_sc_hd__a21o_1
X_07348_ _07349_/A _07349_/B vssd1 vssd1 vccd1 vccd1 _07348_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__09432__A2 _09567_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_412 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07279_ _10570_/A _10567_/A _10571_/A _10664_/A vssd1 vssd1 vccd1 vccd1 _07280_/B
+ sky130_fd_sc_hd__o22a_1
X_09018_ _09018_/A _09018_/B vssd1 vssd1 vccd1 vccd1 _09018_/Y sky130_fd_sc_hd__nor2_1
X_10290_ _10290_/A _10290_/B vssd1 vssd1 vccd1 vccd1 _10292_/C sky130_fd_sc_hd__xor2_1
Xhold171 hold171/A vssd1 vssd1 vccd1 vccd1 hold171/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold160 hold160/A vssd1 vssd1 vccd1 vccd1 hold160/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09196__B2 _07819_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09196__A1 fanout23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold182 hold182/A vssd1 vssd1 vccd1 vccd1 hold182/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold193 hold193/A vssd1 vssd1 vccd1 vccd1 hold193/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12931_ _13154_/B _13155_/A _12887_/X vssd1 vssd1 vccd1 vccd1 _13160_/A sky130_fd_sc_hd__a21o_1
X_12862_ hold266/X hold31/X vssd1 vssd1 vccd1 vccd1 _13224_/B sky130_fd_sc_hd__nand2b_1
X_11813_ _07135_/D _11343_/B _12254_/A1 _10651_/Y _11812_/X vssd1 vssd1 vccd1 vccd1
+ _11813_/X sky130_fd_sc_hd__o221a_1
XANTENNA__06721__A3 _12698_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12793_ _12264_/B _13087_/B2 hold62/X _13128_/A vssd1 vssd1 vccd1 vccd1 _13250_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10805__A2 fanout48/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11744_ _11745_/A _11745_/B vssd1 vssd1 vccd1 vccd1 _11746_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11675_ _11675_/A _11675_/B vssd1 vssd1 vccd1 vccd1 _11676_/B sky130_fd_sc_hd__and2_1
XANTENNA__09959__B1 _12290_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10626_ _10748_/A _10625_/B _10625_/C vssd1 vssd1 vccd1 vccd1 _10626_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_24_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09423__A2 fanout9/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13345_ _13380_/CLK hold85/X vssd1 vssd1 vccd1 vccd1 hold295/A sky130_fd_sc_hd__dfxtp_1
X_10557_ _10557_/A _10557_/B vssd1 vssd1 vccd1 vccd1 _10561_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_24_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13276_ _13378_/CLK hold42/X vssd1 vssd1 vccd1 vccd1 hold41/A sky130_fd_sc_hd__dfxtp_1
X_10488_ _10489_/A _10489_/B vssd1 vssd1 vccd1 vccd1 _10488_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_122_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12227_ _12095_/X _12332_/A _12334_/A vssd1 vssd1 vccd1 vccd1 _12227_/Y sky130_fd_sc_hd__a21oi_1
X_12158_ _12159_/A _12159_/B _12159_/C vssd1 vssd1 vccd1 vccd1 _12160_/A sky130_fd_sc_hd__a21oi_1
Xclkbuf_4_12_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13357_/CLK sky130_fd_sc_hd__clkbuf_8
X_11109_ _11004_/A _11001_/X _11021_/S vssd1 vssd1 vccd1 vccd1 _11109_/X sky130_fd_sc_hd__a21o_1
X_12089_ _12089_/A _12089_/B _12089_/C vssd1 vssd1 vccd1 vccd1 _12090_/B sky130_fd_sc_hd__nand3_1
XANTENNA__09135__S _09142_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06650_ instruction[33] _06694_/B vssd1 vssd1 vccd1 vccd1 _12664_/B sky130_fd_sc_hd__and2_4
XFILLER_0_78_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06581_ _06926_/A _06581_/B vssd1 vssd1 vccd1 vccd1 is_store sky130_fd_sc_hd__nor2_8
XFILLER_0_87_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08320_ _07752_/B fanout87/X fanout82/X _07955_/A vssd1 vssd1 vccd1 vccd1 _08321_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_19_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08251_ _08249_/A _08249_/B _08250_/Y vssd1 vssd1 vccd1 vccd1 _08252_/B sky130_fd_sc_hd__o21ai_2
X_07202_ _10449_/A _07203_/B vssd1 vssd1 vccd1 vccd1 _07208_/A sky130_fd_sc_hd__or2_1
XFILLER_0_55_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08182_ _08721_/B1 _08744_/A2 _08564_/B _08739_/A1 vssd1 vssd1 vccd1 vccd1 _08183_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_27_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07133_ _07133_/A _07133_/B _07133_/C _07133_/D vssd1 vssd1 vccd1 vccd1 _07220_/C
+ sky130_fd_sc_hd__or4_4
XFILLER_0_70_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06779__A3 _12649_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07064_ _12423_/A _07064_/B _07100_/A vssd1 vssd1 vccd1 vccd1 _07066_/B sky130_fd_sc_hd__and3_1
XANTENNA_fanout118_A _12822_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06753__A_N _07089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07966_ _07966_/A _07966_/B vssd1 vssd1 vccd1 vccd1 _07975_/B sky130_fd_sc_hd__xnor2_2
X_06917_ instruction[27] _06921_/B vssd1 vssd1 vccd1 vccd1 _06917_/X sky130_fd_sc_hd__or2_1
X_09705_ _09953_/B _10232_/A vssd1 vssd1 vccd1 vccd1 _10097_/A sky130_fd_sc_hd__or2_1
XANTENNA__07354__A _07485_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09636_ _09636_/A _09636_/B vssd1 vssd1 vccd1 vccd1 _09637_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_65_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07897_ _11564_/A _07897_/B _07897_/C vssd1 vssd1 vccd1 vccd1 _07911_/A sky130_fd_sc_hd__nand3_1
XANTENNA__08153__A2 fanout87/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06848_ _06839_/Y _06847_/X _06647_/B vssd1 vssd1 vccd1 vccd1 _06848_/Y sky130_fd_sc_hd__a21oi_1
X_06779_ _06805_/A _06686_/A _12649_/B _06778_/X vssd1 vssd1 vccd1 vccd1 _06779_/X
+ sky130_fd_sc_hd__a31o_1
X_09567_ _10941_/B _09567_/B vssd1 vssd1 vccd1 vccd1 _09570_/B sky130_fd_sc_hd__or2_1
X_09498_ _09090_/X _09097_/X _09666_/S vssd1 vssd1 vccd1 vccd1 _09498_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_93_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08518_ _08518_/A _08518_/B vssd1 vssd1 vccd1 vccd1 _08540_/A sky130_fd_sc_hd__xor2_1
X_08449_ _08449_/A _08449_/B vssd1 vssd1 vccd1 vccd1 _08457_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_93_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11460__A2 _12150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11460_ _07819_/B _12150_/A _12067_/A fanout24/X vssd1 vssd1 vccd1 vccd1 _11461_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11748__B1 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10411_ _10361_/A _10361_/B _10359_/X vssd1 vssd1 vccd1 vccd1 _10493_/A sky130_fd_sc_hd__a21o_2
X_11391_ _11392_/A _11392_/B vssd1 vssd1 vccd1 vccd1 _11391_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12960__A2 _13213_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13130_ _13130_/A _13130_/B vssd1 vssd1 vccd1 vccd1 _13130_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__07529__A _09716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10420__B1 _11172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10342_ _10342_/A _10342_/B vssd1 vssd1 vccd1 vccd1 _10344_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_21_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13061_ _11470_/B _13087_/B2 hold93/X vssd1 vssd1 vccd1 vccd1 hold94/A sky130_fd_sc_hd__o21a_1
X_10273_ _10780_/A _10270_/X _10271_/X _10272_/Y vssd1 vssd1 vccd1 vccd1 dest_val[7]
+ sky130_fd_sc_hd__a22o_4
X_12012_ _12012_/A _12012_/B _12012_/C vssd1 vssd1 vccd1 vccd1 _12013_/C sky130_fd_sc_hd__nand3_1
XANTENNA__08392__A2 _08393_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12914_ hold244/X hold27/X vssd1 vssd1 vccd1 vccd1 _13096_/B sky130_fd_sc_hd__nand2b_1
X_12845_ hold41/X _12848_/B _12844_/Y _13210_/A vssd1 vssd1 vccd1 vccd1 hold42/A sky130_fd_sc_hd__o211a_1
XFILLER_0_69_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12776_ reg1_val[30] _12782_/A vssd1 vssd1 vccd1 vccd1 _12777_/B sky130_fd_sc_hd__nand2_1
X_11727_ _11727_/A _11973_/B vssd1 vssd1 vccd1 vccd1 _11727_/Y sky130_fd_sc_hd__nand2_1
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11658_ _11770_/A _11658_/B vssd1 vssd1 vccd1 vccd1 _11663_/A sky130_fd_sc_hd__nor2_1
XANTENNA__12400__A1 _08979_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11589_ _11589_/A _11589_/B vssd1 vssd1 vccd1 vccd1 _11591_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_4_727 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10609_ _10611_/A _10611_/B vssd1 vssd1 vccd1 vccd1 _10609_/X sky130_fd_sc_hd__and2_1
XFILLER_0_24_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13328_ _13343_/CLK hold154/X vssd1 vssd1 vccd1 vccd1 hold162/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07958__A2 _07087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13259_ _13355_/CLK hold56/X vssd1 vssd1 vccd1 vccd1 hold55/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07820_ _07033_/A _07033_/B _08671_/B2 vssd1 vssd1 vccd1 vccd1 _07822_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_19_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07751_ _07033_/A _07033_/B _07821_/A vssd1 vssd1 vccd1 vccd1 _07753_/B sky130_fd_sc_hd__a21o_1
X_06702_ _06702_/A _12629_/B vssd1 vssd1 vccd1 vccd1 _06702_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07682_ _08968_/A _08968_/B _07601_/X vssd1 vssd1 vccd1 vccd1 _07685_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_126_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06633_ _12126_/S _06633_/B vssd1 vssd1 vccd1 vccd1 _12110_/A sky130_fd_sc_hd__or2_2
X_09421_ _12798_/A _12316_/B vssd1 vssd1 vccd1 vccd1 _09429_/A sky130_fd_sc_hd__or2_1
XFILLER_0_35_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09352_ _09350_/Y _09351_/Y _11624_/A vssd1 vssd1 vccd1 vccd1 _09352_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_59_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08303_ _08722_/A _08303_/B vssd1 vssd1 vccd1 vccd1 _08370_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09283_ _09283_/A _09283_/B vssd1 vssd1 vccd1 vccd1 _09284_/B sky130_fd_sc_hd__nand2_1
XANTENNA__10650__B1 _10648_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08234_ _08722_/A _08234_/B vssd1 vssd1 vccd1 vccd1 _08287_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__08733__A _08733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13195__A2 _13213_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09399__A1 _07033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08165_ _08752_/A _09396_/B _08166_/B vssd1 vssd1 vccd1 vccd1 _08167_/A sky130_fd_sc_hd__or3_1
XFILLER_0_27_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07116_ _07116_/A _07116_/B vssd1 vssd1 vccd1 vccd1 _07117_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_42_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08096_ _08096_/A _08096_/B vssd1 vssd1 vccd1 vccd1 _08098_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_113_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07047_ _11180_/A _11987_/B _11172_/A vssd1 vssd1 vccd1 vccd1 _07048_/B sky130_fd_sc_hd__or3b_2
XFILLER_0_100_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09571__A1 _10571_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09571__B2 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08998_ _08623_/Y _08997_/Y _09004_/B _08699_/A vssd1 vssd1 vccd1 vccd1 _09000_/A
+ sky130_fd_sc_hd__o211a_1
XANTENNA__10181__A2 _12214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07949_ _07949_/A _07949_/B vssd1 vssd1 vccd1 vccd1 _08033_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__11130__A1 _09354_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout50_A fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10960_ _10833_/A _10961_/C vssd1 vssd1 vccd1 vccd1 _10962_/A sky130_fd_sc_hd__nand2b_1
X_10891_ _11633_/B _11014_/B _13295_/Q vssd1 vssd1 vccd1 vccd1 _10891_/X sky130_fd_sc_hd__a21o_1
X_09619_ _09617_/X _09619_/B vssd1 vssd1 vccd1 vccd1 _09622_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_78_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12630_ _12630_/A _12630_/B vssd1 vssd1 vccd1 vccd1 _12631_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_38_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12561_ _12566_/B _12561_/B vssd1 vssd1 vccd1 vccd1 new_PC[17] sky130_fd_sc_hd__xnor2_4
XFILLER_0_108_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12492_ _12659_/B _12492_/B vssd1 vssd1 vccd1 vccd1 _12493_/B sky130_fd_sc_hd__or2_1
XFILLER_0_65_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09739__A _10449_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11512_ _11702_/A vssd1 vssd1 vccd1 vccd1 _11512_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_19_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13186__A2 _13213_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11443_ _12244_/S _11443_/B vssd1 vssd1 vccd1 vccd1 _11443_/X sky130_fd_sc_hd__or2_1
XFILLER_0_123_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08062__A1 _10537_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13113_ _13113_/A hold259/X vssd1 vssd1 vccd1 vccd1 _13352_/D sky130_fd_sc_hd__and2_1
X_11374_ _09613_/A _12150_/A _12213_/A _09614_/A vssd1 vssd1 vccd1 vccd1 _11375_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08062__B2 _08432_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10325_ _10326_/A _10326_/B vssd1 vssd1 vccd1 vccd1 _10474_/A sky130_fd_sc_hd__nand2b_1
X_10256_ hold242/A _10256_/B vssd1 vssd1 vccd1 vccd1 _10522_/C sky130_fd_sc_hd__or2_1
X_13044_ hold142/X _12788_/A _13080_/B1 hold150/X _13109_/A vssd1 vssd1 vccd1 vccd1
+ hold151/A sky130_fd_sc_hd__o221a_1
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10413__A _10413_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10187_ _10187_/A _10187_/B vssd1 vssd1 vccd1 vccd1 _10190_/A sky130_fd_sc_hd__or2_1
XFILLER_0_88_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09865__A2 _10818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11672__A2 _12150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12828_ _12828_/A _12830_/B vssd1 vssd1 vccd1 vccd1 _12828_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_118_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12759_ reg1_val[26] _12782_/A _12758_/A vssd1 vssd1 vccd1 vccd1 _12761_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_127_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08553__A _08681_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13177__A2 _12789_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07169__A _07169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12385__B1 _12290_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout8 fanout8/A vssd1 vssd1 vccd1 vccd1 fanout8/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__08053__B2 fanout99/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08053__A1 _08436_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09970_ _09974_/A _09970_/B vssd1 vssd1 vccd1 vccd1 _09970_/X sky130_fd_sc_hd__or2_1
XFILLER_0_40_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12137__B1 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08921_ _08922_/A _08922_/B vssd1 vssd1 vccd1 vccd1 _08923_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08356__A2 _09238_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08852_ _08726_/A _08726_/B _08793_/B _08794_/Y vssd1 vssd1 vccd1 vccd1 _08858_/A
+ sky130_fd_sc_hd__o31ai_4
X_07803_ _10537_/A1 fanout99/X _12818_/A _08432_/B vssd1 vssd1 vccd1 vccd1 _07804_/B
+ sky130_fd_sc_hd__o22a_1
X_08783_ _08783_/A _08783_/B vssd1 vssd1 vccd1 vccd1 _08786_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_79_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07734_ _08724_/A _07734_/B vssd1 vssd1 vccd1 vccd1 _07738_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07665_ _07995_/A _07995_/B _07658_/Y vssd1 vssd1 vccd1 vccd1 _08916_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__08728__A _08728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06616_ _06615_/Y _06703_/B1 _06771_/A reg2_val[29] vssd1 vssd1 vccd1 vccd1 _06838_/B
+ sky130_fd_sc_hd__a2bb2o_4
X_09404_ _09404_/A _09404_/B _09404_/C _09404_/D vssd1 vssd1 vccd1 vccd1 _09405_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_0_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07596_ _07597_/A _07597_/B vssd1 vssd1 vccd1 vccd1 _07596_/X sky130_fd_sc_hd__and2_1
XFILLER_0_48_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09335_ _09135_/X _09138_/X _09336_/S vssd1 vssd1 vccd1 vccd1 _09335_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_63_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07619__A1 _10445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07619__B2 _10706_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08463__A _08745_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09266_ _09746_/A _09266_/B _09266_/C vssd1 vssd1 vccd1 vccd1 _09273_/A sky130_fd_sc_hd__and3_1
XFILLER_0_117_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08217_ _11385_/A _08285_/A _08285_/B vssd1 vssd1 vccd1 vccd1 _08238_/A sky130_fd_sc_hd__mux2_1
X_09197_ _09716_/A _09197_/B vssd1 vssd1 vccd1 vccd1 _09199_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_62_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11179__A1 _10574_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11179__B2 _10575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08148_ _08148_/A _08148_/B vssd1 vssd1 vccd1 vccd1 _08149_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08595__A2 _08723_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08079_ _08891_/A _08891_/B vssd1 vssd1 vccd1 vccd1 _08079_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_101_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10110_ _10109_/A _10109_/B _09156_/Y vssd1 vssd1 vccd1 vccd1 _10110_/X sky130_fd_sc_hd__o21a_1
XANTENNA__12128__B1 _12254_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout98_A fanout99/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11090_ _11090_/A _11090_/B vssd1 vssd1 vccd1 vccd1 _11092_/B sky130_fd_sc_hd__xnor2_1
X_10041_ _10040_/A _10040_/B _10040_/C vssd1 vssd1 vccd1 vccd1 _10042_/C sky130_fd_sc_hd__a21oi_1
Xhold31 hold31/A vssd1 vssd1 vccd1 vccd1 hold31/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold20 hold20/A vssd1 vssd1 vccd1 vccd1 hold20/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11351__A1 _09172_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11887__C1 _06924_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold53 hold53/A vssd1 vssd1 vccd1 vccd1 hold53/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 hold42/A vssd1 vssd1 vccd1 vccd1 hold42/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 hold64/A vssd1 vssd1 vccd1 vccd1 hold64/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold86 hold86/A vssd1 vssd1 vccd1 vccd1 hold86/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 hold75/A vssd1 vssd1 vccd1 vccd1 hold75/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 hold97/A vssd1 vssd1 vccd1 vccd1 hold97/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11639__C1 _12307_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11992_ _11992_/A _11992_/B _11992_/C vssd1 vssd1 vccd1 vccd1 _11993_/B sky130_fd_sc_hd__or3_1
XANTENNA__09847__A2 _09821_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10943_ _11470_/A _10943_/B _10943_/C vssd1 vssd1 vccd1 vccd1 _10947_/B sky130_fd_sc_hd__nand3_1
XANTENNA__12851__A1 _12264_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11064__A _12261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10874_ _12031_/A _09007_/X _09009_/D vssd1 vssd1 vccd1 vccd1 _10874_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_128_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12613_ _12611_/A _12604_/B _12608_/A _12608_/B vssd1 vssd1 vccd1 vccd1 _12614_/B
+ sky130_fd_sc_hd__o2bb2a_2
X_12544_ _12544_/A _12544_/B _12544_/C vssd1 vssd1 vccd1 vccd1 _12545_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_93_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07086__A2 _07090_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12475_ _12481_/B _12475_/B vssd1 vssd1 vccd1 vccd1 new_PC[4] sky130_fd_sc_hd__and2_4
XFILLER_0_53_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_6 instruction[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11426_ _11426_/A _11426_/B _11425_/X vssd1 vssd1 vccd1 vccd1 _11427_/B sky130_fd_sc_hd__or3b_4
XFILLER_0_1_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10917__A1 _10570_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11357_ curr_PC[16] curr_PC[17] _11357_/C vssd1 vssd1 vccd1 vccd1 _11550_/B sky130_fd_sc_hd__and3_1
XFILLER_0_6_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10917__B2 _10571_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10308_ _10664_/A fanout16/X _07282_/B _10818_/A vssd1 vssd1 vccd1 vccd1 _10309_/B
+ sky130_fd_sc_hd__o22a_1
X_13027_ _09593_/A _13077_/A2 hold112/X vssd1 vssd1 vccd1 vccd1 _13316_/D sky130_fd_sc_hd__o21a_1
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11288_ _11288_/A _11288_/B vssd1 vssd1 vccd1 vccd1 _11297_/A sky130_fd_sc_hd__xnor2_1
X_10239_ _09653_/A _08994_/A _08994_/B vssd1 vssd1 vccd1 vccd1 _10239_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_89_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09838__A2 _11343_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10797__B _10797_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07450_ _07334_/B _07337_/B _07334_/A vssd1 vssd1 vccd1 vccd1 _07453_/B sky130_fd_sc_hd__o21ba_1
XFILLER_0_76_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07381_ _09746_/A _07381_/B vssd1 vssd1 vccd1 vccd1 _07385_/A sky130_fd_sc_hd__xnor2_1
X_09120_ reg1_val[11] reg1_val[20] _09142_/S vssd1 vssd1 vccd1 vccd1 _09120_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_45_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07077__A2 _10941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09051_ _09056_/A _09065_/C vssd1 vssd1 vccd1 vccd1 _12106_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__12070__A2 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08002_ _08002_/A _08002_/B vssd1 vssd1 vccd1 vccd1 _08004_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_4_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout100_A _11385_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12533__A _12692_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09318__S _09351_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07785__B1 _11558_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09953_ _09953_/A _09953_/B _10232_/A _10368_/A vssd1 vssd1 vccd1 vccd1 _09953_/X
+ sky130_fd_sc_hd__or4_1
X_09884_ _09884_/A _09884_/B vssd1 vssd1 vccd1 vccd1 _09885_/B sky130_fd_sc_hd__xor2_4
X_08904_ _09049_/B _09056_/A vssd1 vssd1 vccd1 vccd1 _08904_/Y sky130_fd_sc_hd__nand2_1
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08835_ _08835_/A _08835_/B vssd1 vssd1 vccd1 vccd1 _08838_/B sky130_fd_sc_hd__xnor2_4
X_08766_ _08766_/A _08766_/B vssd1 vssd1 vccd1 vccd1 _08767_/B sky130_fd_sc_hd__nor2_2
XANTENNA__09829__A2 _09172_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07717_ _07718_/A _07718_/B vssd1 vssd1 vccd1 vccd1 _07717_/X sky130_fd_sc_hd__and2b_1
XANTENNA__12294__C1 _09156_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08697_ _08697_/A _08697_/B vssd1 vssd1 vccd1 vccd1 _09004_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_94_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07648_ _08656_/B _11847_/A _11766_/A _08732_/A2 vssd1 vssd1 vccd1 vccd1 _07649_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_94_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07579_ _07579_/A _07579_/B _07579_/C vssd1 vssd1 vccd1 vccd1 _07580_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_48_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09318_ _09100_/X _09127_/X _09351_/B vssd1 vssd1 vccd1 vccd1 _09318_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_48_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout13_A _12854_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10590_ _10710_/A _10590_/B vssd1 vssd1 vccd1 vccd1 _10700_/A sky130_fd_sc_hd__xnor2_2
X_09249_ _09249_/A _09379_/A _09249_/C vssd1 vssd1 vccd1 vccd1 _09379_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_35_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12260_ fanout12/X fanout9/A fanout5/X _12316_/A vssd1 vssd1 vccd1 vccd1 _12261_/B
+ sky130_fd_sc_hd__o22a_1
X_12191_ hold207/A _12191_/B vssd1 vssd1 vccd1 vccd1 _12248_/B sky130_fd_sc_hd__or2_1
XANTENNA__11021__A0 _09527_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07225__C1 _07135_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11211_ _11211_/A _11211_/B vssd1 vssd1 vccd1 vccd1 _11421_/A sky130_fd_sc_hd__nor2_2
X_11142_ _11138_/X _11141_/Y _11142_/S vssd1 vssd1 vccd1 vccd1 dest_val[14] sky130_fd_sc_hd__mux2_8
XANTENNA__07537__A _11987_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10127__A2 _12404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07528__B1 _11171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11073_ _11073_/A _11073_/B vssd1 vssd1 vccd1 vccd1 _11079_/A sky130_fd_sc_hd__nor2_1
X_10024_ _10024_/A fanout7/X vssd1 vssd1 vccd1 vccd1 _10024_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__13077__A1 _07013_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11975_ _07194_/A _11343_/B _11974_/X _06655_/B vssd1 vssd1 vccd1 vccd1 _11975_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_85_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10926_ _10926_/A _10926_/B vssd1 vssd1 vccd1 vccd1 _10956_/A sky130_fd_sc_hd__xor2_1
XANTENNA__07700__B1 _11923_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10857_ _10859_/A _10859_/B vssd1 vssd1 vccd1 vccd1 _10857_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_27_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08256__A1 _10537_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08256__B2 _08432_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10788_ _10789_/A _10789_/B vssd1 vssd1 vccd1 vccd1 _10913_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_26_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12527_ _12686_/B _12527_/B vssd1 vssd1 vccd1 vccd1 _12528_/B sky130_fd_sc_hd__or2_1
XFILLER_0_42_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11260__B1 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12458_ _12467_/A _12458_/B vssd1 vssd1 vccd1 vccd1 _12460_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_78_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09756__A1 _09568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09756__B2 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11409_ _11410_/A _11410_/B vssd1 vssd1 vccd1 vccd1 _11504_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_22_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09138__S _09142_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12389_ _12389_/A _12389_/B vssd1 vssd1 vccd1 vccd1 _12389_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__09646__B _09647_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06950_ reg1_val[10] reg1_val[11] _07200_/B _07200_/A vssd1 vssd1 vccd1 vccd1 _06951_/B
+ sky130_fd_sc_hd__o31a_2
X_06881_ instruction[2] _06897_/A vssd1 vssd1 vccd1 vccd1 _06881_/X sky130_fd_sc_hd__and2_4
XFILLER_0_94_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12800__B _12818_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_10_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08620_ _09433_/A _08628_/B _08628_/A vssd1 vssd1 vccd1 vccd1 _08621_/C sky130_fd_sc_hd__mux2_1
XFILLER_0_118_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07182__A _07200_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08551_ _09441_/A _08551_/B vssd1 vssd1 vccd1 vccd1 _08558_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__10320__B fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07502_ _07502_/A _07502_/B vssd1 vssd1 vccd1 vccd1 _07517_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_77_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08482_ _08518_/A _08481_/B _08474_/X vssd1 vssd1 vccd1 vccd1 _08493_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__09692__B1 _09167_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07433_ _07433_/A _07433_/B vssd1 vssd1 vccd1 vccd1 _07434_/B sky130_fd_sc_hd__and2_1
XFILLER_0_92_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout148_A _07026_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13240__B2 _06572_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09103_ reg1_val[13] reg1_val[18] _09108_/S vssd1 vssd1 vccd1 vccd1 _09103_/X sky130_fd_sc_hd__mux2_1
X_07364_ reg1_val[29] _07503_/C _07364_/B1 vssd1 vssd1 vccd1 vccd1 _07365_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_115_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09995__B2 _11876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07295_ _09567_/B _11751_/A _11766_/A _09568_/B vssd1 vssd1 vccd1 vccd1 _07296_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_45_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08798__A2 _07087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09034_ _11616_/C _11521_/B _11521_/C _11709_/A vssd1 vssd1 vccd1 vccd1 _11792_/B
+ sky130_fd_sc_hd__and4b_1
XFILLER_0_4_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10990__B _11100_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11554__B2 _11751_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11554__A1 _11766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09936_ _09775_/A _09775_/B _09773_/Y vssd1 vssd1 vccd1 vccd1 _09939_/A sky130_fd_sc_hd__o21a_2
XANTENNA__07076__B _07076_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09572__A _10444_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09867_ _09867_/A _09867_/B vssd1 vssd1 vccd1 vccd1 _09869_/C sky130_fd_sc_hd__xnor2_1
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13059__A1 _11385_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09798_ _09798_/A _09798_/B vssd1 vssd1 vccd1 vccd1 _09799_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__07092__A _11261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08818_ _08817_/B _08817_/C _08817_/A vssd1 vssd1 vccd1 vccd1 _08819_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_68_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10230__B _10231_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08749_ _08749_/A _08749_/B vssd1 vssd1 vccd1 vccd1 _08761_/A sky130_fd_sc_hd__xnor2_1
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11760_ _11908_/A _11760_/B vssd1 vssd1 vccd1 vccd1 _11761_/B sky130_fd_sc_hd__xnor2_1
XTAP_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10711_ _10712_/A _10712_/B vssd1 vssd1 vccd1 vccd1 _10711_/Y sky130_fd_sc_hd__nand2b_1
XTAP_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10657__S _11142_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11691_ _11691_/A _11691_/B vssd1 vssd1 vccd1 vccd1 _11693_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__13231__B2 _12790_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10642_ _11633_/B _10764_/B hold203/A vssd1 vssd1 vccd1 vccd1 _10642_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_82_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11242__B1 _12247_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13361_ _13384_/CLK _13361_/D vssd1 vssd1 vccd1 vccd1 hold279/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10573_ _10572_/B _10572_/C _11269_/A vssd1 vssd1 vccd1 vccd1 _10579_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_8_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13292_ _13299_/CLK _13292_/D vssd1 vssd1 vccd1 vccd1 hold232/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12312_ _12312_/A _12312_/B vssd1 vssd1 vccd1 vccd1 _12312_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__07461__A2 _10570_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12243_ _12243_/A _12243_/B vssd1 vssd1 vccd1 vccd1 _12243_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__09738__A1 fanout59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09738__B2 _10941_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07749__B1 _11766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10753__C1 _09156_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12174_ _06855_/X _12176_/B _12174_/S vssd1 vssd1 vccd1 vccd1 _12175_/B sky130_fd_sc_hd__mux2_1
XANTENNA__08410__A1 _09423_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08410__B2 _07955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11125_ hold279/A _11452_/B1 _11240_/B _12247_/C1 vssd1 vssd1 vccd1 vccd1 _11126_/B
+ sky130_fd_sc_hd__a31o_1
XANTENNA__06972__A1 _11343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11056_ _11056_/A _11056_/B vssd1 vssd1 vccd1 vccd1 _11059_/A sky130_fd_sc_hd__nor2_1
XANTENNA__13208__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10007_ _10211_/B _10007_/B vssd1 vssd1 vccd1 vccd1 _10047_/A sky130_fd_sc_hd__or2_2
XANTENNA__11848__A2 _12214_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_49 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08477__A1 _07885_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11958_ _11959_/A _11959_/B vssd1 vssd1 vccd1 vccd1 _11958_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__08477__B2 _08721_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11889_ _11636_/B _11970_/B hold246/A vssd1 vssd1 vccd1 vccd1 _11889_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_86_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10909_ _10782_/A _10782_/B _10871_/Y _12031_/A vssd1 vssd1 vccd1 vccd1 _10909_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_58_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13222__B2 _12790_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12067__B _12214_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07080_ _07080_/A _07080_/B vssd1 vssd1 vccd1 vccd1 _10148_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_125_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout129 _10167_/A1 vssd1 vssd1 vccd1 vccd1 _08744_/A2 sky130_fd_sc_hd__buf_6
X_07982_ _07808_/A _07706_/B _07704_/Y vssd1 vssd1 vccd1 vccd1 _07989_/A sky130_fd_sc_hd__o21a_1
Xfanout118 _12822_/A vssd1 vssd1 vccd1 vccd1 _08741_/B2 sky130_fd_sc_hd__buf_6
XFILLER_0_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout107 _07524_/A vssd1 vssd1 vccd1 vccd1 _11987_/A sky130_fd_sc_hd__buf_8
X_06933_ _12455_/S _06933_/B vssd1 vssd1 vccd1 vccd1 dest_mask[0] sky130_fd_sc_hd__nand2_8
X_09721_ _11673_/A _09721_/B vssd1 vssd1 vccd1 vccd1 _09722_/B sky130_fd_sc_hd__xnor2_4
X_06864_ _07149_/A _09336_/S vssd1 vssd1 vccd1 vccd1 _08680_/A sky130_fd_sc_hd__nor2_2
X_09652_ _10232_/A _09652_/B vssd1 vssd1 vccd1 vccd1 _09853_/B sky130_fd_sc_hd__xor2_4
XANTENNA__09901__A1 _10445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09901__B2 _10706_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06795_ reg1_val[2] _09974_/A vssd1 vssd1 vccd1 vccd1 _06795_/X sky130_fd_sc_hd__and2_1
X_08603_ _09433_/A _08603_/B vssd1 vssd1 vccd1 vccd1 _08605_/B sky130_fd_sc_hd__xor2_1
X_09583_ _09584_/A _09584_/B vssd1 vssd1 vccd1 vccd1 _09732_/A sky130_fd_sc_hd__nor2_1
XANTENNA__11146__B _12214_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout265_A _12455_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08534_ _08742_/A _08534_/B vssd1 vssd1 vccd1 vccd1 _08573_/A sky130_fd_sc_hd__xnor2_1
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09331__S _09669_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06955__S _10707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08465_ _12802_/A _08741_/A2 _09568_/B _07896_/A vssd1 vssd1 vccd1 vccd1 _08466_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_65_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07416_ _09445_/A _07416_/B vssd1 vssd1 vccd1 vccd1 _07427_/A sky130_fd_sc_hd__xnor2_4
X_08396_ _08598_/A _08396_/B vssd1 vssd1 vccd1 vccd1 _08447_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__11162__A _11564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07347_ _09442_/A _07347_/B vssd1 vssd1 vccd1 vccd1 _07349_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_9_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09567__A _10941_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09017_ _09017_/A _09017_/B vssd1 vssd1 vccd1 vccd1 _11107_/C sky130_fd_sc_hd__xnor2_1
X_07278_ _07278_/A _07278_/B vssd1 vssd1 vccd1 vccd1 _07281_/A sky130_fd_sc_hd__xor2_1
Xhold161 hold161/A vssd1 vssd1 vccd1 vccd1 hold161/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold150 hold150/A vssd1 vssd1 vccd1 vccd1 hold150/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09196__A2 _12810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07087__A _07087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold194 hold194/A vssd1 vssd1 vccd1 vccd1 hold194/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold183 hold183/A vssd1 vssd1 vccd1 vccd1 hold183/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 hold297/A vssd1 vssd1 vccd1 vccd1 hold172/X sky130_fd_sc_hd__buf_1
XANTENNA__09506__S _09669_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout80_A _12832_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09919_ _12810_/A _07262_/A _07262_/B fanout36/X _10413_/A vssd1 vssd1 vccd1 vccd1
+ _09920_/B sky130_fd_sc_hd__o32a_1
X_12930_ _13149_/B _13150_/A _12889_/X vssd1 vssd1 vccd1 vccd1 _13155_/A sky130_fd_sc_hd__a21o_1
X_12861_ hold31/X hold266/X vssd1 vssd1 vccd1 vccd1 _12861_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_87_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11812_ _12307_/B1 _11811_/X _06675_/B vssd1 vssd1 vccd1 vccd1 _11812_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_68_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12792_ hold61/X _12856_/B vssd1 vssd1 vccd1 vccd1 hold62/A sky130_fd_sc_hd__or2_1
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11743_ _12210_/A _11743_/B vssd1 vssd1 vccd1 vccd1 _11745_/B sky130_fd_sc_hd__xnor2_1
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11674_ _11675_/A _11675_/B vssd1 vssd1 vccd1 vccd1 _11768_/B sky130_fd_sc_hd__nor2_1
X_10625_ _10748_/A _10625_/B _10625_/C vssd1 vssd1 vccd1 vccd1 _10625_/X sky130_fd_sc_hd__or3_1
XFILLER_0_64_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13344_ _13380_/CLK hold75/X vssd1 vssd1 vccd1 vccd1 hold82/A sky130_fd_sc_hd__dfxtp_1
X_10556_ _11172_/A _10556_/B vssd1 vssd1 vccd1 vccd1 _10557_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13275_ _13285_/CLK hold20/X vssd1 vssd1 vccd1 vccd1 hold19/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10487_ _10487_/A _10487_/B vssd1 vssd1 vccd1 vccd1 _10489_/B sky130_fd_sc_hd__xnor2_4
X_12226_ _12226_/A _12280_/A vssd1 vssd1 vccd1 vccd1 _12332_/A sky130_fd_sc_hd__nor2_1
XANTENNA__08395__B1 _08727_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12157_ _12157_/A _12157_/B vssd1 vssd1 vccd1 vccd1 _12159_/C sky130_fd_sc_hd__nand2_1
X_11108_ _12031_/A _11107_/B _11107_/C vssd1 vssd1 vccd1 vccd1 _11108_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__10772__A2_N _12404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12088_ _12089_/A _12089_/B _12089_/C vssd1 vssd1 vccd1 vccd1 _12159_/B sky130_fd_sc_hd__a21o_1
XANTENNA__09895__B1 _10022_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11039_ _11040_/A _11040_/B vssd1 vssd1 vccd1 vccd1 _11183_/A sky130_fd_sc_hd__and2_1
XANTENNA__10151__A _10928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06580_ instruction[3] _06581_/B vssd1 vssd1 vccd1 vccd1 is_load sky130_fd_sc_hd__nor2_8
XANTENNA__08556__A _08728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08250_ _08254_/B _08254_/A vssd1 vssd1 vccd1 vccd1 _08250_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_117_527 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07201_ reg1_val[10] _07201_/B vssd1 vssd1 vccd1 vccd1 _07203_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_74_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08181_ _08733_/A _08181_/B vssd1 vssd1 vccd1 vccd1 _08187_/A sky130_fd_sc_hd__xnor2_1
X_07132_ _07133_/A _07133_/B _07133_/C _07133_/D vssd1 vssd1 vccd1 vccd1 _07142_/B
+ sky130_fd_sc_hd__nor4_2
XFILLER_0_70_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06804__A _09343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_755 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07063_ _07095_/A _07089_/A _06964_/A _06964_/B _07074_/B vssd1 vssd1 vccd1 vccd1
+ _07100_/B sky130_fd_sc_hd__o41a_4
XFILLER_0_30_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07189__A1 _09433_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12541__A _12698_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09326__S _09351_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07965_ _08028_/A _08028_/B _07942_/Y vssd1 vssd1 vccd1 vccd1 _07975_/A sky130_fd_sc_hd__a21oi_2
X_06916_ instruction[19] _06884_/Y _06915_/X _06694_/B vssd1 vssd1 vccd1 vccd1 reg2_idx[1]
+ sky130_fd_sc_hd__o211a_4
X_09704_ _09853_/A _09853_/B _09653_/A vssd1 vssd1 vccd1 vccd1 _09704_/X sky130_fd_sc_hd__o21a_1
XANTENNA__11157__A _12210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09635_ _09633_/A _09633_/B _09636_/B vssd1 vssd1 vccd1 vccd1 _09635_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_69_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07896_ _07896_/A _09396_/B vssd1 vssd1 vccd1 vccd1 _07897_/C sky130_fd_sc_hd__or2_1
X_06847_ _06840_/Y _06846_/Y _12293_/A vssd1 vssd1 vccd1 vccd1 _06847_/X sky130_fd_sc_hd__a21o_1
X_06778_ reg2_val[4] _06799_/B vssd1 vssd1 vccd1 vccd1 _06778_/X sky130_fd_sc_hd__and2_2
XANTENNA__08466__A _08742_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09566_ _09566_/A _09566_/B vssd1 vssd1 vccd1 vccd1 _09607_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__11445__B1 _12307_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09497_ _10119_/S _09496_/A _09181_/X vssd1 vssd1 vccd1 vccd1 _09497_/Y sky130_fd_sc_hd__o21ai_2
X_08517_ _08517_/A _08517_/B vssd1 vssd1 vccd1 vccd1 _08543_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_92_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08448_ _08492_/A _08492_/B _08445_/Y vssd1 vssd1 vccd1 vccd1 _08457_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_18_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10410_ _10410_/A _10658_/B vssd1 vssd1 vccd1 vccd1 _10410_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_61_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08379_ _08379_/A _08379_/B vssd1 vssd1 vccd1 vccd1 _08424_/B sky130_fd_sc_hd__xor2_2
XANTENNA__11748__B2 _12067_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11748__A1 _11989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09297__A _09298_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11390_ _11475_/B _11390_/B vssd1 vssd1 vccd1 vccd1 _11392_/B sky130_fd_sc_hd__or2_1
XFILLER_0_104_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10341_ _10341_/A _10341_/B vssd1 vssd1 vccd1 vccd1 _10342_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_103_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13060_ hold137/A _12791_/A _13080_/B1 hold92/X _13128_/A vssd1 vssd1 vccd1 vccd1
+ hold93/A sky130_fd_sc_hd__o221a_1
X_10272_ curr_PC[7] _10403_/C _10780_/A vssd1 vssd1 vccd1 vccd1 _10272_/Y sky130_fd_sc_hd__a21oi_1
X_12011_ _12012_/A _12012_/B _12012_/C vssd1 vssd1 vccd1 vccd1 _12089_/B sky130_fd_sc_hd__a21o_1
XANTENNA__11067__A _12138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11133__C1 _11126_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12913_ hold27/X hold244/X vssd1 vssd1 vccd1 vccd1 _12913_/X sky130_fd_sc_hd__and2b_1
X_12844_ _12844_/A _12848_/B vssd1 vssd1 vccd1 vccd1 _12844_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_84_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07097__C_N _11470_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12775_ reg1_val[30] _12782_/A vssd1 vssd1 vccd1 vccd1 _12777_/A sky130_fd_sc_hd__or2_1
X_11726_ hold275/A _11636_/B _11808_/B _12247_/C1 vssd1 vssd1 vccd1 vccd1 _11726_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__06608__B _12703_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13221__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12626__A _12626_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11657_ _11655_/B _11657_/B vssd1 vssd1 vccd1 vccd1 _11658_/B sky130_fd_sc_hd__and2b_1
X_11588_ _11589_/A _11589_/B vssd1 vssd1 vccd1 vccd1 _11687_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_4_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10608_ _10608_/A _10608_/B vssd1 vssd1 vccd1 vccd1 _10611_/B sky130_fd_sc_hd__xnor2_2
X_13327_ _13343_/CLK _13327_/D vssd1 vssd1 vccd1 vccd1 hold164/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_506 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07958__A3 _07087_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10539_ fanout94/X _12214_/A fanout51/X _10941_/A vssd1 vssd1 vccd1 vccd1 _10540_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_122_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13258_ _13355_/CLK hold52/X vssd1 vssd1 vccd1 vccd1 hold51/A sky130_fd_sc_hd__dfxtp_1
X_13189_ _13189_/A _13189_/B vssd1 vssd1 vccd1 vccd1 _13189_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_110_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12209_ _12261_/A _12209_/B vssd1 vssd1 vccd1 vccd1 _12210_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07750_ _08728_/A _07750_/B vssd1 vssd1 vccd1 vccd1 _07856_/B sky130_fd_sc_hd__xnor2_2
X_06701_ instruction[0] instruction[1] instruction[2] instruction[26] pred_val vssd1
+ vssd1 vccd1 vccd1 _12629_/B sky130_fd_sc_hd__o311a_4
XANTENNA__13192__A _13214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07681_ _07681_/A _07681_/B vssd1 vssd1 vccd1 vccd1 _08968_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_126_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06632_ reg1_val[25] _07169_/A vssd1 vssd1 vccd1 vccd1 _06633_/B sky130_fd_sc_hd__and2b_1
X_09420_ _09420_/A _09420_/B vssd1 vssd1 vccd1 vccd1 _09463_/A sky130_fd_sc_hd__xnor2_1
X_09351_ _12388_/S _09351_/B vssd1 vssd1 vccd1 vccd1 _09351_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_75_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11978__A1 _06924_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09282_ _09283_/A _09283_/B vssd1 vssd1 vccd1 vccd1 _09282_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_47_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08302_ _10537_/A1 _08671_/B2 _07821_/A _08432_/B vssd1 vssd1 vccd1 vccd1 _08303_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_74_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08233_ _10537_/A1 _07752_/B _07955_/A _08432_/B vssd1 vssd1 vccd1 vccd1 _08234_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08843__A1 _08752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13131__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout228_A _12794_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09399__A2 _07033_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08164_ _11385_/A _08164_/B vssd1 vssd1 vccd1 vccd1 _08166_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10402__A1 _12290_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07115_ _09716_/A _07115_/B vssd1 vssd1 vccd1 vccd1 _07116_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_43_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08095_ _08096_/A _08096_/B vssd1 vssd1 vccd1 vccd1 _08763_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_113_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07046_ _11172_/A _11180_/A _11987_/B vssd1 vssd1 vccd1 vccd1 _07048_/A sky130_fd_sc_hd__nand3b_2
XFILLER_0_30_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10166__B1 _10165_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09571__A2 _10589_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08997_ _08625_/A _08625_/B _08995_/B vssd1 vssd1 vccd1 vccd1 _08997_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__09580__A _10448_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07948_ _07949_/A _07949_/B vssd1 vssd1 vccd1 vccd1 _07948_/Y sky130_fd_sc_hd__nor2_1
X_07879_ _07968_/A _07968_/B _07867_/Y vssd1 vssd1 vccd1 vccd1 _07905_/B sky130_fd_sc_hd__a21boi_2
X_10890_ hold189/A _10890_/B vssd1 vssd1 vccd1 vccd1 _11014_/B sky130_fd_sc_hd__or2_1
X_09618_ _09618_/A _09618_/B _09618_/C _09618_/D vssd1 vssd1 vccd1 vccd1 _09619_/B
+ sky130_fd_sc_hd__or4_1
XANTENNA__08196__A _08722_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09549_ _07052_/Y fanout99/X _10567_/A fanout23/X vssd1 vssd1 vccd1 vccd1 _09550_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_38_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12560_ _12623_/A _12554_/B _12566_/A vssd1 vssd1 vccd1 vccd1 _12561_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_81_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12491_ _12659_/B _12492_/B vssd1 vssd1 vccd1 vccd1 _12502_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_81_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12446__A _12626_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11511_ _11511_/A _11511_/B _11421_/B vssd1 vssd1 vccd1 vccd1 _11702_/A sky130_fd_sc_hd__or3b_2
XFILLER_0_123_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11442_ _11442_/A _11442_/B vssd1 vssd1 vccd1 vccd1 _11442_/X sky130_fd_sc_hd__xor2_1
XANTENNA__08047__C1 _09614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11373_ _12210_/A _11373_/B vssd1 vssd1 vccd1 vccd1 _11377_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_1_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13112_ hold258/X _06892_/B _13111_/X _06572_/A vssd1 vssd1 vccd1 vccd1 hold259/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08062__A2 _08721_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10324_ _10324_/A _10324_/B vssd1 vssd1 vccd1 vccd1 _10326_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_104_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10255_ _13290_/Q _10391_/A2 _10389_/B _12401_/B1 vssd1 vssd1 vccd1 vccd1 _10255_/X
+ sky130_fd_sc_hd__a31o_1
X_13043_ _08584_/A _12798_/B hold143/X vssd1 vssd1 vccd1 vccd1 hold144/A sky130_fd_sc_hd__a21boi_1
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10186_ _10186_/A _10186_/B vssd1 vssd1 vccd1 vccd1 _10187_/B sky130_fd_sc_hd__and2_1
XANTENNA__10413__B _12316_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout290 _06799_/B vssd1 vssd1 vccd1 vccd1 _06771_/A sky130_fd_sc_hd__clkbuf_8
XANTENNA_clkbuf_4_15_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08522__B1 _09440_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12827_ hold17/X _12830_/B _12826_/Y _13245_/A vssd1 vssd1 vccd1 vccd1 hold18/A sky130_fd_sc_hd__o211a_1
XFILLER_0_69_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12758_ _12758_/A _12758_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[26] sky130_fd_sc_hd__nor2_8
XFILLER_0_126_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11709_ _11709_/A _11709_/B vssd1 vssd1 vccd1 vccd1 _11709_/X sky130_fd_sc_hd__xor2_1
X_12689_ _12689_/A _12689_/B _12689_/C vssd1 vssd1 vccd1 vccd1 _12690_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_115_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_450 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout9 fanout9/A vssd1 vssd1 vccd1 vccd1 fanout9/X sky130_fd_sc_hd__buf_6
XANTENNA__08053__A2 fanout87/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12137__A1 _12316_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08920_ _08920_/A _08920_/B vssd1 vssd1 vccd1 vccd1 _08922_/B sky130_fd_sc_hd__xor2_1
XANTENNA__12137__B2 fanout12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08851_ _08826_/A _08826_/B _08824_/Y vssd1 vssd1 vccd1 vccd1 _08859_/A sky130_fd_sc_hd__a21o_1
X_07802_ _07805_/B _07805_/C _07805_/A vssd1 vssd1 vccd1 vccd1 _07807_/A sky130_fd_sc_hd__a21o_1
XANTENNA__10323__B _10324_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08782_ _08783_/A _08783_/B vssd1 vssd1 vccd1 vccd1 _08782_/Y sky130_fd_sc_hd__nand2b_1
X_07733_ _08304_/B fanout99/X _08436_/A fanout75/X vssd1 vssd1 vccd1 vccd1 _07734_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__13126__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07664_ _07664_/A _07664_/B vssd1 vssd1 vccd1 vccd1 _07995_/B sky130_fd_sc_hd__xnor2_1
X_06615_ _06635_/A _12698_/B vssd1 vssd1 vccd1 vccd1 _06615_/Y sky130_fd_sc_hd__nor2_1
X_09403_ _09404_/A _09404_/B _09404_/C _09404_/D vssd1 vssd1 vccd1 vccd1 _09403_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_48_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07595_ _07595_/A _07595_/B vssd1 vssd1 vccd1 vccd1 _07597_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_62_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09334_ _09173_/X _09333_/X _09669_/S vssd1 vssd1 vccd1 vccd1 _09334_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_63_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07619__A2 _11065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09265_ _11146_/A _09396_/B vssd1 vssd1 vccd1 vccd1 _09266_/C sky130_fd_sc_hd__or2_1
XFILLER_0_7_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09196_ fanout23/X _12810_/A _12812_/A _07819_/B vssd1 vssd1 vccd1 vccd1 _09197_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_7_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08216_ _08752_/A _08216_/B vssd1 vssd1 vccd1 vccd1 _08285_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_105_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11179__A2 _11989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08147_ _08148_/A _08148_/B vssd1 vssd1 vccd1 vccd1 _08147_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__12128__A1 _07169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08078_ _08078_/A _08078_/B vssd1 vssd1 vccd1 vccd1 _08891_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_30_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10139__B1 _11142_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07029_ reg1_val[20] reg1_val[21] _07254_/B _12726_/B _07364_/B1 vssd1 vssd1 vccd1
+ vccd1 _07030_/B sky130_fd_sc_hd__o41a_2
XANTENNA__06711__B _06988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07095__A _07095_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10040_ _10040_/A _10040_/B _10040_/C vssd1 vssd1 vccd1 vccd1 _10192_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_11_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold10 hold10/A vssd1 vssd1 vccd1 vccd1 hold10/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 hold21/A vssd1 vssd1 vccd1 vccd1 hold21/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 hold32/A vssd1 vssd1 vccd1 vccd1 hold32/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 hold65/A vssd1 vssd1 vccd1 vccd1 hold65/X sky130_fd_sc_hd__clkbuf_2
Xhold54 hold54/A vssd1 vssd1 vccd1 vccd1 hold54/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 hold43/A vssd1 vssd1 vccd1 vccd1 hold43/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 hold87/A vssd1 vssd1 vccd1 vccd1 hold87/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold98 hold98/A vssd1 vssd1 vccd1 vccd1 hold98/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 hold76/A vssd1 vssd1 vccd1 vccd1 hold76/X sky130_fd_sc_hd__dlygate4sd3_1
X_11991_ _11992_/A _11992_/B _11992_/C vssd1 vssd1 vccd1 vccd1 _11993_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_98_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12300__A1 _12429_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10942_ _07154_/A _07154_/B fanout94/X vssd1 vssd1 vccd1 vccd1 _10943_/C sky130_fd_sc_hd__a21o_1
XANTENNA__12851__A2 _13087_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10873_ _10783_/X _10871_/Y _10872_/Y vssd1 vssd1 vccd1 vccd1 _10873_/Y sky130_fd_sc_hd__a21oi_1
X_12612_ _12612_/A _12612_/B vssd1 vssd1 vccd1 vccd1 _12614_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_39_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12543_ _12544_/A _12544_/B _12544_/C vssd1 vssd1 vccd1 vccd1 _12551_/B sky130_fd_sc_hd__a21o_1
XANTENNA__11811__A0 _09527_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12474_ _12474_/A _12474_/B _12474_/C vssd1 vssd1 vccd1 vccd1 _12475_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_81_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12367__A1 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_7 instruction[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11425_ _10499_/A _10499_/B _10499_/C _10992_/X _11424_/B vssd1 vssd1 vccd1 vccd1
+ _11425_/X sky130_fd_sc_hd__a311o_1
XANTENNA__10917__A2 _12150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11356_ _12448_/S _11353_/X _11354_/Y _11355_/X vssd1 vssd1 vccd1 vccd1 dest_val[16]
+ sky130_fd_sc_hd__a22o_4
XFILLER_0_1_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10307_ _10959_/A _10307_/B vssd1 vssd1 vccd1 vccd1 _10314_/A sky130_fd_sc_hd__xnor2_1
X_13026_ hold95/X _12788_/A _13236_/B hold104/X _13109_/A vssd1 vssd1 vccd1 vccd1
+ hold112/A sky130_fd_sc_hd__o221a_1
X_11287_ _11402_/B _11287_/B vssd1 vssd1 vccd1 vccd1 _11288_/B sky130_fd_sc_hd__or2_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11342__A2 _09527_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10238_ _10141_/X _10275_/C _10237_/Y vssd1 vssd1 vccd1 vccd1 _10270_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_83_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10169_ _10169_/A _10169_/B _10169_/C vssd1 vssd1 vccd1 vccd1 _10172_/B sky130_fd_sc_hd__nand3_1
XANTENNA__06994__D _06994_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08564__A _08673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07380_ _10664_/A _10570_/A _10571_/A _10818_/A vssd1 vssd1 vccd1 vccd1 _07381_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_29_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07482__B1 _12834_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09050_ _09045_/B _09049_/Y _09048_/X vssd1 vssd1 vccd1 vccd1 _09065_/C sky130_fd_sc_hd__o21a_1
XFILLER_0_44_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08001_ _07716_/A _07716_/B _07713_/A vssd1 vssd1 vccd1 vccd1 _08002_/B sky130_fd_sc_hd__a21o_1
XANTENNA__12814__A _12814_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09952_ _09952_/A _09952_/B vssd1 vssd1 vccd1 vccd1 _09956_/B sky130_fd_sc_hd__nor2_1
XANTENNA__07785__B2 _08732_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07785__A1 _08656_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08903_ _08901_/X _08903_/B vssd1 vssd1 vccd1 vccd1 _09056_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_0_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09883_ _09884_/A _09884_/B vssd1 vssd1 vccd1 vccd1 _09883_/Y sky130_fd_sc_hd__nand2_1
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08834_ _08834_/A _08834_/B vssd1 vssd1 vccd1 vccd1 _08835_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__09334__S _09669_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08765_ _08765_/A _08765_/B _08765_/C vssd1 vssd1 vccd1 vccd1 _08766_/B sky130_fd_sc_hd__and3_1
XANTENNA__13086__A2 _06572_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07716_ _07716_/A _07716_/B vssd1 vssd1 vccd1 vccd1 _07718_/B sky130_fd_sc_hd__xor2_1
X_08696_ _08695_/A _08993_/A _08695_/B vssd1 vssd1 vccd1 vccd1 _08995_/B sky130_fd_sc_hd__o21ba_2
XFILLER_0_94_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07647_ _07647_/A _07647_/B vssd1 vssd1 vccd1 vccd1 _07664_/A sky130_fd_sc_hd__xnor2_1
X_07578_ _07579_/A _07579_/B _07579_/C vssd1 vssd1 vccd1 vccd1 _07580_/A sky130_fd_sc_hd__o21a_1
X_09317_ _09313_/X _09316_/X _10248_/S vssd1 vssd1 vccd1 vccd1 _09317_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_63_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06706__B _11343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09248_ _09247_/B _09247_/C _09247_/A vssd1 vssd1 vccd1 vccd1 _09249_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_7_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09179_ _09179_/A _09179_/B vssd1 vssd1 vccd1 vccd1 _09182_/A sky130_fd_sc_hd__nand2_1
X_12190_ _12190_/A _12190_/B vssd1 vssd1 vccd1 vccd1 _12190_/X sky130_fd_sc_hd__or2_1
XFILLER_0_114_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11021__A1 _09354_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11210_ _11210_/A _11210_/B _11210_/C vssd1 vssd1 vccd1 vccd1 _11211_/B sky130_fd_sc_hd__and3_1
XFILLER_0_113_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11141_ _11253_/B _11141_/B vssd1 vssd1 vccd1 vccd1 _11141_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07528__A1 _09768_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11072_ _11072_/A _11072_/B vssd1 vssd1 vccd1 vccd1 _11073_/B sky130_fd_sc_hd__and2_1
XANTENNA__07528__B2 _12808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10023_ _10449_/A _10023_/B vssd1 vssd1 vccd1 vccd1 _10027_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__12809__C1 _13128_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11974_ _11973_/A _09527_/B _11973_/Y _12307_/B1 vssd1 vssd1 vccd1 vccd1 _11974_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__09150__B1 _11886_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07700__A1 _08727_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10925_ _11261_/A _10925_/B vssd1 vssd1 vccd1 vccd1 _10926_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__11803__A _11886_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07700__B2 _08727_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10856_ _10858_/A _10858_/B vssd1 vssd1 vccd1 vccd1 _10859_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_85_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08256__A2 _07821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10787_ _11261_/A _10787_/B vssd1 vssd1 vccd1 vccd1 _10789_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__10419__A _11172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12526_ _12686_/B _12527_/B vssd1 vssd1 vccd1 vccd1 _12537_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_81_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11260__A1 _11653_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11260__B2 _08752_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12457_ _12634_/B _12457_/B vssd1 vssd1 vccd1 vccd1 _12458_/B sky130_fd_sc_hd__or2_1
XFILLER_0_78_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09756__A2 _09567_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11408_ _11408_/A _11408_/B vssd1 vssd1 vccd1 vccd1 _11410_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_105_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12388_ _06859_/Y _12387_/X _12388_/S vssd1 vssd1 vccd1 vccd1 _12389_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_22_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11339_ hold271/A _11339_/B vssd1 vssd1 vccd1 vccd1 _11536_/C sky130_fd_sc_hd__or2_1
XFILLER_0_120_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13009_ _13009_/A hold219/X vssd1 vssd1 vccd1 vccd1 _13307_/D sky130_fd_sc_hd__and2_1
XFILLER_0_94_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06880_ instruction[5] _06880_/B vssd1 vssd1 vccd1 vccd1 dest_pred_val sky130_fd_sc_hd__xnor2_4
XFILLER_0_118_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12815__A2 _12818_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08550_ _09423_/B2 _09238_/B _09440_/B1 _07955_/A vssd1 vssd1 vccd1 vccd1 _08551_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_89_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07501_ _07501_/A _07501_/B vssd1 vssd1 vccd1 vccd1 _07502_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__07152__C1 _06838_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08481_ _08474_/X _08481_/B vssd1 vssd1 vccd1 vccd1 _08518_/B sky130_fd_sc_hd__nand2b_1
X_07432_ _07433_/A _07433_/B vssd1 vssd1 vccd1 vccd1 _07434_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_76_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13240__A2 _06892_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09102_ _09100_/X _09101_/X _09330_/S vssd1 vssd1 vccd1 vccd1 _09102_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_91_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07363_ _07363_/A _07363_/B vssd1 vssd1 vccd1 vccd1 _07378_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_17_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11251__B2 _11876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07294_ _07294_/A _07633_/A _07294_/C vssd1 vssd1 vccd1 vccd1 _07308_/A sky130_fd_sc_hd__and3_1
XFILLER_0_45_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08798__A3 _07087_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout210_A _09441_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09033_ _09033_/A _09036_/B vssd1 vssd1 vccd1 vccd1 _11709_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_4_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12200__B1 _06881_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11554__A2 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09935_ _09724_/A _09724_/B _09725_/Y vssd1 vssd1 vccd1 vccd1 _09940_/A sky130_fd_sc_hd__o21ai_4
XFILLER_0_0_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09866_ _11172_/A _09866_/B vssd1 vssd1 vccd1 vccd1 _09867_/B sky130_fd_sc_hd__xor2_1
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09380__B1 _07282_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08817_ _08817_/A _08817_/B _08817_/C vssd1 vssd1 vccd1 vccd1 _08819_/A sky130_fd_sc_hd__and3_1
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13059__A2 _13087_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09797_ _09798_/A _09798_/B vssd1 vssd1 vccd1 vccd1 _09797_/X sky130_fd_sc_hd__and2b_1
XANTENNA__09132__A0 _09343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08748_ _08748_/A _08748_/B vssd1 vssd1 vccd1 vccd1 _08749_/B sky130_fd_sc_hd__nor2_1
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08679_ _12626_/A _09251_/A _08632_/C _09351_/B vssd1 vssd1 vccd1 vccd1 _09364_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10710_ _10710_/A _10710_/B vssd1 vssd1 vccd1 vccd1 _10712_/B sky130_fd_sc_hd__xnor2_2
XTAP_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11690_ _11691_/A _11691_/B vssd1 vssd1 vccd1 vccd1 _11782_/A sky130_fd_sc_hd__nand2_1
XANTENNA__13231__A2 _12789_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10641_ hold232/A _10641_/B vssd1 vssd1 vccd1 vccd1 _10764_/B sky130_fd_sc_hd__or2_1
XFILLER_0_36_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13360_ _13384_/CLK _13360_/D vssd1 vssd1 vccd1 vccd1 hold282/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10572_ _11269_/A _10572_/B _10572_/C vssd1 vssd1 vccd1 vccd1 _10579_/A sky130_fd_sc_hd__and3_1
X_13291_ _13299_/CLK hold222/X vssd1 vssd1 vccd1 vccd1 hold220/A sky130_fd_sc_hd__dfxtp_1
X_12311_ _12295_/Y _12296_/X _12300_/X _12310_/X vssd1 vssd1 vccd1 vccd1 _12312_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_0_23_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12242_ _12240_/Y _12242_/B vssd1 vssd1 vccd1 vccd1 _12243_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__07548__A _09548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09738__A2 _10167_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07749__B2 _08727_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07749__A1 _08727_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12173_ _12110_/A _12108_/X _12126_/S vssd1 vssd1 vccd1 vccd1 _12176_/B sky130_fd_sc_hd__o21ba_1
XANTENNA__08410__A2 _08744_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11124_ _11452_/B1 _11240_/B hold279/A vssd1 vssd1 vccd1 vccd1 _11126_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_101_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11055_ _11055_/A _11055_/B vssd1 vssd1 vccd1 vccd1 _11056_/B sky130_fd_sc_hd__nor2_1
X_10006_ _10211_/A _10004_/Y _09897_/X _09899_/Y vssd1 vssd1 vccd1 vccd1 _10007_/B
+ sky130_fd_sc_hd__o211a_1
X_11957_ _12174_/S _11956_/X _11955_/X vssd1 vssd1 vccd1 vccd1 _11959_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_59_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08477__A2 _08661_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10908_ _11139_/C _10907_/Y _10780_/A _10905_/X vssd1 vssd1 vccd1 vccd1 dest_val[12]
+ sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_58_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11888_ hold252/A _11888_/B vssd1 vssd1 vccd1 vccd1 _11970_/B sky130_fd_sc_hd__or2_1
XFILLER_0_67_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13222__A2 _12789_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10839_ _10839_/A _10839_/B vssd1 vssd1 vccd1 vccd1 _10852_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12509_ _12509_/A _12509_/B _12509_/C vssd1 vssd1 vccd1 vccd1 _12510_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_14_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout119 _11367_/A vssd1 vssd1 vccd1 vccd1 _10418_/A sky130_fd_sc_hd__buf_6
X_07981_ _07981_/A _07981_/B vssd1 vssd1 vccd1 vccd1 _08022_/A sky130_fd_sc_hd__nand2_2
Xfanout108 _12073_/A vssd1 vssd1 vccd1 vccd1 _11172_/A sky130_fd_sc_hd__buf_6
X_06932_ instruction[24] _12341_/A is_load _06771_/B _06931_/X vssd1 vssd1 vccd1 vccd1
+ _06933_/B sky130_fd_sc_hd__a32o_2
X_09720_ fanout30/X _10413_/A _10567_/A _07688_/B vssd1 vssd1 vccd1 vccd1 _09721_/B
+ sky130_fd_sc_hd__o22a_2
X_06863_ instruction[3] instruction[4] vssd1 vssd1 vccd1 vccd1 _09163_/A sky130_fd_sc_hd__or2_4
X_09651_ _09304_/Y _09648_/Y wire3/X _09075_/B _09650_/Y vssd1 vssd1 vccd1 vccd1 _09652_/B
+ sky130_fd_sc_hd__a221oi_4
XANTENNA__09901__A2 _10571_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06794_ _06596_/A _06695_/A _12639_/B _06792_/X vssd1 vssd1 vccd1 vccd1 _06794_/X
+ sky130_fd_sc_hd__a31o_1
X_08602_ _08673_/A _08741_/A2 _09568_/B _08671_/B2 vssd1 vssd1 vccd1 vccd1 _08603_/B
+ sky130_fd_sc_hd__o22a_1
X_09582_ _11384_/A _09582_/B vssd1 vssd1 vccd1 vccd1 _09584_/B sky130_fd_sc_hd__xnor2_1
X_08533_ _08646_/B2 _09567_/B _08617_/B _09423_/B2 vssd1 vssd1 vccd1 vccd1 _08534_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_77_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07921__A _08740_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11443__A _12244_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout258_A _09442_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08464_ _08467_/A _08467_/B vssd1 vssd1 vccd1 vccd1 _08464_/X sky130_fd_sc_hd__or2_1
XFILLER_0_65_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13213__A2 _13213_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07415_ _09444_/A _10941_/B _12852_/A _09236_/B2 vssd1 vssd1 vccd1 vccd1 _07416_/B
+ sky130_fd_sc_hd__o22a_2
X_08395_ _08739_/A1 _08727_/A2 _08727_/B1 _08436_/A vssd1 vssd1 vccd1 vccd1 _08396_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07428__B1 _12836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07346_ _08436_/B _12852_/A _12854_/A _07149_/A vssd1 vssd1 vccd1 vccd1 _07347_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_73_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08752__A _08752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09016_ _10999_/B _10999_/C vssd1 vssd1 vccd1 vccd1 _11107_/B sky130_fd_sc_hd__and2_1
XANTENNA__09567__B _09567_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07277_ _07278_/A _07278_/B vssd1 vssd1 vccd1 vccd1 _07277_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_5_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold140 hold140/A vssd1 vssd1 vccd1 vccd1 hold140/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold162 hold162/A vssd1 vssd1 vccd1 vccd1 hold162/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold151 hold151/A vssd1 vssd1 vccd1 vccd1 hold151/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07087__B _07087_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold195 hold195/A vssd1 vssd1 vccd1 vccd1 hold195/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold184 hold184/A vssd1 vssd1 vccd1 vccd1 hold184/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 hold173/A vssd1 vssd1 vccd1 vccd1 hold173/X sky130_fd_sc_hd__dlygate4sd3_1
X_09918_ _12804_/A _12316_/B vssd1 vssd1 vccd1 vccd1 _09922_/A sky130_fd_sc_hd__or2_1
X_09849_ _09813_/Y _09848_/X _06881_/X vssd1 vssd1 vccd1 vccd1 _09849_/Y sky130_fd_sc_hd__a21oi_2
X_12860_ _12860_/A _12860_/B vssd1 vssd1 vccd1 vccd1 _13229_/A sky130_fd_sc_hd__nor2_1
XANTENNA__10502__A3 _10500_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11811_ _09527_/B _09354_/B _11811_/S vssd1 vssd1 vccd1 vccd1 _11811_/X sky130_fd_sc_hd__mux2_1
X_12791_ _12791_/A _12791_/B vssd1 vssd1 vccd1 vccd1 _12791_/Y sky130_fd_sc_hd__nand2_1
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12449__A _12629_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11742_ fanout29/X _12150_/A _12213_/A fanout27/X vssd1 vssd1 vccd1 vccd1 _11743_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13204__A2 _13213_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11673_ _11673_/A _11673_/B vssd1 vssd1 vccd1 vccd1 _11675_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_64_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10624_ _10624_/A _10624_/B vssd1 vssd1 vccd1 vccd1 _10624_/X sky130_fd_sc_hd__or2_1
XFILLER_0_48_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13343_ _13343_/CLK _13343_/D vssd1 vssd1 vccd1 vccd1 hold72/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08662__A _08728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10555_ _10418_/A fanout23/X _11171_/A _09745_/B vssd1 vssd1 vccd1 vccd1 _10556_/B
+ sky130_fd_sc_hd__o22a_1
X_13274_ _13285_/CLK hold2/X vssd1 vssd1 vccd1 vccd1 hold1/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10486_ _10487_/B _10487_/A vssd1 vssd1 vccd1 vccd1 _10486_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_121_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12225_ _12092_/Y _12160_/A _12160_/B vssd1 vssd1 vccd1 vccd1 _12334_/A sky130_fd_sc_hd__o21ba_1
XFILLER_0_121_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07198__A2 _07200_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08395__B2 _08436_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08395__A1 _08739_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12156_ _12156_/A _12156_/B _12156_/C vssd1 vssd1 vccd1 vccd1 _12157_/B sky130_fd_sc_hd__nand3_1
X_11107_ _12031_/A _11107_/B _11107_/C vssd1 vssd1 vccd1 vccd1 _11107_/X sky130_fd_sc_hd__or3_1
XANTENNA__10432__A _10928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12087_ _12159_/A _12087_/B vssd1 vssd1 vccd1 vccd1 _12089_/C sky130_fd_sc_hd__nand2_1
XANTENNA__09895__A1 _10941_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11038_ _12073_/A _11038_/B vssd1 vssd1 vccd1 vccd1 _11040_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_91_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09895__B2 _09568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_412 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12989_ _13013_/A hold229/X vssd1 vssd1 vccd1 vccd1 _13297_/D sky130_fd_sc_hd__and2_1
XFILLER_0_115_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07200_ _07200_/A _07200_/B vssd1 vssd1 vccd1 vccd1 _07201_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_55_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08180_ _12818_/A _08732_/A2 _08656_/B _12820_/A vssd1 vssd1 vccd1 vccd1 _08181_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12806__B _12818_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07131_ _07210_/A _07131_/B vssd1 vssd1 vccd1 vccd1 _07133_/D sky130_fd_sc_hd__nand2_1
XFILLER_0_55_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_583 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06804__B _09666_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07188__A _09441_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07062_ _07071_/B _07071_/C vssd1 vssd1 vccd1 vccd1 _11384_/A sky130_fd_sc_hd__nand2_8
XFILLER_0_30_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12822__A _12822_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_754 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07964_ _07964_/A _07964_/B vssd1 vssd1 vccd1 vccd1 _08028_/B sky130_fd_sc_hd__xor2_2
X_06915_ instruction[26] _06921_/B vssd1 vssd1 vccd1 vccd1 _06915_/X sky130_fd_sc_hd__or2_1
X_09703_ _10780_/A _09699_/X _09700_/X _09702_/Y vssd1 vssd1 vccd1 vccd1 dest_val[3]
+ sky130_fd_sc_hd__a22o_4
X_07895_ _07099_/A _07099_/B _07955_/A vssd1 vssd1 vccd1 vccd1 _07897_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_4_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06846_ _06846_/A _06846_/B vssd1 vssd1 vccd1 vccd1 _06846_/Y sky130_fd_sc_hd__nand2_1
X_09634_ _09463_/A _09463_/B _09461_/Y vssd1 vssd1 vccd1 vccd1 _09636_/B sky130_fd_sc_hd__o21a_2
XFILLER_0_4_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07651__A _08731_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06777_ _06775_/Y _06777_/B vssd1 vssd1 vccd1 vccd1 _09964_/A sky130_fd_sc_hd__nand2b_1
X_09565_ _09566_/A _09566_/B vssd1 vssd1 vccd1 vccd1 _09565_/X sky130_fd_sc_hd__and2b_1
X_09496_ _09496_/A vssd1 vssd1 vccd1 vccd1 _09496_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_81_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08516_ _08516_/A vssd1 vssd1 vccd1 vccd1 _08707_/A sky130_fd_sc_hd__inv_2
XFILLER_0_108_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08447_ _08447_/A _08447_/B vssd1 vssd1 vccd1 vccd1 _08492_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_37_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08378_ _08376_/A _08376_/B _08377_/X vssd1 vssd1 vccd1 vccd1 _08424_/A sky130_fd_sc_hd__o21bai_2
XANTENNA__11748__A2 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06714__B _06799_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07329_ _10710_/A _07329_/B vssd1 vssd1 vccd1 vccd1 _07333_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_73_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07098__A _11470_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10340_ _10341_/A _10341_/B vssd1 vssd1 vccd1 vccd1 _10340_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_21_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10271_ curr_PC[7] _10403_/C vssd1 vssd1 vccd1 vccd1 _10271_/X sky130_fd_sc_hd__or2_1
XFILLER_0_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10708__B1 _09568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12010_ _12010_/A _12010_/B vssd1 vssd1 vccd1 vccd1 _12012_/C sky130_fd_sc_hd__or2_1
XANTENNA__13122__B2 _12790_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12912_ hold240/X hold88/X vssd1 vssd1 vccd1 vccd1 _13101_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__09760__B _09761_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12843_ hold19/X _12848_/B _12842_/Y _13214_/A vssd1 vssd1 vccd1 vccd1 hold20/A sky130_fd_sc_hd__o211a_1
XFILLER_0_84_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12774_ _12774_/A _12774_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[29] sky130_fd_sc_hd__xnor2_4
X_11725_ _11636_/B _11808_/B hold275/A vssd1 vssd1 vccd1 vccd1 _11725_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_96_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout90 _07178_/Y vssd1 vssd1 vccd1 vccd1 _12820_/A sky130_fd_sc_hd__buf_8
XANTENNA__12626__B _12626_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11656_ _11770_/A vssd1 vssd1 vccd1 vccd1 _11656_/Y sky130_fd_sc_hd__inv_2
X_11587_ _11472_/A _12214_/B _11557_/A _11476_/A vssd1 vssd1 vccd1 vccd1 _11589_/B
+ sky130_fd_sc_hd__o31ai_2
XFILLER_0_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10427__A _11180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10607_ _10608_/A _10608_/B vssd1 vssd1 vccd1 vccd1 _10607_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_101_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13326_ _13343_/CLK hold136/X vssd1 vssd1 vccd1 vccd1 hold134/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10538_ _10707_/A _10538_/B vssd1 vssd1 vccd1 vccd1 _10542_/A sky130_fd_sc_hd__xnor2_1
X_13257_ _13355_/CLK _13257_/D vssd1 vssd1 vccd1 vccd1 hold90/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12208_ _12316_/A fanout9/X fanout4/X fanout56/X vssd1 vssd1 vccd1 vccd1 _12209_/B
+ sky130_fd_sc_hd__o22a_1
X_10469_ _10469_/A _10469_/B vssd1 vssd1 vccd1 vccd1 _10471_/C sky130_fd_sc_hd__xnor2_1
X_13188_ _12875_/X _13188_/B vssd1 vssd1 vccd1 vccd1 _13189_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__11372__B1 _11923_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12139_ _12139_/A _12412_/A vssd1 vssd1 vccd1 vccd1 _12139_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_19_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06700_ _06698_/X _06700_/B vssd1 vssd1 vccd1 vccd1 _11437_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_126_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07680_ _07678_/A _07678_/B _07679_/Y vssd1 vssd1 vccd1 vccd1 _08968_/A sky130_fd_sc_hd__o21ai_4
X_06631_ _07169_/A reg1_val[25] vssd1 vssd1 vccd1 vccd1 _12126_/S sky130_fd_sc_hd__and2b_1
X_09350_ _09350_/A _09350_/B vssd1 vssd1 vccd1 vccd1 _09350_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09281_ _09281_/A _09281_/B vssd1 vssd1 vccd1 vccd1 _09283_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_74_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08301_ _08301_/A _08301_/B vssd1 vssd1 vccd1 vccd1 _08335_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_74_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08232_ _08235_/A _08235_/B vssd1 vssd1 vccd1 vccd1 _08232_/X sky130_fd_sc_hd__or2_1
XFILLER_0_7_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08843__A2 _09614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout123_A _10927_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08163_ _08798_/B2 fanout69/X _08216_/B _07821_/A vssd1 vssd1 vccd1 vccd1 _08164_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08056__B1 _08564_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07114_ fanout23/X _12802_/A _11171_/A _12804_/A vssd1 vssd1 vccd1 vccd1 _07115_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07803__B1 _12818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08094_ _08745_/A _08094_/B vssd1 vssd1 vccd1 vccd1 _08096_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_101_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07045_ reg1_val[24] _07045_/B vssd1 vssd1 vccd1 vccd1 _11987_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_11_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11363__B1 fanout4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08996_ _08996_/A _08996_/B vssd1 vssd1 vccd1 vccd1 _10503_/B sky130_fd_sc_hd__nor2_1
XANTENNA__10072__A _11180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13104__B2 _06572_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09861__A _12076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07947_ _11384_/A _07947_/B vssd1 vssd1 vccd1 vccd1 _07949_/B sky130_fd_sc_hd__xnor2_1
X_07878_ _07878_/A _07878_/B vssd1 vssd1 vccd1 vccd1 _07968_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_92_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06829_ reg1_val[21] _07135_/D vssd1 vssd1 vccd1 vccd1 _06829_/Y sky130_fd_sc_hd__nand2_1
X_09617_ _09618_/A _09618_/B _09618_/C _09618_/D vssd1 vssd1 vccd1 vccd1 _09617_/X
+ sky130_fd_sc_hd__o22a_1
X_09548_ _09548_/A _09548_/B vssd1 vssd1 vccd1 vccd1 _09552_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout36_A _07282_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09479_ _09480_/A _09480_/B vssd1 vssd1 vccd1 vccd1 _09479_/X sky130_fd_sc_hd__and2_1
XFILLER_0_66_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11510_ _11316_/A _11416_/X _11511_/B vssd1 vssd1 vccd1 vccd1 _11510_/X sky130_fd_sc_hd__a21o_1
X_12490_ reg1_val[7] curr_PC[7] _12622_/S vssd1 vssd1 vccd1 vccd1 _12492_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_80_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11441_ _11439_/Y _11441_/B vssd1 vssd1 vccd1 vccd1 _11442_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_34_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08047__B1 _08752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10929__B1 _10575_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11372_ fanout29/X _11847_/A _11923_/A fanout27/X vssd1 vssd1 vccd1 vccd1 _11373_/B
+ sky130_fd_sc_hd__o22a_1
X_13111_ hold291/A _13110_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13111_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_104_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10323_ _10324_/A _10324_/B vssd1 vssd1 vccd1 vccd1 _10416_/A sky130_fd_sc_hd__or2_1
XFILLER_0_21_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09547__B1 _07263_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10254_ _10391_/A2 _10389_/B _13290_/Q vssd1 vssd1 vccd1 vccd1 _10254_/Y sky130_fd_sc_hd__a21oi_1
X_13042_ hold145/A _12788_/A _13236_/B hold142/X _13109_/A vssd1 vssd1 vccd1 vccd1
+ hold143/A sky130_fd_sc_hd__o221a_1
XFILLER_0_100_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10185_ _10186_/A _10186_/B vssd1 vssd1 vccd1 vccd1 _10187_/A sky130_fd_sc_hd__nor2_1
Xfanout280 hold65/X vssd1 vssd1 vccd1 vccd1 _12790_/A sky130_fd_sc_hd__clkbuf_8
Xfanout291 _06584_/X vssd1 vssd1 vccd1 vccd1 _06799_/B sky130_fd_sc_hd__buf_4
XANTENNA__08522__A1 _12802_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10710__A _10710_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08522__B2 _07896_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12826_ _12826_/A _12830_/B vssd1 vssd1 vccd1 vccd1 _12826_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_69_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12757_ _12766_/A _12766_/B _12757_/C vssd1 vssd1 vccd1 vccd1 _12758_/B sky130_fd_sc_hd__and3_2
XFILLER_0_126_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11708_ _11616_/B _11616_/C _11874_/A vssd1 vssd1 vccd1 vccd1 _11709_/B sky130_fd_sc_hd__o21a_1
X_12688_ _12689_/A _12689_/B _12689_/C vssd1 vssd1 vccd1 vccd1 _12695_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_37_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13031__B1 _09594_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11639_ _11638_/A _09527_/B _11638_/Y _12307_/B1 vssd1 vssd1 vccd1 vccd1 _11639_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_37_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10157__A _12076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13309_ _13314_/CLK hold182/X vssd1 vssd1 vccd1 vccd1 hold223/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07261__A1 _12076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12137__A2 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11345__B1 _11344_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09538__B1 _06881_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08850_ _08817_/A _08817_/C _08817_/B vssd1 vssd1 vccd1 vccd1 _08861_/A sky130_fd_sc_hd__a21bo_2
X_07801_ _07800_/B _07800_/C _08724_/A vssd1 vssd1 vccd1 vccd1 _07805_/C sky130_fd_sc_hd__o21ai_1
XANTENNA__06772__B1 _12429_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08781_ _08211_/A _08211_/B _08209_/X vssd1 vssd1 vccd1 vccd1 _08783_/B sky130_fd_sc_hd__a21o_1
X_07732_ _08740_/A _07732_/B vssd1 vssd1 vccd1 vccd1 _07738_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07663_ _07729_/A _07729_/B vssd1 vssd1 vccd1 vccd1 _07995_/A sky130_fd_sc_hd__nor2_1
X_06614_ instruction[39] _06634_/B vssd1 vssd1 vccd1 vccd1 _12698_/B sky130_fd_sc_hd__and2_4
X_09402_ _09401_/B _09401_/C _11987_/A vssd1 vssd1 vccd1 vccd1 _09404_/D sky130_fd_sc_hd__a21oi_1
X_09333_ _09132_/X _09134_/X _09336_/S vssd1 vssd1 vccd1 vccd1 _09333_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_75_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07594_ _07595_/A _07595_/B vssd1 vssd1 vccd1 vccd1 _09192_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_47_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12547__A _12703_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout240_A _09147_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09264_ _11065_/A _10570_/A vssd1 vssd1 vccd1 vccd1 _09266_/B sky130_fd_sc_hd__or2_1
XFILLER_0_35_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13022__B1 _13213_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09195_ _09548_/A _09195_/B vssd1 vssd1 vccd1 vccd1 _09199_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__10067__A _11261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08215_ _08215_/A _08215_/B vssd1 vssd1 vccd1 vccd1 _08285_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_62_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09777__B1 _10963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08146_ _08146_/A _08146_/B vssd1 vssd1 vccd1 vccd1 _08148_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_120_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08077_ _08075_/B _08872_/B _08075_/A vssd1 vssd1 vccd1 vccd1 _08891_/A sky130_fd_sc_hd__o21ba_1
XFILLER_0_30_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12128__A2 _11343_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07028_ reg1_val[21] _07028_/B vssd1 vssd1 vccd1 vccd1 _07028_/X sky130_fd_sc_hd__xor2_1
XANTENNA__11887__A1 _11886_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold22 hold22/A vssd1 vssd1 vccd1 vccd1 hold22/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold11 hold11/A vssd1 vssd1 vccd1 vccd1 hold11/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07343__A_N _06838_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09591__A _09898_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold44 hold44/A vssd1 vssd1 vccd1 vccd1 hold44/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 hold33/A vssd1 vssd1 vccd1 vccd1 hold33/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 hold55/A vssd1 vssd1 vccd1 vccd1 hold55/X sky130_fd_sc_hd__dlygate4sd3_1
X_08979_ _12423_/A _08980_/B vssd1 vssd1 vccd1 vccd1 _08979_/X sky130_fd_sc_hd__and2_2
Xhold66 hold66/A vssd1 vssd1 vccd1 vccd1 hold66/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 hold88/A vssd1 vssd1 vccd1 vccd1 hold88/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 hold77/A vssd1 vssd1 vccd1 vccd1 hold77/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 hold99/A vssd1 vssd1 vccd1 vccd1 hold99/X sky130_fd_sc_hd__dlygate4sd3_1
X_11990_ _12065_/A _11990_/B vssd1 vssd1 vccd1 vccd1 _11992_/C sky130_fd_sc_hd__xnor2_1
X_10941_ _10941_/A _10941_/B vssd1 vssd1 vccd1 vccd1 _10943_/B sky130_fd_sc_hd__or2_1
XFILLER_0_97_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12611_ _12611_/A _12611_/B vssd1 vssd1 vccd1 vccd1 _12612_/B sky130_fd_sc_hd__nor2_1
X_10872_ _10783_/X _10871_/Y _11707_/A vssd1 vssd1 vccd1 vccd1 _10872_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__12457__A _12634_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12542_ _12551_/A _12542_/B vssd1 vssd1 vccd1 vccd1 _12544_/C sky130_fd_sc_hd__nand2_1
XANTENNA__11811__A1 _09354_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12473_ _12474_/A _12474_/B _12474_/C vssd1 vssd1 vccd1 vccd1 _12481_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_53_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09768__B1 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11424_ _11424_/A _11424_/B vssd1 vssd1 vccd1 vccd1 _11426_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_62_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_8 reg1_val[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08440__B1 _08727_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11355_ curr_PC[16] _11357_/C _11142_/S vssd1 vssd1 vccd1 vccd1 _11355_/X sky130_fd_sc_hd__o21a_1
XANTENNA__07286__A _09442_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11286_ _11285_/B _11286_/B vssd1 vssd1 vccd1 vccd1 _11287_/B sky130_fd_sc_hd__and2b_1
X_10306_ _10567_/A fanout9/X fanout5/X _10413_/A vssd1 vssd1 vccd1 vccd1 _10307_/B
+ sky130_fd_sc_hd__o22a_1
X_13025_ _13242_/A hold96/X vssd1 vssd1 vccd1 vccd1 _13315_/D sky130_fd_sc_hd__and2_1
X_10237_ _10141_/X _10275_/C _12290_/A vssd1 vssd1 vccd1 vccd1 _10237_/Y sky130_fd_sc_hd__a21oi_1
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06710__A_N _06988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10168_ _10449_/A _10168_/B vssd1 vssd1 vccd1 vccd1 _10169_/C sky130_fd_sc_hd__xor2_1
XFILLER_0_83_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10099_ _09482_/X _09645_/X _09646_/X _10368_/A _10496_/A vssd1 vssd1 vccd1 vccd1
+ _10100_/B sky130_fd_sc_hd__a2111oi_2
XFILLER_0_88_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12809_ hold51/X _12856_/B _12808_/Y _13128_/A vssd1 vssd1 vccd1 vccd1 hold52/A sky130_fd_sc_hd__o211a_1
XANTENNA__08564__B _08564_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12055__A1 _11876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10066__B1 fanout66/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07482__A1 _10445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07482__B2 _10706_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08000_ _08000_/A _08000_/B vssd1 vssd1 vccd1 vccd1 _08002_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_4_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12814__B _12818_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08580__A _08728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10615__A _10615_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07196__A _10165_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09951_ _09300_/X _09482_/X _09483_/X _10232_/A _10368_/A vssd1 vssd1 vccd1 vccd1
+ _09952_/B sky130_fd_sc_hd__a2111oi_2
XFILLER_0_40_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07785__A2 _08038_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08902_ _08901_/A _08901_/B _08901_/C vssd1 vssd1 vccd1 vccd1 _08903_/B sky130_fd_sc_hd__a21o_1
XANTENNA__12830__A _12830_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09882_ _08632_/A _08632_/B _12264_/B _09772_/B _09770_/X vssd1 vssd1 vccd1 vccd1
+ _09884_/B sky130_fd_sc_hd__a41o_2
XFILLER_0_57_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout190_A _09127_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06745__B1 _06744_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08833_ _08834_/A _08834_/B vssd1 vssd1 vccd1 vccd1 _08833_/X sky130_fd_sc_hd__or2_1
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08764_ _08765_/A _08765_/B _08765_/C vssd1 vssd1 vccd1 vccd1 _08766_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__08498__B1 _08564_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07715_ _07833_/A _07715_/B vssd1 vssd1 vccd1 vccd1 _07716_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08695_ _08695_/A _08695_/B vssd1 vssd1 vccd1 vccd1 _08993_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_73_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07170__B1 _09440_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07646_ _07642_/A _07642_/B _07991_/A vssd1 vssd1 vccd1 vccd1 _07666_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_48_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07577_ _07577_/A _07577_/B vssd1 vssd1 vccd1 vccd1 _07579_/C sky130_fd_sc_hd__xnor2_1
X_09316_ _09314_/X _09315_/X _09663_/S vssd1 vssd1 vccd1 vccd1 _09316_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_75_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09247_ _09247_/A _09247_/B _09247_/C vssd1 vssd1 vccd1 vccd1 _09379_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_44_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09178_ _11118_/A _09181_/B vssd1 vssd1 vccd1 vccd1 _09179_/B sky130_fd_sc_hd__or2_2
XFILLER_0_90_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09586__A _09906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08129_ _08140_/A vssd1 vssd1 vccd1 vccd1 _08129_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_120_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11140_ curr_PC[13] _11139_/C curr_PC[14] vssd1 vssd1 vccd1 vccd1 _11141_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_31_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07528__A2 fanout23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11071_ _11072_/A _11072_/B vssd1 vssd1 vccd1 vccd1 _11073_/A sky130_fd_sc_hd__nor2_1
X_10022_ _09568_/A _10167_/A1 _10022_/B1 fanout13/X vssd1 vssd1 vccd1 vccd1 _10023_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_98_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11973_ _11973_/A _11973_/B vssd1 vssd1 vccd1 vccd1 _11973_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_58_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10924_ _11653_/A _10571_/B fanout51/X fanout66/X vssd1 vssd1 vccd1 vccd1 _10925_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__13234__B1 _12789_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07700__A2 _11847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10855_ _10987_/B _10855_/B vssd1 vssd1 vccd1 vccd1 _10859_/A sky130_fd_sc_hd__nand2_2
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12525_ reg1_val[12] curr_PC[12] _12586_/S vssd1 vssd1 vccd1 vccd1 _12527_/B sky130_fd_sc_hd__mux2_1
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_384 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10786_ _07087_/A _07087_/B _10570_/B _10571_/B fanout66/X vssd1 vssd1 vccd1 vccd1
+ _10787_/B sky130_fd_sc_hd__o32a_1
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08661__B1 _08673_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11260__A2 _12213_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12456_ _12634_/B _12457_/B vssd1 vssd1 vccd1 vccd1 _12467_/A sky130_fd_sc_hd__nand2_1
X_12387_ _06621_/B _12341_/B _06621_/A vssd1 vssd1 vccd1 vccd1 _12387_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10435__A _10959_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11407_ _11408_/A _11408_/B vssd1 vssd1 vccd1 vccd1 _11504_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__12634__B _12634_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11338_ _11247_/X _11337_/Y _12244_/S vssd1 vssd1 vccd1 vccd1 _11338_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_104_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06632__B _07169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11965__S _12244_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_9_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13355_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11269_ _11269_/A _11269_/B vssd1 vssd1 vccd1 vccd1 _11272_/A sky130_fd_sc_hd__xnor2_1
X_13008_ hold192/X _13016_/A2 _13016_/B1 hold218/X vssd1 vssd1 vccd1 vccd1 hold219/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_94_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06727__B1 _06726_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07500_ _07500_/A _07500_/B vssd1 vssd1 vccd1 vccd1 _07501_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_77_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08480_ _08474_/A _08474_/B _08474_/C vssd1 vssd1 vccd1 vccd1 _08481_/B sky130_fd_sc_hd__a21o_1
X_07431_ _10165_/A _07431_/B vssd1 vssd1 vccd1 vccd1 _07433_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_43_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07362_ _07362_/A _07362_/B vssd1 vssd1 vccd1 vccd1 _07363_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_9_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09101_ reg1_val[14] reg1_val[17] _09108_/S vssd1 vssd1 vccd1 vccd1 _09101_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_72_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07293_ _12138_/A _07293_/B vssd1 vssd1 vccd1 vccd1 _07294_/C sky130_fd_sc_hd__or2_1
X_09032_ _09036_/A _09032_/B vssd1 vssd1 vccd1 vccd1 _11616_/C sky130_fd_sc_hd__xnor2_2
XFILLER_0_32_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07919__A _08742_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold300 hold300/A vssd1 vssd1 vccd1 vccd1 hold300/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07207__A1 _07131_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07207__B2 _07220_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11471__A1_N _07099_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09934_ _09799_/A _09799_/B _09797_/X vssd1 vssd1 vccd1 vccd1 _09941_/A sky130_fd_sc_hd__a21o_1
X_09865_ fanout23/X _10818_/A _10963_/A _11171_/A vssd1 vssd1 vccd1 vccd1 _09866_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07654__A _08728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09380__A1 _12804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09380__B2 _09768_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08816_ _08815_/B _08815_/C _08815_/A vssd1 vssd1 vccd1 vccd1 _08817_/C sky130_fd_sc_hd__o21ai_1
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06733__A3 _12686_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09796_ _09624_/A _09624_/B _09625_/X vssd1 vssd1 vccd1 vccd1 _09798_/B sky130_fd_sc_hd__a21o_1
X_08747_ _08746_/B _08747_/B vssd1 vssd1 vccd1 vccd1 _08748_/B sky130_fd_sc_hd__and2b_1
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08678_ _08678_/A _08678_/B vssd1 vssd1 vccd1 vccd1 _08983_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_68_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07629_ _07629_/A _07629_/B vssd1 vssd1 vccd1 vccd1 _07631_/B sky130_fd_sc_hd__xor2_2
XTAP_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06717__B _06981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10640_ _12244_/S _10638_/X _10639_/Y _09172_/B vssd1 vssd1 vccd1 vccd1 _10640_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_95_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10571_ _10571_/A _10571_/B vssd1 vssd1 vccd1 vccd1 _10572_/C sky130_fd_sc_hd__or2_1
X_12310_ _12305_/Y _12306_/X _12309_/Y _12303_/X vssd1 vssd1 vccd1 vccd1 _12310_/X
+ sky130_fd_sc_hd__o211a_1
X_13290_ _13299_/CLK hold159/X vssd1 vssd1 vccd1 vccd1 _13290_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07829__A _11758_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10450__B1 _10449_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12241_ reg1_val[27] curr_PC[27] vssd1 vssd1 vccd1 vccd1 _12242_/B sky130_fd_sc_hd__nand2_1
XANTENNA__07749__A2 _11847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12172_ _12290_/A _12172_/B _12172_/C vssd1 vssd1 vccd1 vccd1 _12172_/X sky130_fd_sc_hd__or3_1
X_11123_ hold282/A _11123_/B vssd1 vssd1 vccd1 vccd1 _11240_/B sky130_fd_sc_hd__or2_1
XANTENNA__12470__A _12644_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11054_ _11055_/A _11055_/B vssd1 vssd1 vccd1 vccd1 _11056_/A sky130_fd_sc_hd__and2_1
XFILLER_0_64_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10005_ _09897_/X _09899_/Y _10211_/A _10004_/Y vssd1 vssd1 vccd1 vccd1 _10211_/B
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_64_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07382__B1 _10567_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12258__A1 _06882_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11956_ _11880_/A _11877_/X _11894_/A vssd1 vssd1 vccd1 vccd1 _11956_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_86_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10907_ curr_PC[12] _10906_/B _11142_/S vssd1 vssd1 vccd1 vccd1 _10907_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_59_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12629__B _12629_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11887_ _11886_/A _10528_/Y _11886_/Y _06924_/X vssd1 vssd1 vccd1 vccd1 _11887_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_39_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10838_ _10838_/A _10838_/B vssd1 vssd1 vccd1 vccd1 _10839_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10769_ hold269/A _10769_/B vssd1 vssd1 vccd1 vccd1 _10893_/B sky130_fd_sc_hd__or2_1
XFILLER_0_82_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08634__B1 _09442_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12508_ _12509_/A _12509_/B _12509_/C vssd1 vssd1 vccd1 vccd1 _12516_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_81_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12439_ _09108_/S _09147_/X _12433_/Y _12438_/X vssd1 vssd1 vccd1 vccd1 _12439_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_81_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10165__A _10165_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07980_ _07978_/A _07978_/B _07979_/Y vssd1 vssd1 vccd1 vccd1 _08912_/A sky130_fd_sc_hd__a21bo_2
XANTENNA__07070__C1 _11163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout109 _09716_/A vssd1 vssd1 vccd1 vccd1 _12073_/A sky130_fd_sc_hd__buf_8
X_06931_ instruction[40] _06589_/X _06929_/X _06930_/Y vssd1 vssd1 vccd1 vccd1 _06931_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__09362__A1 _09442_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09650_ _09300_/X _09482_/X _09483_/X vssd1 vssd1 vccd1 vccd1 _09650_/Y sky130_fd_sc_hd__a21oi_2
X_06862_ instruction[6] _06861_/Y _06853_/X vssd1 vssd1 vccd1 vccd1 _06862_/Y sky130_fd_sc_hd__a21boi_1
X_08601_ _08627_/A _08627_/B _08601_/C vssd1 vssd1 vccd1 vccd1 _08606_/A sky130_fd_sc_hd__nand3_1
X_06793_ _06805_/A _06695_/A _12639_/B _06792_/X vssd1 vssd1 vccd1 vccd1 _09503_/S
+ sky130_fd_sc_hd__a31oi_4
XANTENNA__06715__A3 _12703_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09581_ _10941_/A _09745_/B _11558_/A fanout94/X vssd1 vssd1 vccd1 vccd1 _09582_/B
+ sky130_fd_sc_hd__o22a_1
X_08532_ _08538_/A _08538_/B vssd1 vssd1 vccd1 vccd1 _08532_/X sky130_fd_sc_hd__and2_1
XFILLER_0_77_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08463_ _08745_/A _08463_/B vssd1 vssd1 vccd1 vccd1 _08467_/B sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout153_A _08722_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07414_ _07460_/B _07414_/B vssd1 vssd1 vccd1 vccd1 _07438_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_107_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08394_ _08394_/A _08394_/B _08394_/C vssd1 vssd1 vccd1 vccd1 _08394_/X sky130_fd_sc_hd__and3_1
XFILLER_0_64_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07428__A1 _10589_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07428__B2 _08507_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07345_ _07345_/A _07345_/B vssd1 vssd1 vccd1 vccd1 _07345_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_0_73_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07276_ _10422_/A _07276_/B vssd1 vssd1 vccd1 vccd1 _07278_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07649__A _08733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08752__B _08752_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09015_ _09015_/A _09015_/B vssd1 vssd1 vccd1 vccd1 _10999_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_103_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold141 hold141/A vssd1 vssd1 vccd1 vccd1 hold141/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold152 hold162/X vssd1 vssd1 vccd1 vccd1 hold152/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold130 hold130/A vssd1 vssd1 vccd1 vccd1 hold130/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold174 hold174/A vssd1 vssd1 vccd1 vccd1 hold174/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold185 hold185/A vssd1 vssd1 vccd1 vccd1 hold185/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold163 hold163/A vssd1 vssd1 vccd1 vccd1 hold163/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12290__A _12290_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold196 hold196/A vssd1 vssd1 vccd1 vccd1 hold196/X sky130_fd_sc_hd__dlygate4sd3_1
X_09917_ _10959_/A _09917_/B _09917_/C vssd1 vssd1 vccd1 vccd1 _09923_/B sky130_fd_sc_hd__or3_1
X_09848_ _09814_/Y _09815_/X _09847_/X vssd1 vssd1 vccd1 vccd1 _09848_/X sky130_fd_sc_hd__o21a_1
XANTENNA_fanout66_A _08752_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09779_ _11146_/A _11653_/A _08752_/B _11294_/A vssd1 vssd1 vccd1 vccd1 _09780_/B
+ sky130_fd_sc_hd__o22a_1
X_11810_ hold252/A _11636_/B _11888_/B _11809_/Y _12247_/C1 vssd1 vssd1 vccd1 vccd1
+ _11810_/X sky130_fd_sc_hd__a311o_1
X_12790_ _12790_/A _12790_/B vssd1 vssd1 vccd1 vccd1 _12790_/Y sky130_fd_sc_hd__nor2_1
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11741_ _12261_/A _11741_/B vssd1 vssd1 vccd1 vccd1 _11745_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__11999__B1 fanout12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10671__B1 _12213_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11672_ fanout27/X _12150_/A _12067_/A fanout29/X vssd1 vssd1 vccd1 vccd1 _11673_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09758__B fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10623_ _10624_/A _10624_/B vssd1 vssd1 vccd1 vccd1 _10623_/Y sky130_fd_sc_hd__nand2_1
X_13342_ _13355_/CLK hold115/X vssd1 vssd1 vccd1 vccd1 hold128/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10554_ _10557_/A vssd1 vssd1 vccd1 vccd1 _10554_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_122_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13273_ _13371_/CLK hold4/X vssd1 vssd1 vccd1 vccd1 hold3/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10485_ _10485_/A _10485_/B vssd1 vssd1 vccd1 vccd1 _10487_/B sky130_fd_sc_hd__xnor2_2
X_12224_ _12222_/Y _12224_/B vssd1 vssd1 vccd1 vccd1 _12414_/A sky130_fd_sc_hd__nand2b_2
XFILLER_0_102_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08395__A2 _08727_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12155_ _12156_/A _12156_/B _12156_/C vssd1 vssd1 vccd1 vccd1 _12157_/A sky130_fd_sc_hd__a21o_1
X_11106_ _11034_/Y _11650_/B _11105_/Y vssd1 vssd1 vccd1 vccd1 _11106_/Y sky130_fd_sc_hd__a21oi_1
X_12086_ _12086_/A _12086_/B vssd1 vssd1 vccd1 vccd1 _12087_/B sky130_fd_sc_hd__or2_1
XANTENNA__09895__A2 _10167_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11037_ _11171_/A fanout48/X _10930_/B fanout23/X vssd1 vssd1 vccd1 vccd1 _11038_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_91_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12988_ hold212/X _13004_/A2 _13006_/B1 hold205/X vssd1 vssd1 vccd1 vccd1 hold229/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11939_ _11939_/A _11939_/B vssd1 vssd1 vccd1 vccd1 _11940_/B sky130_fd_sc_hd__and2_1
XANTENNA__09949__A _09949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10662__B1 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07130_ _07130_/A _11343_/A vssd1 vssd1 vccd1 vccd1 _07133_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_55_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07061_ _07071_/B _07071_/C vssd1 vssd1 vccd1 vccd1 _07485_/A sky130_fd_sc_hd__and2_4
XFILLER_0_2_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09684__A _12341_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12822__B _12830_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09834__D hold260/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07963_ _08076_/A _08076_/B _07953_/X vssd1 vssd1 vccd1 vccd1 _08028_/A sky130_fd_sc_hd__a21o_1
X_06914_ instruction[18] _06884_/Y _06913_/X _06694_/B vssd1 vssd1 vccd1 vccd1 reg2_idx[0]
+ sky130_fd_sc_hd__o211a_4
XANTENNA__07346__B1 _12854_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09702_ _10780_/A _09997_/C vssd1 vssd1 vccd1 vccd1 _09702_/Y sky130_fd_sc_hd__nor2_1
X_07894_ _07902_/A _07902_/B vssd1 vssd1 vccd1 vccd1 _07903_/A sky130_fd_sc_hd__and2_1
X_06845_ _12176_/A _06844_/X _06841_/X vssd1 vssd1 vccd1 vccd1 _06846_/B sky130_fd_sc_hd__a21o_1
X_09633_ _09633_/A _09633_/B vssd1 vssd1 vccd1 vccd1 _09636_/A sky130_fd_sc_hd__nand2_2
XANTENNA__07932__A _08731_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09564_ _09564_/A _09564_/B vssd1 vssd1 vccd1 vccd1 _09566_/B sky130_fd_sc_hd__xor2_2
X_06776_ reg1_val[5] _06960_/C vssd1 vssd1 vccd1 vccd1 _06777_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_78_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08515_ _09010_/A _09010_/B vssd1 vssd1 vccd1 vccd1 _08516_/A sky130_fd_sc_hd__nor2_1
XANTENNA__11445__A2 _09527_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09495_ _11118_/A _09976_/B _09177_/Y vssd1 vssd1 vccd1 vccd1 _09496_/A sky130_fd_sc_hd__a21oi_2
X_08446_ _08474_/A _08446_/B vssd1 vssd1 vccd1 vccd1 _08492_/A sky130_fd_sc_hd__xor2_1
XANTENNA__09859__A _11180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08763__A _11758_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08377_ _08385_/B _08385_/A vssd1 vssd1 vccd1 vccd1 _08377_/X sky130_fd_sc_hd__and2b_1
X_07328_ _10589_/A _12832_/A _12834_/A _08507_/B vssd1 vssd1 vccd1 vccd1 _07329_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_46_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09271__B1 _11987_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07098__B _11470_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07259_ reg1_val[28] _07259_/B vssd1 vssd1 vccd1 vccd1 _07263_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09594__A _09594_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10270_ _10270_/A _10270_/B _10270_/C _10270_/D vssd1 vssd1 vccd1 vccd1 _10270_/X
+ sky130_fd_sc_hd__or4_2
XANTENNA__10708__A1 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10708__B2 _10948_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11905__B1 _12316_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06730__B _07074_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13122__A2 _12789_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12911_ hold88/X hold240/X vssd1 vssd1 vccd1 vccd1 _12911_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_69_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11364__A _12261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12842_ _12842_/A _12848_/B vssd1 vssd1 vccd1 vccd1 _12842_/Y sky130_fd_sc_hd__nand2_1
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12773_ _12773_/A _12773_/B vssd1 vssd1 vccd1 vccd1 _12774_/B sky130_fd_sc_hd__or2_2
X_11724_ hold293/A _11724_/B vssd1 vssd1 vccd1 vccd1 _11808_/B sky130_fd_sc_hd__or2_1
XANTENNA__10644__A0 _09527_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09769__A _12264_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08673__A _08673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11655_ _11657_/B _11655_/B vssd1 vssd1 vccd1 vccd1 _11770_/A sky130_fd_sc_hd__and2b_1
XANTENNA__06905__B _06921_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout80 _12832_/A vssd1 vssd1 vccd1 vccd1 _10574_/B sky130_fd_sc_hd__clkbuf_8
XANTENNA__07289__A _09445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout91 _11564_/A vssd1 vssd1 vccd1 vccd1 _11269_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_0_4_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11586_ _11469_/A _11469_/B _11466_/A vssd1 vssd1 vccd1 vccd1 _11589_/A sky130_fd_sc_hd__a21o_1
X_10606_ _10606_/A _10606_/B vssd1 vssd1 vccd1 vccd1 _10608_/B sky130_fd_sc_hd__xor2_2
X_13325_ _13343_/CLK _13325_/D vssd1 vssd1 vccd1 vccd1 hold150/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10537_ _10537_/A1 _09568_/A fanout13/X _10706_/B2 vssd1 vssd1 vccd1 vccd1 _10538_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_110_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13256_ _13355_/CLK hold36/X vssd1 vssd1 vccd1 vccd1 hold35/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12149__B1 fanout4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10468_ _10469_/A _10469_/B vssd1 vssd1 vccd1 vccd1 _10468_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_122_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12207_ _12317_/A _12207_/B vssd1 vssd1 vccd1 vccd1 _12212_/A sky130_fd_sc_hd__xnor2_1
X_13187_ _13210_/A hold276/X vssd1 vssd1 vccd1 vccd1 _13367_/D sky130_fd_sc_hd__and2_1
X_10399_ _10390_/Y _10391_/X _10398_/Y _10113_/A _10397_/X vssd1 vssd1 vccd1 vccd1
+ _10399_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_86_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11372__B2 fanout27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11372__A1 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12138_ _12138_/A _12138_/B vssd1 vssd1 vccd1 vccd1 _12142_/A sky130_fd_sc_hd__xnor2_1
X_12069_ _11989_/A _12214_/B _12065_/A _11993_/A vssd1 vssd1 vccd1 vccd1 _12084_/A
+ sky130_fd_sc_hd__o31a_1
XANTENNA__07328__B1 _12834_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07752__A _09614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06630_ reg2_val[25] _06771_/A _06703_/B1 _06629_/Y vssd1 vssd1 vccd1 vccd1 _07169_/A
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_126_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06630__A2_N _06771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09280_ _09280_/A _09280_/B vssd1 vssd1 vccd1 vccd1 _09281_/B sky130_fd_sc_hd__xor2_1
X_08300_ _08300_/A _08300_/B vssd1 vssd1 vccd1 vccd1 _08381_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_47_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08231_ _08724_/A _08231_/B vssd1 vssd1 vccd1 vccd1 _08235_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_117_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09253__B1 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08162_ _08752_/A _09396_/B vssd1 vssd1 vccd1 vccd1 _08162_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__08056__B2 _12820_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08056__A1 _12818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07113_ _07113_/A _07113_/B vssd1 vssd1 vccd1 vccd1 _07116_/A sky130_fd_sc_hd__xor2_1
XANTENNA__07803__B2 _08432_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07803__A1 _10537_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08093_ _08436_/A _08744_/A2 _08564_/B fanout99/X vssd1 vssd1 vccd1 vccd1 _08094_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_15_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07044_ _07044_/A _07044_/B vssd1 vssd1 vccd1 vccd1 _09598_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_30_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11363__A1 _11558_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11363__B2 _11472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08995_ _08995_/A _08995_/B vssd1 vssd1 vccd1 vccd1 _08996_/B sky130_fd_sc_hd__xor2_2
XANTENNA__13104__A2 _06892_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07946_ _07896_/A fanout69/X _08216_/B _08723_/B1 vssd1 vssd1 vccd1 vccd1 _07947_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07319__B1 _11171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07662__A _10449_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08758__A _11564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07877_ _07943_/A _07875_/X _07872_/X vssd1 vssd1 vccd1 vccd1 _07968_/A sky130_fd_sc_hd__o21ai_2
X_06828_ reg1_val[22] _07135_/B vssd1 vssd1 vccd1 vccd1 _06828_/Y sky130_fd_sc_hd__nand2_1
X_09616_ _09615_/B _09615_/C _11987_/A vssd1 vssd1 vccd1 vccd1 _09618_/D sky130_fd_sc_hd__a21oi_1
X_06759_ _07080_/A reg1_val[7] vssd1 vssd1 vccd1 vccd1 _06759_/X sky130_fd_sc_hd__and2b_1
X_09547_ _09768_/A1 fanout16/X _07263_/Y _12808_/A vssd1 vssd1 vccd1 vccd1 _09548_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_78_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09478_ _09478_/A _09478_/B vssd1 vssd1 vccd1 vccd1 _09480_/B sky130_fd_sc_hd__xnor2_4
XANTENNA_fanout29_A fanout30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_11_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13380_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_93_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08429_ _08429_/A _08429_/B vssd1 vssd1 vccd1 vccd1 _08451_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_53_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11440_ reg1_val[17] curr_PC[17] vssd1 vssd1 vccd1 vccd1 _11441_/B sky130_fd_sc_hd__nand2_1
XANTENNA__09244__B1 _09593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11371_ _11371_/A _11371_/B vssd1 vssd1 vccd1 vccd1 _11398_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_116_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13110_ _13110_/A _13110_/B vssd1 vssd1 vccd1 vccd1 _13110_/Y sky130_fd_sc_hd__xnor2_1
X_10322_ _10320_/X _10321_/Y _10449_/A vssd1 vssd1 vccd1 vccd1 _10324_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_34_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13041_ _07217_/B _12798_/B hold146/X vssd1 vssd1 vccd1 vccd1 hold147/A sky130_fd_sc_hd__a21boi_1
XANTENNA__09547__A1 _09768_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10253_ hold157/A _10253_/B vssd1 vssd1 vccd1 vccd1 _10389_/B sky130_fd_sc_hd__or2_1
XANTENNA__09547__B2 _12808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10184_ _11384_/A _10184_/B vssd1 vssd1 vccd1 vccd1 _10186_/B sky130_fd_sc_hd__xnor2_1
Xfanout270 _06686_/A vssd1 vssd1 vccd1 vccd1 _06702_/A sky130_fd_sc_hd__clkbuf_8
Xfanout292 _06596_/A vssd1 vssd1 vccd1 vccd1 _06805_/A sky130_fd_sc_hd__buf_6
Xfanout281 _07200_/A vssd1 vssd1 vccd1 vccd1 _07364_/B1 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_88_327 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08522__A2 _09238_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12825_ hold13/X _12818_/B _12824_/Y _13245_/A vssd1 vssd1 vccd1 vccd1 hold14/A sky130_fd_sc_hd__o211a_1
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12756_ _12766_/B _12757_/C _12766_/A vssd1 vssd1 vccd1 vccd1 _12758_/A sky130_fd_sc_hd__a21oi_4
XANTENNA__06635__B _12680_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11707_ _11707_/A _11707_/B vssd1 vssd1 vccd1 vccd1 _11707_/Y sky130_fd_sc_hd__nand2_1
X_12687_ _12687_/A _12695_/A vssd1 vssd1 vccd1 vccd1 _12689_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_21_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11638_ _11638_/A _11973_/B vssd1 vssd1 vccd1 vccd1 _11638_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_71_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13308_ _13314_/CLK hold209/X vssd1 vssd1 vccd1 vccd1 hold207/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11569_ _11569_/A _11569_/B vssd1 vssd1 vccd1 vccd1 _11570_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_12_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07261__A2 _07263_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11345__A1 _09167_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13239_ hold172/X hold63/X _13109_/A _13238_/X vssd1 vssd1 vccd1 vccd1 hold64/A sky130_fd_sc_hd__o211a_1
XFILLER_0_20_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11269__A _11269_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11896__A2 _11343_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07800_ _08724_/A _07800_/B _07800_/C vssd1 vssd1 vccd1 vccd1 _07805_/B sky130_fd_sc_hd__or3_1
X_08780_ _08780_/A _08780_/B vssd1 vssd1 vccd1 vccd1 _08783_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__09173__S _09351_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07731_ _08741_/B2 fanout87/X fanout82/X _08732_/A1 vssd1 vssd1 vccd1 vccd1 _07732_/B
+ sky130_fd_sc_hd__o22a_1
X_07662_ _10449_/A _07662_/B vssd1 vssd1 vccd1 vccd1 _07729_/B sky130_fd_sc_hd__xnor2_1
X_06613_ _12402_/S _06613_/B vssd1 vssd1 vccd1 vccd1 _12389_/A sky130_fd_sc_hd__nor2_2
X_07593_ _07593_/A _07593_/B vssd1 vssd1 vccd1 vccd1 _07595_/B sky130_fd_sc_hd__xnor2_2
X_09401_ _11987_/A _09401_/B _09401_/C vssd1 vssd1 vccd1 vccd1 _09404_/C sky130_fd_sc_hd__and3_1
XANTENNA__12828__A _12828_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09332_ _09328_/X _09970_/B _09974_/A vssd1 vssd1 vccd1 vccd1 _09332_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_118_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09263_ _07449_/A _07449_/B _07446_/A vssd1 vssd1 vccd1 vccd1 _09281_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__09202__A _11673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09194_ _12802_/A fanout16/X _07282_/B _12804_/A vssd1 vssd1 vccd1 vccd1 _09195_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_62_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09226__B1 _12836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08214_ _08214_/A _08214_/B vssd1 vssd1 vccd1 vccd1 _08249_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_28_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09777__B2 _09613_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09777__A1 _11065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08145_ _08169_/A _08169_/B vssd1 vssd1 vccd1 vccd1 _08148_/A sky130_fd_sc_hd__or2_1
X_08076_ _08076_/A _08076_/B vssd1 vssd1 vccd1 vccd1 _08872_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_30_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07027_ reg1_val[20] _07254_/B _12726_/B _07364_/B1 vssd1 vssd1 vccd1 vccd1 _07028_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_3_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold23 hold23/A vssd1 vssd1 vccd1 vccd1 hold23/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold12 hold12/A vssd1 vssd1 vccd1 vccd1 hold12/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 hold45/A vssd1 vssd1 vccd1 vccd1 hold45/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 hold34/A vssd1 vssd1 vccd1 vccd1 hold34/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 hold56/A vssd1 vssd1 vccd1 vccd1 hold56/X sky130_fd_sc_hd__dlygate4sd3_1
X_08978_ _09706_/A _08978_/B vssd1 vssd1 vccd1 vccd1 _09542_/A sky130_fd_sc_hd__xor2_2
Xhold89 hold89/A vssd1 vssd1 vccd1 vccd1 hold89/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11639__A2 _09527_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold67 hold67/A vssd1 vssd1 vccd1 vccd1 hold67/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 hold78/A vssd1 vssd1 vccd1 vccd1 hold78/X sky130_fd_sc_hd__dlygate4sd3_1
X_07929_ _11908_/A _07929_/B vssd1 vssd1 vccd1 vccd1 _07940_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_97_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10940_ _11076_/B _10940_/B vssd1 vssd1 vccd1 vccd1 _10954_/A sky130_fd_sc_hd__nor2_1
X_12610_ _12611_/A _12611_/B vssd1 vssd1 vccd1 vccd1 _12612_/A sky130_fd_sc_hd__and2_1
X_10871_ _10871_/A _10871_/B vssd1 vssd1 vccd1 vccd1 _10871_/Y sky130_fd_sc_hd__nand2_2
X_12541_ _12698_/B _12541_/B vssd1 vssd1 vccd1 vccd1 _12542_/B sky130_fd_sc_hd__or2_1
XFILLER_0_93_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09217__B1 _09568_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12472_ _12481_/A _12472_/B vssd1 vssd1 vccd1 vccd1 _12474_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_19_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09768__B2 _07026_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09768__A1 _09768_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11423_ _11423_/A _11608_/A vssd1 vssd1 vccd1 vccd1 _11424_/B sky130_fd_sc_hd__or2_1
XFILLER_0_123_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09766__B _12316_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_9 reg1_val[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08440__B2 _08739_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08440__A1 _08721_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11354_ curr_PC[16] _11357_/C vssd1 vssd1 vccd1 vccd1 _11354_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11285_ _11286_/B _11285_/B vssd1 vssd1 vccd1 vccd1 _11402_/B sky130_fd_sc_hd__and2b_1
X_10305_ _10480_/B _10305_/B vssd1 vssd1 vccd1 vccd1 _10344_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_21_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13024_ hold95/X _06892_/B _12798_/B reg1_val[0] vssd1 vssd1 vccd1 vccd1 hold96/A
+ sky130_fd_sc_hd__a22o_1
X_10236_ _10741_/A _10236_/B vssd1 vssd1 vccd1 vccd1 _10275_/C sky130_fd_sc_hd__xnor2_4
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10167_ _10167_/A1 fanout13/X fanout6/X _07222_/Y vssd1 vssd1 vccd1 vccd1 _10168_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_89_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10098_ _09806_/X _09947_/X _09948_/X vssd1 vssd1 vccd1 vccd1 _10100_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_89_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12808_ _12808_/A _12856_/B vssd1 vssd1 vccd1 vccd1 _12808_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_57_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10066__A1 _10418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11271__B fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10168__A _10449_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12739_ _12746_/C _12739_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[22] sky130_fd_sc_hd__xnor2_4
XANTENNA__10066__B2 _09745_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07482__A2 _12832_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09759__B2 _09897_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09950_ _09645_/X _09806_/X _09807_/X vssd1 vssd1 vccd1 vccd1 _09952_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__07785__A3 _08038_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08901_ _08901_/A _08901_/B _08901_/C vssd1 vssd1 vccd1 vccd1 _08901_/X sky130_fd_sc_hd__and3_1
XFILLER_0_0_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12830__B _12830_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09881_ _09881_/A _09881_/B vssd1 vssd1 vccd1 vccd1 _09884_/A sky130_fd_sc_hd__xor2_4
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08195__B1 _07955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08832_ _08834_/A _08834_/B vssd1 vssd1 vccd1 vccd1 _08832_/X sky130_fd_sc_hd__and2_1
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08763_ _11758_/A _08763_/B vssd1 vssd1 vccd1 vccd1 _08765_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__08498__A1 _08798_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07714_ _10148_/A _09609_/B _09396_/B _07089_/Y vssd1 vssd1 vccd1 vccd1 _07715_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08498__B2 _08646_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08694_ _08653_/A _08653_/B _08693_/X vssd1 vssd1 vccd1 vccd1 _08993_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_79_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07170__A1 _09238_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07170__B2 _12844_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07645_ _07990_/A _07990_/B vssd1 vssd1 vccd1 vccd1 _07991_/A sky130_fd_sc_hd__and2_1
XANTENNA__13243__B2 _06572_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07576_ _07363_/A _07363_/B _07361_/X vssd1 vssd1 vccd1 vccd1 _07581_/A sky130_fd_sc_hd__o21ai_4
XANTENNA__09447__B1 _10930_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09315_ _09093_/X _09095_/X _09330_/S vssd1 vssd1 vccd1 vccd1 _09315_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_48_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09246_ _09245_/A _09245_/B _09237_/Y vssd1 vssd1 vccd1 vccd1 _09247_/C sky130_fd_sc_hd__o21bai_1
XFILLER_0_105_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09177_ _11118_/A _09181_/B vssd1 vssd1 vccd1 vccd1 _09177_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_50_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10806__A _11180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07225__A2 _07220_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08128_ _08728_/A _08128_/B vssd1 vssd1 vccd1 vccd1 _08140_/A sky130_fd_sc_hd__xnor2_2
X_08059_ _08055_/A _08055_/B _08808_/A vssd1 vssd1 vccd1 vccd1 _08067_/A sky130_fd_sc_hd__o21ba_2
XANTENNA_fanout96_A _12818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11070_ _11070_/A _11070_/B vssd1 vssd1 vccd1 vccd1 _11072_/B sky130_fd_sc_hd__xnor2_1
X_10021_ _10021_/A _10021_/B vssd1 vssd1 vccd1 vccd1 _10029_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_11_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07933__B1 _08656_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11972_ hold265/A _11636_/B _12046_/B _12247_/C1 vssd1 vssd1 vccd1 vccd1 _11972_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_98_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10923_ _10923_/A _10923_/B vssd1 vssd1 vccd1 vccd1 _10926_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_128_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10854_ _10854_/A _10854_/B _10854_/C vssd1 vssd1 vccd1 vccd1 _10855_/B sky130_fd_sc_hd__or3_1
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12524_ _12530_/B _12524_/B vssd1 vssd1 vccd1 vccd1 new_PC[11] sky130_fd_sc_hd__and2_4
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10785_ _11470_/A _10785_/B vssd1 vssd1 vccd1 vccd1 _10789_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12915__B hold260/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08681__A _08681_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08661__A1 _08673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08661__B2 _08671_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06913__B _06921_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12455_ reg1_val[2] curr_PC[2] _12455_/S vssd1 vssd1 vccd1 vccd1 _12457_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_81_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12386_ _12382_/Y _12384_/X _12385_/Y vssd1 vssd1 vccd1 vccd1 _12386_/X sky130_fd_sc_hd__o21a_1
X_11406_ _11301_/A _11301_/B _11304_/A vssd1 vssd1 vccd1 vccd1 _11408_/B sky130_fd_sc_hd__a21bo_1
X_11337_ _11337_/A _11337_/B vssd1 vssd1 vccd1 vccd1 _11337_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_22_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10508__C1 _11624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11268_ _10570_/A _12316_/A fanout12/X _10571_/A vssd1 vssd1 vccd1 vccd1 _11269_/B
+ sky130_fd_sc_hd__o22a_1
X_13007_ _13013_/A hold193/X vssd1 vssd1 vccd1 vccd1 hold194/A sky130_fd_sc_hd__and2_1
X_10219_ _10218_/A _10218_/B _10220_/A vssd1 vssd1 vccd1 vccd1 _10219_/X sky130_fd_sc_hd__a21bo_1
X_11199_ _11086_/A _11086_/B _11084_/X vssd1 vssd1 vccd1 vccd1 _11201_/B sky130_fd_sc_hd__a21bo_1
XANTENNA__07924__B1 _08564_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07152__A1 _07144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11484__B1 _11923_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07430_ _12842_/A _09567_/B _09568_/B _12844_/A vssd1 vssd1 vccd1 vccd1 _07431_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_76_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07361_ _07362_/A _07362_/B vssd1 vssd1 vccd1 vccd1 _07361_/X sky130_fd_sc_hd__or2_1
XFILLER_0_43_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09100_ reg1_val[15] reg1_val[16] _09108_/S vssd1 vssd1 vccd1 vccd1 _09100_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_72_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08101__B1 _08656_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07292_ _07292_/A _07292_/B _07293_/B vssd1 vssd1 vccd1 vccd1 _07633_/A sky130_fd_sc_hd__or3b_1
X_09031_ _08344_/A _09026_/A _09026_/B _09030_/X vssd1 vssd1 vccd1 vccd1 _09032_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_5_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold301 hold301/A vssd1 vssd1 vccd1 vccd1 hold70/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09933_ _09791_/A _09790_/B _09788_/Y vssd1 vssd1 vccd1 vccd1 _09943_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_110_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09864_ _09864_/A _09864_/B vssd1 vssd1 vccd1 vccd1 _09867_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09380__A2 fanout16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08815_ _08815_/A _08815_/B _08815_/C vssd1 vssd1 vccd1 vccd1 _08817_/B sky130_fd_sc_hd__or3_1
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09795_ _09607_/A _09607_/B _09605_/X vssd1 vssd1 vccd1 vccd1 _09798_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_68_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08746_ _08747_/B _08746_/B vssd1 vssd1 vccd1 vccd1 _08748_/A sky130_fd_sc_hd__and2b_1
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07143__A1 _07144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08677_ _08678_/A _08677_/B _08677_/C vssd1 vssd1 vccd1 vccd1 _08677_/X sky130_fd_sc_hd__and3_1
XFILLER_0_68_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07628_ _07628_/A _07628_/B vssd1 vssd1 vccd1 vccd1 _07631_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_67_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07559_ _07557_/Y _07559_/B vssd1 vssd1 vccd1 vccd1 _07560_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_119_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10570_ _10570_/A _10570_/B vssd1 vssd1 vccd1 vccd1 _10572_/B sky130_fd_sc_hd__or2_1
XFILLER_0_17_750 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09229_ _11385_/A _09229_/B vssd1 vssd1 vccd1 vccd1 _09231_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_17_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12240_ reg1_val[27] curr_PC[27] vssd1 vssd1 vccd1 vccd1 _12240_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_16_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12171_ _12170_/A _12287_/A _12170_/B vssd1 vssd1 vccd1 vccd1 _12172_/C sky130_fd_sc_hd__a21oi_1
XFILLER_0_31_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11122_ _11886_/A _11117_/X _11121_/Y _09172_/B vssd1 vssd1 vccd1 vccd1 _11137_/B
+ sky130_fd_sc_hd__o211a_1
XANTENNA__11367__A _11367_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11053_ _11180_/A _11053_/B vssd1 vssd1 vccd1 vccd1 _11055_/B sky130_fd_sc_hd__xnor2_1
X_10004_ _07035_/Y _12264_/B _09907_/Y _09911_/A vssd1 vssd1 vccd1 vccd1 _10004_/Y
+ sky130_fd_sc_hd__a211oi_1
XANTENNA__07382__B2 fanout66/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07382__A1 _11653_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10269__A1 _09111_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11955_ _11880_/A _11878_/X _06828_/Y _12423_/A vssd1 vssd1 vccd1 vccd1 _11955_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_59_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10906_ curr_PC[12] _10906_/B vssd1 vssd1 vccd1 vccd1 _11139_/C sky130_fd_sc_hd__and2_1
XFILLER_0_104_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11886_ _11886_/A _11886_/B vssd1 vssd1 vccd1 vccd1 _11886_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_73_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12966__B1 _13213_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10837_ _10838_/A _10838_/B vssd1 vssd1 vccd1 vccd1 _10976_/B sky130_fd_sc_hd__nand2_1
X_10768_ _12307_/B1 _10767_/X _06737_/B vssd1 vssd1 vccd1 vccd1 _10768_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_109_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12507_ _12516_/A _12507_/B vssd1 vssd1 vccd1 vccd1 _12509_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_125_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12438_ _08980_/B _09158_/Y _12430_/A _09152_/Y _12437_/X vssd1 vssd1 vccd1 vccd1
+ _12438_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_54_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10699_ _10700_/A _10700_/B vssd1 vssd1 vccd1 vccd1 _10699_/X sky130_fd_sc_hd__and2_1
XFILLER_0_2_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12369_ fanout13/X _12316_/B _12366_/Y _12418_/S vssd1 vssd1 vccd1 vccd1 _12372_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_2_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06930_ instruction[6] is_load vssd1 vssd1 vccd1 vccd1 _06930_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__11277__A _12317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06861_ _08980_/B _12423_/B _06852_/Y vssd1 vssd1 vccd1 vccd1 _06861_/Y sky130_fd_sc_hd__o21ai_1
X_08600_ _09897_/A _08600_/B vssd1 vssd1 vccd1 vccd1 _08601_/C sky130_fd_sc_hd__xnor2_1
X_06792_ reg2_val[2] _06799_/B vssd1 vssd1 vccd1 vccd1 _06792_/X sky130_fd_sc_hd__and2_2
X_09580_ _10448_/A _09580_/B vssd1 vssd1 vccd1 vccd1 _09584_/A sky130_fd_sc_hd__xnor2_1
X_08531_ _08560_/A _08529_/Y _08526_/Y vssd1 vssd1 vccd1 vccd1 _08538_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_89_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08462_ _08646_/B2 _08744_/A2 _08564_/B _09423_/B2 vssd1 vssd1 vccd1 vccd1 _08463_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_54_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07413_ _07413_/A _07413_/B vssd1 vssd1 vccd1 vccd1 _07414_/B sky130_fd_sc_hd__nand2_1
XANTENNA__12836__A _12836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08393_ _08645_/A _08393_/B _08393_/C vssd1 vssd1 vccd1 vccd1 _08394_/C sky130_fd_sc_hd__or3_1
XANTENNA_fanout146_A _07036_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07428__A2 _12834_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07344_ _07142_/Y _07343_/Y _07220_/B vssd1 vssd1 vccd1 vccd1 _07345_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_73_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07275_ _11653_/A _12810_/A fanout66/X _10413_/A vssd1 vssd1 vccd1 vccd1 _07276_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_72_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09014_ _09013_/A _09013_/B _09015_/A vssd1 vssd1 vccd1 vccd1 _09014_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_0_41_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold120 hold120/A vssd1 vssd1 vccd1 vccd1 hold120/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold142 hold142/A vssd1 vssd1 vccd1 vccd1 hold142/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold153 hold153/A vssd1 vssd1 vccd1 vccd1 hold153/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold131 hold131/A vssd1 vssd1 vccd1 vccd1 hold131/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold175 hold175/A vssd1 vssd1 vccd1 vccd1 hold175/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold186 hold186/A vssd1 vssd1 vccd1 vccd1 hold186/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold164 hold164/A vssd1 vssd1 vccd1 vccd1 hold164/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold197 hold234/X vssd1 vssd1 vccd1 vccd1 hold197/X sky130_fd_sc_hd__dlygate4sd3_1
X_09916_ _09917_/B _09917_/C _10959_/A vssd1 vssd1 vccd1 vccd1 _09923_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__09880__A _11269_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09847_ _10113_/A _09821_/X _09846_/X _09819_/Y vssd1 vssd1 vccd1 vccd1 _09847_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold260_A hold260/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09778_ _11180_/A _09778_/B vssd1 vssd1 vccd1 vccd1 _09782_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__09091__S _09666_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout59_A _12848_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08729_ _08736_/A vssd1 vssd1 vccd1 vccd1 _08729_/Y sky130_fd_sc_hd__inv_2
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11740_ _11923_/A fanout9/X fanout4/X _11847_/A vssd1 vssd1 vccd1 vccd1 _11741_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11999__B2 fanout27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11999__A1 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10671__B2 fanout94/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10671__A1 _10941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11671_ _11768_/A _11671_/B vssd1 vssd1 vccd1 vccd1 _11675_/A sky130_fd_sc_hd__or2_1
XFILLER_0_63_130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10622_ _11102_/A _10622_/B vssd1 vssd1 vccd1 vccd1 _10624_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_36_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13341_ _13355_/CLK hold69/X vssd1 vssd1 vccd1 vccd1 _13341_/Q sky130_fd_sc_hd__dfxtp_1
X_10553_ _10928_/A _10553_/B vssd1 vssd1 vccd1 vccd1 _10557_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_8_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13272_ _13371_/CLK hold10/X vssd1 vssd1 vccd1 vccd1 hold9/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11796__S _12423_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10484_ _10484_/A _10484_/B vssd1 vssd1 vccd1 vccd1 _10485_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_122_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12223_ _12277_/B _12221_/X _12154_/A _12157_/A vssd1 vssd1 vccd1 vccd1 _12224_/B
+ sky130_fd_sc_hd__o211ai_2
X_12154_ _12154_/A _12154_/B vssd1 vssd1 vccd1 vccd1 _12156_/C sky130_fd_sc_hd__nand2_1
X_11105_ _11034_/Y _11650_/B _11707_/A vssd1 vssd1 vccd1 vccd1 _11105_/Y sky130_fd_sc_hd__o21ai_1
X_12085_ _12086_/A _12086_/B vssd1 vssd1 vccd1 vccd1 _12159_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08552__B1 _08038_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11036_ _12210_/A _11036_/B vssd1 vssd1 vccd1 vccd1 _11040_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__06746__A_N _07095_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12987_ _13013_/A hold213/X vssd1 vssd1 vccd1 vccd1 hold214/A sky130_fd_sc_hd__and2_1
XANTENNA__06638__B _07140_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11938_ _11939_/A _11939_/B vssd1 vssd1 vccd1 vccd1 _11940_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_86_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09949__B _09949_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11869_ _11517_/B _11868_/Y _11867_/Y vssd1 vssd1 vccd1 vccd1 _11870_/B sky130_fd_sc_hd__a21oi_2
XANTENNA__10662__B2 _11146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10662__A1 _11065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10414__A1 _10413_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07060_ reg1_val[16] _07364_/B1 _07069_/B reg1_val[17] vssd1 vssd1 vccd1 vccd1 _07071_/C
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_27_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_30 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07485__A _07485_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10623__B _10624_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09701_ curr_PC[3] _09701_/B vssd1 vssd1 vccd1 vccd1 _09997_/C sky130_fd_sc_hd__and2_1
X_07962_ _07962_/A _07962_/B vssd1 vssd1 vccd1 vccd1 _08076_/B sky130_fd_sc_hd__xnor2_2
X_06913_ instruction[25] _06921_/B vssd1 vssd1 vccd1 vccd1 _06913_/X sky130_fd_sc_hd__or2_1
XANTENNA__07346__A1 _08436_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07893_ _07890_/B _07915_/B _07890_/A vssd1 vssd1 vccd1 vccd1 _07902_/B sky130_fd_sc_hd__o21bai_1
XANTENNA__07346__B2 _07149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06844_ _12110_/A _06843_/X _06842_/X vssd1 vssd1 vccd1 vccd1 _06844_/X sky130_fd_sc_hd__a21o_1
X_09632_ _09391_/A _09391_/B _09392_/Y vssd1 vssd1 vccd1 vccd1 _09637_/A sky130_fd_sc_hd__o21ai_4
XFILLER_0_78_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09563_ _09405_/B _09408_/B _09403_/X vssd1 vssd1 vccd1 vccd1 _09564_/B sky130_fd_sc_hd__a21o_1
X_06775_ reg1_val[5] _06960_/C vssd1 vssd1 vccd1 vccd1 _06775_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_fanout263_A _12455_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08514_ _08514_/A _08514_/B vssd1 vssd1 vccd1 vccd1 _09010_/B sky130_fd_sc_hd__xnor2_1
X_09494_ _10250_/S _09334_/X _09176_/B vssd1 vssd1 vccd1 vccd1 _09976_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__10653__A1 _09152_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08445_ _08474_/A _08446_/B vssd1 vssd1 vccd1 vccd1 _08445_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_105_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08376_ _08376_/A _08376_/B vssd1 vssd1 vccd1 vccd1 _08385_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_46_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11470__A _11470_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07327_ _07325_/A _07325_/B _07326_/X vssd1 vssd1 vccd1 vccd1 _07394_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_45_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07258_ _07254_/B _07254_/C _12765_/B _07364_/B1 vssd1 vssd1 vccd1 vccd1 _07259_/B
+ sky130_fd_sc_hd__o31a_2
XFILLER_0_5_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07189_ _09433_/A _10024_/A _07187_/Y vssd1 vssd1 vccd1 vccd1 _07189_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_103_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09086__S _09108_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10708__A2 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11905__B2 fanout27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11905__A1 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12910_ _12908_/X _12910_/B vssd1 vssd1 vccd1 vccd1 _13106_/A sky130_fd_sc_hd__nand2b_1
X_12841_ hold1/X _12848_/B _12840_/Y _13210_/A vssd1 vssd1 vccd1 vccd1 hold2/A sky130_fd_sc_hd__o211a_1
XFILLER_0_69_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12772_ _12772_/A _12772_/B vssd1 vssd1 vccd1 vccd1 _12774_/A sky130_fd_sc_hd__nand2_2
X_11723_ _11723_/A _11723_/B vssd1 vssd1 vccd1 vccd1 _11723_/X sky130_fd_sc_hd__or2_1
XANTENNA__10644__A1 _09354_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08673__B _08673_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11380__A _12073_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11654_ _11758_/A _11654_/B vssd1 vssd1 vccd1 vccd1 _11655_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_92_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout81 _07210_/Y vssd1 vssd1 vccd1 vccd1 _12832_/A sky130_fd_sc_hd__buf_4
XFILLER_0_64_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout92 _07833_/A vssd1 vssd1 vccd1 vccd1 _11564_/A sky130_fd_sc_hd__buf_8
Xfanout70 _07819_/B vssd1 vssd1 vccd1 vccd1 _11171_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_37_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10605_ _10484_/A _10484_/B _10482_/X vssd1 vssd1 vccd1 vccd1 _10606_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_52_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11585_ _11486_/A _11486_/B _11487_/X vssd1 vssd1 vccd1 vccd1 _11591_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_24_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13324_ _13343_/CLK hold144/X vssd1 vssd1 vccd1 vccd1 hold142/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07273__B1 _08216_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12149__A1 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10536_ _10416_/A _10415_/B _10415_/A vssd1 vssd1 vccd1 vccd1 _10551_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_122_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13255_ _13355_/CLK hold50/X vssd1 vssd1 vccd1 vccd1 hold49/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12149__B2 _12213_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10467_ _11470_/A _10467_/B vssd1 vssd1 vccd1 vccd1 _10469_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__06921__B _06921_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12206_ fanout16/X fanout12/X fanout8/X _07282_/B vssd1 vssd1 vccd1 vccd1 _12207_/B
+ sky130_fd_sc_hd__o22a_1
X_13186_ hold275/X _13213_/A2 _13185_/X _13213_/B2 vssd1 vssd1 vccd1 vccd1 hold276/A
+ sky130_fd_sc_hd__a22o_1
X_10398_ _10252_/S _10251_/X _09181_/X vssd1 vssd1 vccd1 vccd1 _10398_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_102_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11372__A2 _11847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12137_ _12316_/A fanout15/X fanout36/X fanout12/X vssd1 vssd1 vccd1 vccd1 _12138_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07328__A1 _10589_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12068_ _12068_/A _12068_/B vssd1 vssd1 vccd1 vccd1 _12086_/A sky130_fd_sc_hd__xnor2_1
X_11019_ hold282/A _11341_/B _11123_/B _09837_/A vssd1 vssd1 vccd1 vccd1 _11019_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__07328__B2 _08507_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07752__B _07752_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11555__A _12261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11290__A _12261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08230_ fanout75/X _08798_/B2 _07821_/A _08304_/B vssd1 vssd1 vccd1 vccd1 _08231_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_43_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09253__A1 _09423_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09253__B2 _12798_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08056__A2 _08744_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08161_ _08161_/A _08161_/B vssd1 vssd1 vccd1 vccd1 _08253_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__07264__B1 _07282_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07112_ _07113_/A _07113_/B vssd1 vssd1 vccd1 vccd1 _07112_/X sky130_fd_sc_hd__and2_1
XANTENNA__07803__A2 fanout99/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08092_ _08742_/A _08092_/B vssd1 vssd1 vccd1 vccd1 _08096_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_15_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07043_ _11231_/S _07044_/B vssd1 vssd1 vccd1 vccd1 _07043_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_0_43_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout109_A _09716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11363__A2 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08104__A _08731_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08994_ _08994_/A _08994_/B vssd1 vssd1 vccd1 vccd1 _08996_/A sky130_fd_sc_hd__or2_1
XANTENNA__07319__A1 _12804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07945_ _08722_/A _07945_/B vssd1 vssd1 vccd1 vccd1 _07949_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__13156__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07319__B2 _09768_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09615_ _11987_/A _09615_/B _09615_/C vssd1 vssd1 vccd1 vccd1 _09618_/C sky130_fd_sc_hd__and3_1
X_07876_ _07876_/A _07876_/B vssd1 vssd1 vccd1 vccd1 _07943_/B sky130_fd_sc_hd__xor2_1
X_06827_ _11623_/A _11619_/B _06680_/X vssd1 vssd1 vccd1 vccd1 _06827_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_92_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06758_ _06805_/A _06702_/A _12664_/B _06757_/X vssd1 vssd1 vccd1 vccd1 _07080_/A
+ sky130_fd_sc_hd__a31o_4
X_09546_ _09460_/A _09458_/Y _09457_/Y vssd1 vssd1 vccd1 vccd1 _09560_/A sky130_fd_sc_hd__a21o_2
XFILLER_0_66_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09477_ _09478_/B _09478_/A vssd1 vssd1 vccd1 vccd1 _09477_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_108_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06689_ reg1_val[18] _07131_/B vssd1 vssd1 vccd1 vccd1 _06689_/X sky130_fd_sc_hd__and2_1
XFILLER_0_93_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08428_ _08428_/A _08428_/B vssd1 vssd1 vccd1 vccd1 _08451_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13040__A2 _12788_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08359_ _08681_/A _08359_/B vssd1 vssd1 vccd1 vccd1 _08364_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_18_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11370_ _11370_/A _11370_/B vssd1 vssd1 vccd1 vccd1 _11371_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_104_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10321_ _10321_/A fanout7/X vssd1 vssd1 vccd1 vccd1 _10321_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_61_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06741__B _07100_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13040_ hold155/A _12788_/A _13236_/B hold145/X _13109_/A vssd1 vssd1 vccd1 vccd1
+ hold146/A sky130_fd_sc_hd__o221a_1
XANTENNA__09547__A2 fanout16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10252_ _10249_/X _10251_/X _10252_/S vssd1 vssd1 vccd1 vccd1 _10252_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_100_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10183_ _10941_/A fanout48/X _10570_/B fanout94/X vssd1 vssd1 vccd1 vccd1 _10184_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12839__C1 _13214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout282 _06940_/X vssd1 vssd1 vccd1 vccd1 _07200_/A sky130_fd_sc_hd__clkbuf_8
Xfanout271 _06686_/A vssd1 vssd1 vccd1 vccd1 _06695_/A sky130_fd_sc_hd__clkbuf_4
Xfanout260 _07123_/Y vssd1 vssd1 vccd1 vccd1 _09442_/A sky130_fd_sc_hd__buf_12
XANTENNA__11106__A2 _11650_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11375__A _11908_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout293 _13009_/A vssd1 vssd1 vccd1 vccd1 _13013_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_88_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12824_ _12824_/A _12830_/B vssd1 vssd1 vccd1 vccd1 _12824_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_96_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12755_ reg1_val[24] reg1_val[25] _12782_/A vssd1 vssd1 vccd1 vccd1 _12757_/C sky130_fd_sc_hd__o21ai_2
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11706_ _11874_/A _12169_/A _11822_/A vssd1 vssd1 vccd1 vccd1 _11707_/B sky130_fd_sc_hd__a21o_1
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12686_ reg1_val[12] _12686_/B vssd1 vssd1 vccd1 vccd1 _12695_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_37_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11637_ _11636_/B _11724_/B hold293/A vssd1 vssd1 vccd1 vccd1 _11637_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_4_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07246__B1 _12830_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11568_ _11568_/A _11568_/B vssd1 vssd1 vccd1 vccd1 _11569_/B sky130_fd_sc_hd__nand2_1
X_13307_ _13307_/CLK _13307_/D vssd1 vssd1 vccd1 vccd1 hold218/A sky130_fd_sc_hd__dfxtp_1
X_10519_ _11633_/B _10641_/B hold232/A vssd1 vssd1 vccd1 vccd1 _10519_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_97_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12653__B _12654_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06651__B _12664_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11499_ _11499_/A _11499_/B vssd1 vssd1 vccd1 vccd1 _11501_/B sky130_fd_sc_hd__xnor2_1
X_13238_ hold297/X _06892_/B _12783_/Y _06572_/A vssd1 vssd1 vccd1 vccd1 _13238_/X
+ sky130_fd_sc_hd__a22o_1
X_13169_ _12881_/X _13169_/B vssd1 vssd1 vccd1 vccd1 _13170_/B sky130_fd_sc_hd__nand2b_1
X_07730_ _07995_/A _07730_/B vssd1 vssd1 vccd1 vccd1 _07741_/A sky130_fd_sc_hd__or2_1
XANTENNA__09171__B1 _09169_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07661_ _11367_/A _10167_/A1 _10022_/B1 _09745_/B vssd1 vssd1 vccd1 vccd1 _07662_/B
+ sky130_fd_sc_hd__o22a_1
X_06612_ reg1_val[30] _06612_/B vssd1 vssd1 vccd1 vccd1 _06613_/B sky130_fd_sc_hd__nor2_1
X_07592_ _07593_/A _07593_/B vssd1 vssd1 vccd1 vccd1 _09192_/A sky130_fd_sc_hd__nand2b_1
X_09400_ _09400_/A _10818_/A vssd1 vssd1 vccd1 vccd1 _09401_/C sky130_fd_sc_hd__or2_1
XFILLER_0_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12828__B _12830_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09331_ _09329_/X _09330_/X _09669_/S vssd1 vssd1 vccd1 vccd1 _09970_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_87_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09262_ _09262_/A _09262_/B vssd1 vssd1 vccd1 vccd1 _09283_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_63_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12844__A _12844_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09193_ _09209_/B _07492_/B _07501_/B _07502_/B _07502_/A vssd1 vssd1 vccd1 vccd1
+ _09208_/A sky130_fd_sc_hd__a32o_2
XANTENNA__09226__B2 _10706_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09226__A1 _10445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07003__A _12210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08213_ _08213_/A _08213_/B vssd1 vssd1 vccd1 vccd1 _08252_/A sky130_fd_sc_hd__xor2_1
XANTENNA_fanout226_A _12794_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07237__B1 _10941_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09777__A2 _10575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08144_ _08728_/A _08144_/B vssd1 vssd1 vccd1 vccd1 _08169_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_102_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10364__A _10364_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08075_ _08075_/A _08075_/B vssd1 vssd1 vccd1 vccd1 _08872_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_3_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07026_ _07026_/A _07026_/B vssd1 vssd1 vccd1 vccd1 _07026_/X sky130_fd_sc_hd__and2_2
XFILLER_0_101_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10544__B1 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold13 hold13/A vssd1 vssd1 vccd1 vccd1 hold13/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 hold24/A vssd1 vssd1 vccd1 vccd1 hold24/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 hold46/A vssd1 vssd1 vccd1 vccd1 hold46/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13089__A2 fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold35 hold35/A vssd1 vssd1 vccd1 vccd1 hold35/X sky130_fd_sc_hd__dlygate4sd3_1
X_08977_ _08977_/A _08977_/B vssd1 vssd1 vccd1 vccd1 _08978_/B sky130_fd_sc_hd__nand2_1
Xhold57 hold57/A vssd1 vssd1 vccd1 vccd1 hold57/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 hold79/A vssd1 vssd1 vccd1 vccd1 hold79/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09354__C_N _09343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold68 hold68/A vssd1 vssd1 vccd1 vccd1 hold68/X sky130_fd_sc_hd__dlygate4sd3_1
X_07928_ _08752_/A _09613_/A _09614_/A _08798_/B2 vssd1 vssd1 vccd1 vccd1 _07929_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_97_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07859_ _12818_/A fanout87/X fanout82/X _12820_/A vssd1 vssd1 vccd1 vccd1 _07860_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12049__A0 _11973_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10870_ _11100_/A _10870_/B _10870_/C _10870_/D vssd1 vssd1 vccd1 vccd1 _10871_/B
+ sky130_fd_sc_hd__nand4_1
XANTENNA__11923__A _11923_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09529_ _09835_/B _09528_/X hold240/A vssd1 vssd1 vccd1 vccd1 _09529_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout41_A _12834_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06736__B _06963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12540_ _12698_/B _12541_/B vssd1 vssd1 vccd1 vccd1 _12551_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_66_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09217__A1 _12846_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09217__B2 _12848_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12471_ _12644_/B _12471_/B vssd1 vssd1 vccd1 vccd1 _12472_/B sky130_fd_sc_hd__or2_1
XFILLER_0_123_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09768__A2 fanout9/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11422_ _11421_/A _11212_/Y _11421_/B _11420_/A vssd1 vssd1 vccd1 vccd1 _11426_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_123_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08440__A2 _08661_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11353_ _11876_/A _11327_/Y _11328_/X _11352_/X _11326_/X vssd1 vssd1 vccd1 vccd1
+ _11353_/X sky130_fd_sc_hd__a311o_1
X_11284_ _12210_/A _11284_/B vssd1 vssd1 vccd1 vccd1 _11285_/B sky130_fd_sc_hd__xnor2_1
X_10304_ _10303_/B _10304_/B vssd1 vssd1 vccd1 vccd1 _10305_/B sky130_fd_sc_hd__and2b_1
X_13023_ _13214_/A hold119/X vssd1 vssd1 vccd1 vccd1 hold120/A sky130_fd_sc_hd__and2_1
X_10235_ _09652_/B _10232_/X _10233_/X _10234_/X vssd1 vssd1 vccd1 vccd1 _10236_/B
+ sky130_fd_sc_hd__o211a_1
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10166_ _10165_/B _10165_/C _10165_/A vssd1 vssd1 vccd1 vccd1 _10169_/B sky130_fd_sc_hd__a21o_1
XANTENNA__12827__A2 _12830_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10097_ _10097_/A _10368_/A _10496_/A vssd1 vssd1 vccd1 vccd1 _10097_/X sky130_fd_sc_hd__or3_2
XFILLER_0_16_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12807_ _07035_/Y _13087_/B2 hold91/X _13128_/A vssd1 vssd1 vccd1 vccd1 _13257_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_69_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12648__B _12649_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10999_ _11792_/A _10999_/B _10999_/C vssd1 vssd1 vccd1 vccd1 _10999_/X sky130_fd_sc_hd__or3_1
XFILLER_0_9_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10449__A _10449_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12738_ _12730_/Y _12734_/B _12732_/B vssd1 vssd1 vccd1 vccd1 _12739_/B sky130_fd_sc_hd__o21ai_4
XFILLER_0_29_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10066__A2 _07087_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12669_ reg1_val[9] _12669_/B vssd1 vssd1 vccd1 vccd1 _12677_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_115_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07219__B1 _07220_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07758__A _12073_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10184__A _11384_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09880_ _11269_/A _09880_/B vssd1 vssd1 vccd1 vccd1 _09881_/B sky130_fd_sc_hd__xnor2_2
X_08900_ _08900_/A _08900_/B vssd1 vssd1 vccd1 vccd1 _08901_/C sky130_fd_sc_hd__xor2_1
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10526__B1 _10523_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08831_ _08831_/A _08831_/B vssd1 vssd1 vccd1 vccd1 _08834_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_0_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08195__B2 _10537_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08195__A1 _08432_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11727__B _11973_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08762_ _08760_/Y _08762_/B vssd1 vssd1 vccd1 vccd1 _08767_/A sky130_fd_sc_hd__and2b_1
XANTENNA__08498__A2 _08744_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08693_ _08653_/A _08653_/B _08660_/Y _08989_/A _08690_/B vssd1 vssd1 vccd1 vccd1
+ _08693_/X sky130_fd_sc_hd__a221o_1
X_07713_ _07713_/A _07713_/B vssd1 vssd1 vccd1 vccd1 _07716_/A sky130_fd_sc_hd__nor2_1
XANTENNA_fanout176_A _09444_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07644_ _09716_/A _07644_/B vssd1 vssd1 vccd1 vccd1 _07990_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__11743__A _12210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07170__A2 _12842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13243__A2 _06892_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07575_ _07582_/B vssd1 vssd1 vccd1 vccd1 _07575_/Y sky130_fd_sc_hd__inv_2
XANTENNA__09447__B2 _10445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09447__A1 _10706_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09314_ _09092_/X _09111_/X _09351_/B vssd1 vssd1 vccd1 vccd1 _09314_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_36_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09245_ _09245_/A _09245_/B _09237_/Y vssd1 vssd1 vccd1 vccd1 _09247_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_75_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06572__A _06572_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09176_ _09176_/A _09176_/B vssd1 vssd1 vccd1 vccd1 _09179_/A sky130_fd_sc_hd__and2_1
XFILLER_0_71_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10094__A _10096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08127_ _08732_/A1 _08727_/A2 _08727_/B1 _10927_/A1 vssd1 vssd1 vccd1 vccd1 _08128_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_114_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08058_ _08807_/B _08058_/B vssd1 vssd1 vccd1 vccd1 _08808_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07009_ reg1_val[25] _07009_/B vssd1 vssd1 vccd1 vccd1 _07009_/X sky130_fd_sc_hd__xor2_1
XANTENNA__08499__A _08584_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10020_ _09881_/A _09881_/B _09877_/X vssd1 vssd1 vccd1 vccd1 _10021_/B sky130_fd_sc_hd__a21o_1
XANTENNA_fanout89_A _07178_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07933__A1 _11367_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07933__B2 _11472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11971_ _11636_/B _12046_/B hold265/A vssd1 vssd1 vccd1 vccd1 _11971_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__11653__A _11653_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10922_ _10922_/A _10922_/B vssd1 vssd1 vccd1 vccd1 _10923_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_98_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13234__A2 _12790_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10853_ _10854_/A _10854_/B _10854_/C vssd1 vssd1 vccd1 vccd1 _10987_/B sky130_fd_sc_hd__o21ai_2
XANTENNA__11245__A1 _12307_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10784_ _10941_/A fanout59/X _10941_/B fanout94/X vssd1 vssd1 vccd1 vccd1 _10785_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_27_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12523_ _12523_/A _12523_/B _12523_/C vssd1 vssd1 vccd1 vccd1 _12524_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_94_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12484__A _12654_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08661__A2 _08661_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12454_ _12460_/B _12454_/B vssd1 vssd1 vccd1 vccd1 new_PC[1] sky130_fd_sc_hd__and2_4
XFILLER_0_62_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12385_ _12382_/Y _12384_/X _12290_/A vssd1 vssd1 vccd1 vccd1 _12385_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_34_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11405_ _11405_/A _11405_/B vssd1 vssd1 vccd1 vccd1 _11408_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_120_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11336_ _11334_/Y _11336_/B vssd1 vssd1 vccd1 vccd1 _11337_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_104_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13006_ hold225/A _13016_/A2 _13006_/B1 hold192/X vssd1 vssd1 vccd1 vccd1 hold193/A
+ sky130_fd_sc_hd__a22o_1
X_11267_ _11267_/A _11267_/B vssd1 vssd1 vccd1 vccd1 _11275_/A sky130_fd_sc_hd__nand2_1
X_10218_ _10218_/A _10218_/B vssd1 vssd1 vccd1 vccd1 _10220_/B sky130_fd_sc_hd__and2_1
X_11198_ _11198_/A _11198_/B vssd1 vssd1 vccd1 vccd1 _11201_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__07924__A1 _12820_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07924__B2 _08741_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10149_ _10149_/A _10149_/B vssd1 vssd1 vccd1 vccd1 _10178_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__11563__A _11908_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07152__A2 _07343_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11484__B2 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11484__A1 fanout27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07360_ _07360_/A _07360_/B vssd1 vssd1 vccd1 vccd1 _07362_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_128_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08101__B2 _08732_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08101__A1 _08741_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_252 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12394__A _12394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07291_ _07647_/A _07647_/B vssd1 vssd1 vccd1 vccd1 _07292_/B sky130_fd_sc_hd__and2b_1
X_09030_ _08341_/Y _08715_/B _08342_/X vssd1 vssd1 vccd1 vccd1 _09030_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_45_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold302 hold302/A vssd1 vssd1 vccd1 vccd1 hold302/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10118__S _11118_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09932_ _09932_/A _09932_/B vssd1 vssd1 vccd1 vccd1 _09945_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_40_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09863_ _09863_/A _09863_/B vssd1 vssd1 vccd1 vccd1 _09864_/B sky130_fd_sc_hd__nor2_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09794_ _09560_/A _09560_/B _09559_/A vssd1 vssd1 vccd1 vccd1 _09799_/A sky130_fd_sc_hd__a21o_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08814_ _08813_/B _08813_/C _08813_/A vssd1 vssd1 vccd1 vccd1 _08815_/C sky130_fd_sc_hd__a21oi_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08745_ _08745_/A _08745_/B vssd1 vssd1 vccd1 vccd1 _08747_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07951__A _08724_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11473__A _11557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08676_ _08677_/B _08677_/C _08678_/A vssd1 vssd1 vccd1 vccd1 _08685_/A sky130_fd_sc_hd__a21oi_1
XTAP_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07627_ _07627_/A _08918_/A vssd1 vssd1 vccd1 vccd1 _07669_/A sky130_fd_sc_hd__or2_1
X_07558_ _07558_/A _07558_/B vssd1 vssd1 vccd1 vccd1 _07559_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_48_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09089__S _09108_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07489_ _08724_/A _07489_/B vssd1 vssd1 vccd1 vccd1 _07491_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_118_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09228_ _12826_/A fanout69/X _08216_/B _12828_/A vssd1 vssd1 vccd1 vccd1 _09229_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_8_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09159_ _09168_/A _09159_/B vssd1 vssd1 vccd1 vccd1 _09159_/X sky130_fd_sc_hd__or2_1
XFILLER_0_90_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09817__S _12388_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12170_ _12170_/A _12170_/B _12287_/A vssd1 vssd1 vccd1 vccd1 _12172_/B sky130_fd_sc_hd__and3_1
XFILLER_0_32_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11121_ _12394_/A _11121_/B vssd1 vssd1 vccd1 vccd1 _11121_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_7_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13152__B2 _13246_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11367__B _12214_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11052_ _10575_/A _11989_/A _10570_/B _10574_/A vssd1 vssd1 vccd1 vccd1 _11053_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__06709__A2 _06587_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10003_ _09907_/Y _09911_/A _07035_/Y _10959_/A vssd1 vssd1 vccd1 vccd1 _10211_/A
+ sky130_fd_sc_hd__o211a_1
XANTENNA__07382__A2 _10413_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11383__A _11758_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11954_ _11953_/A _11953_/B _11953_/Y _11876_/A vssd1 vssd1 vccd1 vccd1 _11954_/X
+ sky130_fd_sc_hd__o211a_1
X_11885_ _11885_/A _11885_/B vssd1 vssd1 vccd1 vccd1 _11886_/B sky130_fd_sc_hd__xnor2_1
X_10905_ _10874_/Y _10875_/X _10904_/X _10873_/Y vssd1 vssd1 vccd1 vccd1 _10905_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_58_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10836_ _10976_/A _10836_/B vssd1 vssd1 vccd1 vccd1 _10838_/B sky130_fd_sc_hd__and2_1
XFILLER_0_94_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10767_ _09527_/B _09354_/B _10767_/S vssd1 vssd1 vccd1 vccd1 _10767_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_109_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12506_ _12669_/B _12506_/B vssd1 vssd1 vccd1 vccd1 _12507_/B sky130_fd_sc_hd__or2_1
XFILLER_0_42_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10698_ _10580_/B _10583_/B _10578_/X vssd1 vssd1 vccd1 vccd1 _10700_/B sky130_fd_sc_hd__a21o_1
X_12437_ reg1_val[31] _07064_/B _11973_/B _12436_/X _12404_/A vssd1 vssd1 vccd1 vccd1
+ _12437_/X sky130_fd_sc_hd__a311o_1
XANTENNA__07101__A _11385_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12368_ _12368_/A vssd1 vssd1 vccd1 vccd1 _12418_/S sky130_fd_sc_hd__inv_2
X_12299_ _12429_/B _12299_/B vssd1 vssd1 vccd1 vccd1 _12299_/Y sky130_fd_sc_hd__nor2_1
X_11319_ _11319_/A _11514_/A vssd1 vssd1 vccd1 vccd1 _11319_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__11558__A _11558_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10462__A _11163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06860_ _12389_/A _06859_/Y _06837_/Y vssd1 vssd1 vccd1 vccd1 _12423_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__12351__C1 _06924_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11154__B1 fanout4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06791_ _06789_/Y _06791_/B vssd1 vssd1 vccd1 vccd1 _09686_/B sky130_fd_sc_hd__nand2b_2
XFILLER_0_89_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11457__A1 _09156_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08530_ _08530_/A _08530_/B vssd1 vssd1 vccd1 vccd1 _08560_/B sky130_fd_sc_hd__xnor2_1
X_08461_ _09441_/A _08461_/B vssd1 vssd1 vccd1 vccd1 _08467_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_54_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07412_ _07413_/A _07413_/B vssd1 vssd1 vccd1 vccd1 _07460_/B sky130_fd_sc_hd__or2_1
XFILLER_0_9_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08392_ _08393_/B _08393_/C _08645_/A vssd1 vssd1 vccd1 vccd1 _08394_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_58_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07343_ _06838_/B _07343_/B vssd1 vssd1 vccd1 vccd1 _07343_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_70_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08086__B1 _08617_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout139_A _12810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07274_ _07485_/A _07274_/B vssd1 vssd1 vccd1 vccd1 _07278_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_45_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09013_ _09013_/A _09013_/B vssd1 vssd1 vccd1 vccd1 _09015_/B sky130_fd_sc_hd__nor2_1
XANTENNA__07011__A _09716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12852__A _12852_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold110 hold110/A vssd1 vssd1 vccd1 vccd1 hold110/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout306_A _06574_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold132 hold132/A vssd1 vssd1 vccd1 vccd1 hold132/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold121 hold121/A vssd1 vssd1 vccd1 vccd1 hold121/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold143 hold143/A vssd1 vssd1 vccd1 vccd1 hold143/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold176 hold176/A vssd1 vssd1 vccd1 vccd1 hold176/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold165 hold165/A vssd1 vssd1 vccd1 vccd1 hold165/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold154 hold154/A vssd1 vssd1 vccd1 vccd1 hold154/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11468__A _11908_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold198 hold198/A vssd1 vssd1 vccd1 vccd1 hold198/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold187 hold187/A vssd1 vssd1 vccd1 vccd1 hold187/X sky130_fd_sc_hd__dlygate4sd3_1
X_09915_ _12808_/A _10797_/B vssd1 vssd1 vccd1 vccd1 _09917_/C sky130_fd_sc_hd__nor2_1
X_09846_ _09828_/Y _09830_/Y _09832_/Y _09833_/X _09845_/X vssd1 vssd1 vccd1 vccd1
+ _09846_/X sky130_fd_sc_hd__o221a_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12299__A _12429_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06989_ _12822_/A fanout74/X _10948_/B2 _12824_/A vssd1 vssd1 vccd1 vccd1 _06990_/B
+ sky130_fd_sc_hd__o22a_1
X_09777_ _11065_/A _10575_/A _10963_/A _09613_/A vssd1 vssd1 vccd1 vccd1 _09778_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11448__A1 _09152_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08728_ _08728_/A _08728_/B vssd1 vssd1 vccd1 vccd1 _08736_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_96_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08659_ _08689_/A _08689_/B _08689_/C vssd1 vssd1 vccd1 vccd1 _08690_/A sky130_fd_sc_hd__o21a_1
XANTENNA__11999__A2 _12316_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10671__A2 _12150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11670_ _11670_/A _11670_/B vssd1 vssd1 vccd1 vccd1 _11671_/B sky130_fd_sc_hd__and2_1
XANTENNA__06698__A_N _07130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06744__B _06799_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10621_ _09489_/B _10097_/X _10617_/X _10618_/Y _10620_/Y vssd1 vssd1 vccd1 vccd1
+ _10622_/B sky130_fd_sc_hd__o311ai_4
XANTENNA__11650__B _11650_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09401__A _11987_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13340_ _13340_/CLK _13340_/D vssd1 vssd1 vccd1 vccd1 hold67/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11142__S _11142_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10552_ _10963_/A fanout16/X _07282_/B _11065_/A vssd1 vssd1 vccd1 vccd1 _10553_/B
+ sky130_fd_sc_hd__o22a_1
X_13271_ _13376_/CLK hold16/X vssd1 vssd1 vccd1 vccd1 hold15/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12222_ _12154_/A _12157_/A _12277_/B _12221_/X vssd1 vssd1 vccd1 vccd1 _12222_/Y
+ sky130_fd_sc_hd__a211oi_1
X_10483_ _10483_/A _10483_/B vssd1 vssd1 vccd1 vccd1 _10484_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_20_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12153_ _12153_/A _12153_/B vssd1 vssd1 vccd1 vccd1 _12154_/B sky130_fd_sc_hd__nand2_1
XANTENNA__10282__A _11261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11104_ _11318_/A _11104_/B vssd1 vssd1 vccd1 vccd1 _11650_/B sky130_fd_sc_hd__xor2_4
X_12084_ _12084_/A _12084_/B vssd1 vssd1 vccd1 vccd1 _12086_/B sky130_fd_sc_hd__xnor2_1
X_11035_ fanout29/X _11558_/A _10575_/B fanout27/X vssd1 vssd1 vccd1 vccd1 _11036_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08552__A1 _08730_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08552__B2 _12808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06919__B _06921_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12986_ _13295_/Q _13004_/A2 _13006_/B1 hold212/X vssd1 vssd1 vccd1 vccd1 hold213/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_86_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11937_ _11854_/A _11852_/X _11851_/Y vssd1 vssd1 vccd1 vccd1 _11939_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_24_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06935__A _12455_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11868_ _11868_/A _12024_/B vssd1 vssd1 vccd1 vccd1 _11868_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__10662__A2 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11799_ reg1_val[21] curr_PC[21] vssd1 vssd1 vccd1 vccd1 _11800_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_55_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10819_ _10820_/B _10820_/A vssd1 vssd1 vccd1 vccd1 _10819_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_27_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06654__B _07194_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10414__A2 _12316_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07766__A _08724_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07961_ _08031_/A vssd1 vssd1 vccd1 vccd1 _08076_/A sky130_fd_sc_hd__inv_2
X_06912_ instruction[15] _06884_/Y _06911_/X _06634_/B vssd1 vssd1 vccd1 vccd1 reg1_idx[4]
+ sky130_fd_sc_hd__o211a_4
X_09700_ curr_PC[3] _09701_/B vssd1 vssd1 vccd1 vccd1 _09700_/X sky130_fd_sc_hd__or2_1
XANTENNA__07346__A2 _12852_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07892_ _08724_/A _07892_/B vssd1 vssd1 vccd1 vccd1 _07915_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__10920__A _11180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06843_ reg1_val[24] _07140_/C vssd1 vssd1 vccd1 vccd1 _06843_/X sky130_fd_sc_hd__and2_1
X_09631_ _09467_/A _09467_/B _09466_/A vssd1 vssd1 vccd1 vccd1 _09641_/A sky130_fd_sc_hd__a21o_2
X_06774_ reg1_val[5] _06774_/B vssd1 vssd1 vccd1 vccd1 _06774_/X sky130_fd_sc_hd__and2_1
XANTENNA__06829__B _07135_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09562_ _09439_/A _09438_/Y _09434_/Y vssd1 vssd1 vccd1 vccd1 _09564_/A sky130_fd_sc_hd__a21o_1
XANTENNA__07006__A _09666_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08513_ _08494_/A _08494_/B _08512_/Y vssd1 vssd1 vccd1 vccd1 _09010_/A sky130_fd_sc_hd__a21bo_1
XANTENNA_fanout256_A _08436_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09493_ _08983_/A _08985_/A _09653_/A _09163_/X _09492_/Y vssd1 vssd1 vccd1 vccd1
+ _09493_/X sky130_fd_sc_hd__a311o_1
XANTENNA__11751__A _11751_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08444_ _08444_/A _08444_/B vssd1 vssd1 vccd1 vccd1 _08446_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_92_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08375_ _08372_/A _08372_/B _08374_/Y vssd1 vssd1 vccd1 vccd1 _08385_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__11470__B _11470_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07326_ _07398_/B _07398_/A vssd1 vssd1 vccd1 vccd1 _07326_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_60_101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07257_ _12317_/A vssd1 vssd1 vccd1 vccd1 _12138_/A sky130_fd_sc_hd__inv_4
XFILLER_0_5_250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07188_ _09441_/A _07188_/B vssd1 vssd1 vccd1 vccd1 _10024_/A sky130_fd_sc_hd__nand2_1
XANTENNA__11905__A2 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06793__B1 _06792_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09829_ _12394_/A _09172_/B _09152_/Y vssd1 vssd1 vccd1 vccd1 _09830_/A sky130_fd_sc_hd__a21o_1
X_12840_ _12840_/A _12848_/B vssd1 vssd1 vccd1 vccd1 _12840_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_96_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12771_ reg1_val[29] _12782_/A vssd1 vssd1 vccd1 vccd1 _12772_/B sky130_fd_sc_hd__or2_1
X_11722_ hold210/A _11450_/B _11805_/B _11968_/B1 vssd1 vssd1 vccd1 vccd1 _11723_/B
+ sky130_fd_sc_hd__a31o_1
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11653_ _11653_/A fanout8/X vssd1 vssd1 vccd1 vccd1 _11654_/B sky130_fd_sc_hd__nor2_1
Xfanout60 _07145_/X vssd1 vssd1 vccd1 vccd1 _12848_/A sky130_fd_sc_hd__buf_4
Xfanout82 _08507_/B vssd1 vssd1 vccd1 vccd1 fanout82/X sky130_fd_sc_hd__buf_6
Xfanout71 _07052_/Y vssd1 vssd1 vccd1 vccd1 _07819_/B sky130_fd_sc_hd__buf_8
X_10604_ _10604_/A _10604_/B vssd1 vssd1 vccd1 vccd1 _10606_/A sky130_fd_sc_hd__or2_2
X_13323_ _13343_/CLK hold147/X vssd1 vssd1 vccd1 vccd1 hold145/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout93 _07833_/A vssd1 vssd1 vccd1 vccd1 _09746_/A sky130_fd_sc_hd__buf_4
X_11584_ _11489_/A _11489_/B _11479_/A vssd1 vssd1 vccd1 vccd1 _11596_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__12492__A _12659_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07273__A1 fanout69/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07273__B2 _10963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10535_ _10485_/A _10485_/B _10486_/X vssd1 vssd1 vccd1 vccd1 _10612_/A sky130_fd_sc_hd__a21o_2
X_13254_ _13380_/CLK _13254_/D vssd1 vssd1 vccd1 vccd1 hold88/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12149__A2 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10466_ _10941_/A _10571_/B fanout51/X fanout94/X vssd1 vssd1 vccd1 vccd1 _10467_/B
+ sky130_fd_sc_hd__o22a_1
X_13185_ hold293/A _13184_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13185_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_122_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12205_ _12170_/B _12287_/A _12170_/A vssd1 vssd1 vccd1 vccd1 _12205_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_60_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10397_ _06756_/B _09354_/B _10392_/Y _06754_/Y _10396_/X vssd1 vssd1 vccd1 vccd1
+ _10397_/X sky130_fd_sc_hd__o221a_1
X_12136_ _12066_/B _12068_/B _12066_/A vssd1 vssd1 vccd1 vccd1 _12148_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_19_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12067_ _12067_/A _12214_/B vssd1 vssd1 vccd1 vccd1 _12068_/B sky130_fd_sc_hd__nor2_1
X_11018_ _11341_/B _11123_/B hold282/A vssd1 vssd1 vccd1 vccd1 _11018_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__07328__A2 _12832_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12969_ _13009_/A hold235/X vssd1 vssd1 vccd1 vccd1 _13287_/D sky130_fd_sc_hd__and2_1
XFILLER_0_75_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09976__A _11118_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08160_ _08161_/A _08161_/B vssd1 vssd1 vccd1 vccd1 _08160_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_28_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12793__C1 _13128_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09253__A2 fanout9/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07111_ _11987_/A _07111_/B vssd1 vssd1 vccd1 vccd1 _07113_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_28_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07264__B2 _08671_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07264__A1 _12794_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08091_ _12818_/A _08741_/A2 _08617_/B _12820_/A vssd1 vssd1 vccd1 vccd1 _08092_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07042_ _10248_/S _09666_/S _09351_/B _07064_/B _12341_/A vssd1 vssd1 vccd1 vccd1
+ _07044_/B sky130_fd_sc_hd__o311a_2
XANTENNA__07496__A _09897_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09187__S _11343_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11899__A1 _11624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08993_ _08993_/A _08993_/B vssd1 vssd1 vccd1 vccd1 _08994_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_11_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07944_ _10537_/A1 _08739_/A1 _08436_/A _08432_/B vssd1 vssd1 vccd1 vccd1 _07945_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09216__A _09431_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07319__A2 fanout23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09713__B1 _07282_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07875_ _07876_/A _07876_/B vssd1 vssd1 vccd1 vccd1 _07875_/X sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_4_2_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06826_ _06693_/X _11524_/B _06689_/X vssd1 vssd1 vccd1 vccd1 _11619_/B sky130_fd_sc_hd__a21o_1
XANTENNA__11520__B1 _12290_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09614_ _09614_/A _10963_/A vssd1 vssd1 vccd1 vccd1 _09615_/C sky130_fd_sc_hd__or2_1
X_09545_ _09476_/A _09476_/B _09477_/Y vssd1 vssd1 vccd1 vccd1 _09644_/A sky130_fd_sc_hd__o21ai_4
X_06757_ reg2_val[7] _06799_/B vssd1 vssd1 vccd1 vccd1 _06757_/X sky130_fd_sc_hd__and2_1
X_06688_ _06686_/Y _06703_/B1 _06720_/B reg2_val[18] vssd1 vssd1 vccd1 vccd1 _06691_/B
+ sky130_fd_sc_hd__a2bb2o_2
X_09476_ _09476_/A _09476_/B vssd1 vssd1 vccd1 vccd1 _09478_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__11481__A _12317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08427_ _09023_/A vssd1 vssd1 vccd1 vccd1 _08427_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_19_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08358_ _12818_/A _08436_/B _12820_/A _07149_/A vssd1 vssd1 vccd1 vccd1 _08359_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_46_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07309_ _07309_/A _07309_/B vssd1 vssd1 vccd1 vccd1 _07602_/B sky130_fd_sc_hd__xnor2_4
X_08289_ _08345_/A _08345_/B vssd1 vssd1 vccd1 vccd1 _08346_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_34_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13201__A _13214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10320_ _10320_/A fanout7/X vssd1 vssd1 vccd1 vccd1 _10320_/X sky130_fd_sc_hd__or2_1
XFILLER_0_21_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10251_ _09179_/A _10250_/X _11118_/A vssd1 vssd1 vccd1 vccd1 _10251_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10011__B1 _08507_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10182_ _10448_/A _10182_/B vssd1 vssd1 vccd1 vccd1 _10186_/A sky130_fd_sc_hd__xnor2_1
Xfanout250 _12247_/C1 vssd1 vssd1 vccd1 vccd1 _09837_/A sky130_fd_sc_hd__buf_4
XFILLER_0_100_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout283 _12611_/A vssd1 vssd1 vccd1 vccd1 _12623_/A sky130_fd_sc_hd__buf_8
Xfanout272 _06635_/A vssd1 vssd1 vccd1 vccd1 _06686_/A sky130_fd_sc_hd__clkbuf_4
Xfanout294 _06578_/Y vssd1 vssd1 vccd1 vccd1 _13009_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_88_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12823_ hold23/X _12830_/B _12822_/Y _13245_/A vssd1 vssd1 vccd1 vccd1 hold24/A sky130_fd_sc_hd__o211a_1
XANTENNA__11814__A1 _09111_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12754_ _12754_/A _12754_/B vssd1 vssd1 vccd1 vccd1 _12766_/B sky130_fd_sc_hd__or2_1
XFILLER_0_96_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11705_ _11874_/A _12169_/A _11822_/A vssd1 vssd1 vccd1 vccd1 _11705_/X sky130_fd_sc_hd__and3_1
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12685_ reg1_val[12] _12686_/B vssd1 vssd1 vccd1 vccd1 _12687_/A sky130_fd_sc_hd__or2_1
X_11636_ hold293/A _11636_/B _11724_/B vssd1 vssd1 vccd1 vccd1 _11636_/X sky130_fd_sc_hd__and3_1
XFILLER_0_71_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07246__A1 _12828_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07246__B2 _08507_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11567_ _11568_/A _11568_/B vssd1 vssd1 vccd1 vccd1 _11569_/A sky130_fd_sc_hd__or2_1
XFILLER_0_21_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13306_ _13307_/CLK hold194/X vssd1 vssd1 vccd1 vccd1 hold192/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10518_ hold220/A _10518_/B vssd1 vssd1 vccd1 vccd1 _10641_/B sky130_fd_sc_hd__or2_1
XANTENNA__11330__S _12174_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13237_ hold63/X _13246_/B2 _13109_/A _13236_/Y vssd1 vssd1 vccd1 vccd1 hold66/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_52_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11498_ _11499_/B _11499_/A vssd1 vssd1 vccd1 vccd1 _11599_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_122_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10449_ _10449_/A _10449_/B _10449_/C vssd1 vssd1 vccd1 vccd1 _10449_/X sky130_fd_sc_hd__and3_1
XFILLER_0_20_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13168_ _13245_/A _13168_/B vssd1 vssd1 vccd1 vccd1 _13363_/D sky130_fd_sc_hd__and2_1
XFILLER_0_0_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_384 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12119_ hold254/A _12119_/B vssd1 vssd1 vccd1 vccd1 _12187_/B sky130_fd_sc_hd__or2_1
X_13099_ hold240/X _06892_/B _13098_/X _06572_/A vssd1 vssd1 vccd1 vccd1 hold241/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11566__A _11758_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09171__A1 hold260/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07660_ _10165_/A _07660_/B vssd1 vssd1 vccd1 vccd1 _07729_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_46_98 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06611_ reg1_val[30] _06612_/B vssd1 vssd1 vccd1 vccd1 _12402_/S sky130_fd_sc_hd__and2_1
X_07591_ _07394_/A _07394_/B _07392_/X vssd1 vssd1 vccd1 vccd1 _07593_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_1_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09330_ _09124_/X _09126_/X _09330_/S vssd1 vssd1 vccd1 vccd1 _09330_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_75_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09261_ _09260_/B _09260_/C _09260_/A vssd1 vssd1 vccd1 vccd1 _09262_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_117_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08212_ _08213_/A _08213_/B vssd1 vssd1 vccd1 vccd1 _08212_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__06759__A_N _07080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09192_ _09192_/A _09192_/B vssd1 vssd1 vccd1 vccd1 _09299_/A sky130_fd_sc_hd__nand2_4
XANTENNA__09226__A2 _12834_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07237__B2 _07149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07237__A1 _12848_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout121_A _08432_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08143_ _08741_/B2 _08727_/A2 _08727_/B1 _08732_/A1 vssd1 vssd1 vccd1 vccd1 _08144_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__13021__A _13214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout219_A _13213_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06842__B _07169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08074_ _08073_/A _08073_/B _08073_/C vssd1 vssd1 vccd1 vccd1 _08075_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_16_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07025_ _07074_/B _06964_/A _07023_/X _06774_/B vssd1 vssd1 vccd1 vccd1 _07026_/B
+ sky130_fd_sc_hd__a211o_1
XANTENNA__10364__B _10364_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08115__A _08740_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10544__A1 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold14 hold14/A vssd1 vssd1 vccd1 vccd1 hold14/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10544__B2 _10948_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold25 hold25/A vssd1 vssd1 vccd1 vccd1 hold25/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 hold47/A vssd1 vssd1 vccd1 vccd1 hold47/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 hold36/A vssd1 vssd1 vccd1 vccd1 hold36/X sky130_fd_sc_hd__dlygate4sd3_1
X_08976_ _09485_/B _09649_/B _08975_/Y _09487_/C _09487_/B vssd1 vssd1 vccd1 vccd1
+ _08977_/B sky130_fd_sc_hd__o32a_1
Xhold58 hold58/A vssd1 vssd1 vccd1 vccd1 hold58/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold69 hold69/A vssd1 vssd1 vccd1 vccd1 hold69/X sky130_fd_sc_hd__dlygate4sd3_1
X_07927_ _08029_/A _07926_/Y _07922_/Y vssd1 vssd1 vccd1 vccd1 _07940_/A sky130_fd_sc_hd__a21oi_2
X_07858_ _08742_/A _07858_/B vssd1 vssd1 vccd1 vccd1 _07862_/A sky130_fd_sc_hd__xnor2_1
X_06809_ _09350_/A _09350_/B _06802_/X vssd1 vssd1 vccd1 vccd1 _06809_/X sky130_fd_sc_hd__a21o_1
XANTENNA__11923__B _12412_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07789_ _07790_/A _07790_/B vssd1 vssd1 vccd1 vccd1 _07789_/X sky130_fd_sc_hd__or2_1
X_09528_ hold244/A hold260/A vssd1 vssd1 vccd1 vccd1 _09528_/X sky130_fd_sc_hd__or2_1
XFILLER_0_78_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout34_A _12264_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09459_ _09459_/A _09459_/B vssd1 vssd1 vccd1 vccd1 _09460_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_108_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09217__A2 _09567_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12470_ _12644_/B _12471_/B vssd1 vssd1 vccd1 vccd1 _12481_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_47_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11421_ _11421_/A _11421_/B vssd1 vssd1 vccd1 vccd1 _11608_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_104_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11352_ _09156_/Y _11331_/X _11332_/Y _11351_/X vssd1 vssd1 vccd1 vccd1 _11352_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_22_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10303_ _10304_/B _10303_/B vssd1 vssd1 vccd1 vccd1 _10480_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_104_386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11283_ fanout27/X _11847_/A _11766_/A fanout29/X vssd1 vssd1 vccd1 vccd1 _11284_/B
+ sky130_fd_sc_hd__o22a_1
X_13022_ hold215/A _13213_/B2 _13213_/A2 hold118/X vssd1 vssd1 vccd1 vccd1 hold119/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__06739__B1 _06738_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10234_ _09645_/X _09806_/X _09807_/X _10496_/A _10617_/A vssd1 vssd1 vccd1 vccd1
+ _10234_/X sky130_fd_sc_hd__a2111o_1
XANTENNA__07864__A _08745_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10165_ _10165_/A _10165_/B _10165_/C vssd1 vssd1 vccd1 vccd1 _10169_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_83_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10096_ _10096_/A _10096_/B vssd1 vssd1 vccd1 vccd1 _10617_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_89_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12806_ hold90/X _12818_/B vssd1 vssd1 vccd1 vccd1 hold91/A sky130_fd_sc_hd__or2_1
XFILLER_0_97_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10998_ _10909_/X _10996_/Y _10997_/Y vssd1 vssd1 vccd1 vccd1 _10998_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_8_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12737_ _12737_/A _12737_/B vssd1 vssd1 vccd1 vccd1 _12746_/C sky130_fd_sc_hd__nand2_2
XFILLER_0_84_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12668_ reg1_val[9] _12669_/B vssd1 vssd1 vccd1 vccd1 _12675_/B sky130_fd_sc_hd__or2_1
X_11619_ _12174_/S _11619_/B vssd1 vssd1 vccd1 vccd1 _11623_/B sky130_fd_sc_hd__or2_1
XANTENNA__07219__A1 _07220_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12664__B _12664_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12599_ reg1_val[23] curr_PC[23] _12622_/S vssd1 vssd1 vccd1 vccd1 _12600_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_53_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07774__A _11758_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09916__B1 _10959_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10526__B2 _10524_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08830_ _08831_/A _08831_/B vssd1 vssd1 vccd1 vccd1 _08864_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_0_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08195__A2 _07896_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06745__A3 _12673_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08761_ _08761_/A _08761_/B vssd1 vssd1 vccd1 vccd1 _08762_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_79_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08692_ _08629_/X _08638_/Y _08622_/B _08626_/Y vssd1 vssd1 vccd1 vccd1 _08695_/B
+ sky130_fd_sc_hd__o211a_1
X_07712_ _07712_/A _07712_/B vssd1 vssd1 vccd1 vccd1 _07713_/B sky130_fd_sc_hd__nor2_1
XANTENNA__10829__A2 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07643_ _12798_/A fanout24/X _07819_/B _09423_/B2 vssd1 vssd1 vccd1 vccd1 _07644_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11239__C1 _09169_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout169_A _09568_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09313_ _09311_/X _09312_/X _09666_/S vssd1 vssd1 vccd1 vccd1 _09313_/X sky130_fd_sc_hd__mux2_1
X_07574_ _07574_/A _07574_/B vssd1 vssd1 vccd1 vccd1 _07582_/B sky130_fd_sc_hd__or2_2
XANTENNA__09447__A2 fanout48/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09244_ _09242_/B _09242_/C _09593_/A vssd1 vssd1 vccd1 vccd1 _09244_/X sky130_fd_sc_hd__a21o_1
X_09175_ _09974_/A _09181_/B vssd1 vssd1 vccd1 vccd1 _09176_/B sky130_fd_sc_hd__or2_2
XFILLER_0_90_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12203__A1 _12455_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08126_ _08130_/A _08130_/B vssd1 vssd1 vccd1 vccd1 _08126_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_120_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06969__B1 _11343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10094__B _10096_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08057_ _08745_/A _08057_/B vssd1 vssd1 vccd1 vccd1 _08807_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_113_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07008_ reg1_val[24] _07254_/B _07254_/C _07364_/B1 vssd1 vssd1 vccd1 vccd1 _07009_/B
+ sky130_fd_sc_hd__o31a_1
XANTENNA__07933__A2 _08732_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08959_ _08959_/A _08959_/B vssd1 vssd1 vccd1 vccd1 _08960_/B sky130_fd_sc_hd__xnor2_2
X_11970_ hold246/A _11970_/B vssd1 vssd1 vccd1 vccd1 _12046_/B sky130_fd_sc_hd__or2_1
XFILLER_0_98_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07146__B1 _09236_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11653__B fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10921_ _10922_/A _10922_/B vssd1 vssd1 vccd1 vccd1 _10923_/A sky130_fd_sc_hd__and2_1
XANTENNA__06747__B _07095_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10852_ _10852_/A _10852_/B vssd1 vssd1 vccd1 vccd1 _10854_/C sky130_fd_sc_hd__xor2_1
XANTENNA__08646__B1 _08673_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10783_ _11792_/A _10783_/B vssd1 vssd1 vccd1 vccd1 _10783_/X sky130_fd_sc_hd__or2_1
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12522_ _12523_/A _12523_/B _12523_/C vssd1 vssd1 vccd1 vccd1 _12530_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_93_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12453_ _12453_/A _12453_/B vssd1 vssd1 vccd1 vccd1 _12454_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_35_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12384_ _12287_/A _12287_/B _12383_/X _12170_/A vssd1 vssd1 vccd1 vccd1 _12384_/X
+ sky130_fd_sc_hd__o31a_1
X_11404_ _11404_/A _11404_/B vssd1 vssd1 vccd1 vccd1 _11405_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_22_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11335_ reg1_val[16] curr_PC[16] vssd1 vssd1 vccd1 vccd1 _11336_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_105_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11266_ _11266_/A _11266_/B vssd1 vssd1 vccd1 vccd1 _11267_/B sky130_fd_sc_hd__or2_1
X_13005_ _13009_/A hold226/X vssd1 vssd1 vccd1 vccd1 hold227/A sky130_fd_sc_hd__and2_1
XFILLER_0_120_676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10217_ _10047_/A _10047_/B _10045_/Y vssd1 vssd1 vccd1 vccd1 _10220_/A sky130_fd_sc_hd__o21ai_4
XFILLER_0_94_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11197_ _11197_/A _11197_/B vssd1 vssd1 vccd1 vccd1 _11198_/B sky130_fd_sc_hd__and2_1
XANTENNA__06727__A3 _12692_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07924__A2 _08744_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10148_ _10148_/A _12316_/B vssd1 vssd1 vccd1 vccd1 _10149_/B sky130_fd_sc_hd__or2_1
X_10079_ _10079_/A _10079_/B vssd1 vssd1 vccd1 vccd1 _10092_/A sky130_fd_sc_hd__xor2_4
XANTENNA__11844__A _12261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06938__A _12423_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12659__B _12659_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06657__B _12659_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11484__A2 _11989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_354 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07290_ _07290_/A _07290_/B vssd1 vssd1 vccd1 vccd1 _07647_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_45_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08101__A2 _08732_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12197__B1 _12254_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold303 hold303/A vssd1 vssd1 vccd1 vccd1 hold303/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09931_ _09931_/A _09931_/B vssd1 vssd1 vccd1 vccd1 _09932_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_13_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09862_ _09863_/A _09863_/B vssd1 vssd1 vccd1 vccd1 _09864_/A sky130_fd_sc_hd__and2_1
XFILLER_0_0_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09793_ _09637_/A _09637_/B _09635_/X vssd1 vssd1 vccd1 vccd1 _09800_/A sky130_fd_sc_hd__a21bo_1
X_08813_ _08813_/A _08813_/B _08813_/C vssd1 vssd1 vccd1 vccd1 _08815_/B sky130_fd_sc_hd__and3_1
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout286_A _06587_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08744_ fanout99/X _08744_/A2 _08564_/B _12818_/A vssd1 vssd1 vccd1 vccd1 _08745_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12121__B1 _12247_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08675_ _08728_/A _08678_/B vssd1 vssd1 vccd1 vccd1 _08677_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_67_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07626_ _08917_/B _07626_/B vssd1 vssd1 vccd1 vccd1 _08918_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_88_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07557_ _07558_/A _07558_/B vssd1 vssd1 vccd1 vccd1 _07557_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07488_ _12828_/A fanout74/X _10948_/B2 _12830_/A vssd1 vssd1 vccd1 vccd1 _07489_/B
+ sky130_fd_sc_hd__o22a_1
X_09227_ _10707_/A _09227_/B vssd1 vssd1 vccd1 vccd1 _09231_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_16_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09158_ _09168_/A _09159_/B vssd1 vssd1 vccd1 vccd1 _09158_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_90_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09894__A _10165_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09089_ reg1_val[2] reg1_val[29] _09108_/S vssd1 vssd1 vccd1 vccd1 _09089_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_32_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08109_ _08110_/A _08110_/B vssd1 vssd1 vccd1 vccd1 _08111_/A sky130_fd_sc_hd__nand2_1
X_11120_ _10119_/S _09368_/Y _11119_/X vssd1 vssd1 vccd1 vccd1 _11121_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_102_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08303__A _08722_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13152__A2 _06890_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06658__A2_N _06771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11051_ _11269_/A _11051_/B vssd1 vssd1 vccd1 vccd1 _11055_/A sky130_fd_sc_hd__xnor2_1
X_10002_ _09941_/A _09941_/B _09942_/Y vssd1 vssd1 vccd1 vccd1 _10093_/A sky130_fd_sc_hd__a21bo_2
X_11953_ _11953_/A _11953_/B vssd1 vssd1 vccd1 vccd1 _11953_/Y sky130_fd_sc_hd__nand2_1
X_10904_ _09156_/Y _10878_/Y _10879_/X _10903_/X vssd1 vssd1 vccd1 vccd1 _10904_/X
+ sky130_fd_sc_hd__a31o_1
X_11884_ _11800_/A _11802_/B _11800_/B vssd1 vssd1 vccd1 vccd1 _11885_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_67_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10835_ _10835_/A _10835_/B _10835_/C vssd1 vssd1 vccd1 vccd1 _10836_/B sky130_fd_sc_hd__or3_1
XANTENNA__10426__B1 _10574_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10766_ hold189/A _11450_/B _10890_/B _11968_/B1 vssd1 vssd1 vccd1 vccd1 _10766_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_109_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12505_ _12669_/B _12506_/B vssd1 vssd1 vccd1 vccd1 _12516_/A sky130_fd_sc_hd__nand2_1
XANTENNA__12179__B1 _09163_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10697_ _10546_/A _10546_/B _10543_/A vssd1 vssd1 vccd1 vccd1 _10701_/A sky130_fd_sc_hd__o21bai_2
XFILLER_0_112_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12436_ reg1_val[31] _07064_/B _09154_/Y vssd1 vssd1 vccd1 vccd1 _12436_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_82_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07101__B _11470_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06940__B _12341_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12367_ fanout13/X _12366_/Y _12365_/X vssd1 vssd1 vccd1 vccd1 _12368_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_10_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09347__A1 _12254_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12298_ reg1_val[28] _12348_/C vssd1 vssd1 vccd1 vccd1 _12298_/Y sky130_fd_sc_hd__xnor2_1
X_11318_ _11318_/A _11421_/A vssd1 vssd1 vccd1 vccd1 _11514_/A sky130_fd_sc_hd__nand2_1
XANTENNA__11558__B _12214_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11249_ _11249_/A _11249_/B _11249_/C vssd1 vssd1 vccd1 vccd1 _11250_/C sky130_fd_sc_hd__or3_1
XANTENNA__07358__B1 _12824_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11154__A1 _10418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11154__B2 _11294_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11574__A _12073_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06790_ reg1_val[3] _11010_/S vssd1 vssd1 vccd1 vccd1 _06791_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_89_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_4_7_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08460_ _08723_/B1 _08732_/A2 _08656_/B _07885_/B vssd1 vssd1 vccd1 vccd1 _08461_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_54_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08391_ _12626_/A _08391_/B _08391_/C vssd1 vssd1 vccd1 vccd1 _08393_/C sky130_fd_sc_hd__and3_1
X_07411_ _11163_/A _07411_/B vssd1 vssd1 vccd1 vccd1 _07413_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_58_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07342_ _09441_/A _07342_/B vssd1 vssd1 vccd1 vccd1 _07349_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_58_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10918__A _11269_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10417__B1 _11294_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08086__B2 _12818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08086__A1 fanout99/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07273_ fanout69/X _10818_/A _08216_/B _10963_/A vssd1 vssd1 vccd1 vccd1 _07274_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_116_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09012_ _09000_/A _09004_/Y _09008_/A _08590_/B _09006_/A vssd1 vssd1 vccd1 vccd1
+ _09013_/B sky130_fd_sc_hd__o2111a_1
XFILLER_0_60_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07011__B _07013_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold100 hold100/A vssd1 vssd1 vccd1 vccd1 hold100/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11749__A _12317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout201_A _12830_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold133 hold133/A vssd1 vssd1 vccd1 vccd1 hold133/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold111 hold111/A vssd1 vssd1 vccd1 vccd1 hold111/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold144 hold144/A vssd1 vssd1 vccd1 vccd1 hold144/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold122 hold122/A vssd1 vssd1 vccd1 vccd1 hold122/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold177 hold177/A vssd1 vssd1 vccd1 vccd1 hold177/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold166 hold299/X vssd1 vssd1 vccd1 vccd1 hold166/X sky130_fd_sc_hd__buf_1
Xhold155 hold155/A vssd1 vssd1 vccd1 vccd1 hold155/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08123__A _08733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold199 hold199/A vssd1 vssd1 vccd1 vccd1 hold199/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold188 hold188/A vssd1 vssd1 vccd1 vccd1 hold188/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09914_ _07510_/A _12366_/B _07036_/X vssd1 vssd1 vccd1 vccd1 _09917_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09845_ _06870_/C _09527_/B _09838_/X _09844_/X vssd1 vssd1 vccd1 vccd1 _09845_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_95_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06988_ _06988_/A _06988_/B vssd1 vssd1 vccd1 vccd1 _12824_/A sky130_fd_sc_hd__xnor2_4
X_09776_ _09556_/A _09556_/B _09553_/A vssd1 vssd1 vccd1 vccd1 _09787_/A sky130_fd_sc_hd__o21ai_2
X_08727_ _11367_/A _08727_/A2 _08727_/B1 _11472_/A vssd1 vssd1 vccd1 vccd1 _08728_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08658_ _08733_/A _08666_/B _08657_/Y vssd1 vssd1 vccd1 vccd1 _08689_/C sky130_fd_sc_hd__a21o_1
Xclkbuf_4_8_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13340_/CLK sky130_fd_sc_hd__clkbuf_8
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07521__B1 _12802_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07609_ _07610_/A _07610_/B vssd1 vssd1 vccd1 vccd1 _07624_/B sky130_fd_sc_hd__nand2_1
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08589_ _08589_/A _08589_/B _08589_/C vssd1 vssd1 vccd1 vccd1 _08590_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_64_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10828__A _11164_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10620_ _10365_/Y _10616_/Y _10619_/Y vssd1 vssd1 vccd1 vccd1 _10620_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__11650__C _11650_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07202__A _10449_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10551_ _10551_/A _10551_/B vssd1 vssd1 vccd1 vccd1 _10597_/A sky130_fd_sc_hd__xor2_2
X_13270_ _13365_/CLK hold22/X vssd1 vssd1 vccd1 vccd1 hold21/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10482_ _10480_/A _10480_/B _10483_/B vssd1 vssd1 vccd1 vccd1 _10482_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_122_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12221_ _12277_/A _12219_/Y _12146_/A _12147_/Y vssd1 vssd1 vccd1 vccd1 _12221_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_121_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06760__B _07080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12152_ _12153_/A _12153_/B vssd1 vssd1 vccd1 vccd1 _12154_/A sky130_fd_sc_hd__or2_1
X_11103_ _10622_/B _11102_/Y _11515_/A vssd1 vssd1 vccd1 vccd1 _11104_/B sky130_fd_sc_hd__a21oi_2
X_12083_ _12084_/A _12084_/B vssd1 vssd1 vccd1 vccd1 _12156_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__11136__A1 _12254_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11034_ _12170_/A _11034_/B vssd1 vssd1 vccd1 vccd1 _11034_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__08552__A2 _12810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12985_ _13013_/A hold190/X vssd1 vssd1 vccd1 vccd1 hold191/A sky130_fd_sc_hd__and2_1
XFILLER_0_115_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11936_ _11936_/A _11936_/B vssd1 vssd1 vccd1 vccd1 _11939_/A sky130_fd_sc_hd__xnor2_1
X_11867_ _11699_/Y _12024_/B _11865_/Y vssd1 vssd1 vccd1 vccd1 _11867_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_0_24_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13061__A1 _11470_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11798_ reg1_val[21] curr_PC[21] vssd1 vssd1 vccd1 vccd1 _11800_/A sky130_fd_sc_hd__or2_1
XFILLER_0_67_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10818_ _10818_/A _12316_/B vssd1 vssd1 vccd1 vccd1 _10820_/B sky130_fd_sc_hd__or2_1
X_10749_ _10748_/A _10748_/B _10748_/C vssd1 vssd1 vccd1 vccd1 _10749_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_55_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12672__B _12673_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12419_ _12419_/A _12419_/B vssd1 vssd1 vccd1 vccd1 _12419_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_11_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07960_ _08030_/A _08030_/B _08030_/C vssd1 vssd1 vccd1 vccd1 _08031_/A sky130_fd_sc_hd__a21o_1
X_06911_ instruction[22] _06921_/B vssd1 vssd1 vccd1 vccd1 _06911_/X sky130_fd_sc_hd__or2_1
XFILLER_0_65_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07891_ fanout75/X _08721_/B1 _08739_/A1 _08304_/B vssd1 vssd1 vccd1 vccd1 _07892_/B
+ sky130_fd_sc_hd__o22a_1
X_06842_ reg1_val[25] _07169_/A vssd1 vssd1 vccd1 vccd1 _06842_/X sky130_fd_sc_hd__and2_1
X_09630_ _09630_/A _09630_/B vssd1 vssd1 vccd1 vccd1 _09643_/A sky130_fd_sc_hd__xor2_4
XANTENNA__07751__B1 _07821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06773_ reg2_val[5] _06771_/A _12429_/B vssd1 vssd1 vccd1 vccd1 _06960_/C sky130_fd_sc_hd__a21o_2
XFILLER_0_65_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09561_ _09456_/A _09456_/B _09453_/A vssd1 vssd1 vccd1 vccd1 _09566_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_77_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08512_ _08517_/A _08517_/B vssd1 vssd1 vccd1 vccd1 _08512_/Y sky130_fd_sc_hd__nand2b_1
X_09492_ _08985_/A _09653_/A _08985_/B vssd1 vssd1 vccd1 vccd1 _09492_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_77_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08443_ _08443_/A _08443_/B vssd1 vssd1 vccd1 vccd1 _08444_/B sky130_fd_sc_hd__nand2_1
XANTENNA__11751__B _12214_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08374_ _08428_/A _08428_/B vssd1 vssd1 vccd1 vccd1 _08374_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_46_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11470__C fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07325_ _07325_/A _07325_/B vssd1 vssd1 vccd1 vccd1 _07398_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__11063__B1 fanout4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07256_ reg1_val[29] _07256_/B vssd1 vssd1 vccd1 vccd1 _07256_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_116_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06580__B _06581_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07187_ _09433_/A _07187_/B vssd1 vssd1 vccd1 vccd1 _07187_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_60_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09828_ _09147_/S _09827_/X _09825_/X vssd1 vssd1 vccd1 vccd1 _09828_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__10322__S _10449_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09759_ _07163_/X fanout7/X _09758_/X _09897_/A vssd1 vssd1 vccd1 vccd1 _09761_/B
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA_fanout64_A _09396_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12770_ reg1_val[29] _12782_/A vssd1 vssd1 vccd1 vccd1 _12772_/A sky130_fd_sc_hd__nand2_1
X_11721_ _11450_/B _11805_/B hold210/A vssd1 vssd1 vccd1 vccd1 _11723_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__06755__B _07089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13043__A1 _08584_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11652_ _11908_/A _11652_/B vssd1 vssd1 vccd1 vccd1 _11657_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_126_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout83 _07208_/Y vssd1 vssd1 vccd1 vccd1 _08507_/B sky130_fd_sc_hd__buf_8
Xfanout72 _09614_/A vssd1 vssd1 vccd1 vccd1 _10575_/A sky130_fd_sc_hd__clkbuf_8
Xfanout50 fanout51/X vssd1 vssd1 vccd1 vccd1 _12067_/A sky130_fd_sc_hd__clkbuf_8
X_10603_ _10603_/A _10603_/B _10603_/C vssd1 vssd1 vccd1 vccd1 _10604_/B sky130_fd_sc_hd__nor3_1
Xfanout61 _12214_/A vssd1 vssd1 vccd1 vccd1 _12150_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_107_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13322_ _13343_/CLK _13322_/D vssd1 vssd1 vccd1 vccd1 hold155/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11583_ _11583_/A _11583_/B vssd1 vssd1 vccd1 vccd1 _11598_/A sky130_fd_sc_hd__and2_1
Xfanout94 _08216_/B vssd1 vssd1 vccd1 vccd1 fanout94/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__06771__A _06771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07273__A2 _10818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10534_ _10490_/A _10490_/B _10488_/Y vssd1 vssd1 vccd1 vccd1 _10615_/A sky130_fd_sc_hd__o21a_2
XFILLER_0_10_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13253_ _13380_/CLK hold28/X vssd1 vssd1 vccd1 vccd1 hold27/A sky130_fd_sc_hd__dfxtp_1
X_10465_ _10465_/A _10465_/B vssd1 vssd1 vccd1 vccd1 _10469_/A sky130_fd_sc_hd__xnor2_1
X_13184_ _13184_/A _13184_/B vssd1 vssd1 vccd1 vccd1 _13184_/Y sky130_fd_sc_hd__xnor2_1
X_10396_ _07089_/A _12404_/A _10394_/Y _10395_/X vssd1 vssd1 vccd1 vccd1 _10396_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_12204_ curr_PC[27] _12204_/B vssd1 vssd1 vccd1 vccd1 _12204_/X sky130_fd_sc_hd__xor2_1
X_12135_ _06881_/X _12132_/X _12134_/Y vssd1 vssd1 vccd1 vccd1 dest_val[25] sky130_fd_sc_hd__o21ai_4
XANTENNA__12857__A1 _12412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12066_ _12066_/A _12066_/B vssd1 vssd1 vccd1 vccd1 _12068_/A sky130_fd_sc_hd__nand2_1
X_11017_ hold287/A _11017_/B vssd1 vssd1 vccd1 vccd1 _11123_/B sky130_fd_sc_hd__or2_1
XANTENNA__07733__B1 _08436_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12968_ hold197/X _13004_/A2 _13016_/B1 hold187/X vssd1 vssd1 vccd1 vccd1 hold235/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12899_ hold55/X hold294/A vssd1 vssd1 vccd1 vccd1 _12899_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_59_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11919_ _12012_/B _11919_/B vssd1 vssd1 vccd1 vccd1 _11936_/A sky130_fd_sc_hd__and2_1
XFILLER_0_117_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07110_ _10574_/A _09768_/A1 _10575_/A _12808_/A vssd1 vssd1 vccd1 vccd1 _07111_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_55_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07264__A2 fanout16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08090_ _08146_/A _08146_/B vssd1 vssd1 vccd1 vccd1 _08098_/A sky130_fd_sc_hd__or2_2
XFILLER_0_27_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07041_ _07041_/A _07041_/B vssd1 vssd1 vccd1 vccd1 _07629_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_2_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08992_ _10105_/B _10106_/A vssd1 vssd1 vccd1 vccd1 _08994_/A sky130_fd_sc_hd__nand2_1
XANTENNA__10931__A _12073_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08401__A _10444_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07943_ _07943_/A _07943_/B vssd1 vssd1 vccd1 vccd1 _07962_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__13019__A _13214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09713__A1 _12808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09713__B2 _12810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07874_ _08728_/A _07874_/B vssd1 vssd1 vccd1 vccd1 _07943_/A sky130_fd_sc_hd__xnor2_2
X_06825_ _11437_/A _06824_/Y _06697_/X vssd1 vssd1 vccd1 vccd1 _11524_/B sky130_fd_sc_hd__a21o_1
X_09613_ _09613_/A _10818_/A vssd1 vssd1 vccd1 vccd1 _09615_/B sky130_fd_sc_hd__or2_1
XFILLER_0_78_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06756_ _06754_/Y _06756_/B vssd1 vssd1 vccd1 vccd1 _10378_/A sky130_fd_sc_hd__nand2b_2
X_09544_ _09481_/A _09481_/B _09479_/X vssd1 vssd1 vccd1 vccd1 _09647_/A sky130_fd_sc_hd__a21oi_4
XFILLER_0_93_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06687_ reg2_val[18] _06720_/B _06703_/B1 _06686_/Y vssd1 vssd1 vccd1 vccd1 _07131_/B
+ sky130_fd_sc_hd__o2bb2a_2
X_09475_ _09292_/A _09292_/B _09290_/Y vssd1 vssd1 vccd1 vccd1 _09476_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_38_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08426_ _08426_/A _08426_/B vssd1 vssd1 vccd1 vccd1 _09023_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_74_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08357_ _09441_/A _08357_/B vssd1 vssd1 vccd1 vccd1 _08364_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_33_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11587__A1 _11472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07308_ _07308_/A _07308_/B vssd1 vssd1 vccd1 vccd1 _07602_/A sky130_fd_sc_hd__or2_2
XANTENNA__07687__A _11908_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08288_ _08288_/A _08288_/B vssd1 vssd1 vccd1 vccd1 _08345_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_104_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07239_ _12846_/A _09236_/B2 _12844_/A _09444_/A vssd1 vssd1 vccd1 vccd1 _07240_/B
+ sky130_fd_sc_hd__o22a_2
X_10250_ _09666_/X _09669_/X _10250_/S vssd1 vssd1 vccd1 vccd1 _10250_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10011__B2 _10941_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10011__A1 fanout59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10181_ _10445_/A _12214_/A fanout59/X _10706_/B2 vssd1 vssd1 vccd1 vccd1 _10182_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_100_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout240 _09147_/S vssd1 vssd1 vccd1 vccd1 _10119_/S sky130_fd_sc_hd__clkbuf_8
XANTENNA__09407__A _10422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout251 _09168_/X vssd1 vssd1 vccd1 vccd1 _12247_/C1 sky130_fd_sc_hd__buf_4
Xfanout273 _12788_/A vssd1 vssd1 vccd1 vccd1 _12791_/A sky130_fd_sc_hd__buf_4
Xfanout262 _12455_/S vssd1 vssd1 vccd1 vccd1 _10780_/A sky130_fd_sc_hd__buf_6
Xfanout295 _13210_/A vssd1 vssd1 vccd1 vccd1 _13214_/A sky130_fd_sc_hd__clkbuf_4
Xfanout284 _06587_/X vssd1 vssd1 vccd1 vccd1 _12611_/A sky130_fd_sc_hd__buf_4
X_12822_ _12822_/A _12830_/B vssd1 vssd1 vccd1 vccd1 _12822_/Y sky130_fd_sc_hd__nand2_1
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12753_ reg1_val[26] _12782_/A vssd1 vssd1 vccd1 vccd1 _12766_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_29_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11704_ _11866_/A _11704_/B vssd1 vssd1 vccd1 vccd1 _11822_/A sky130_fd_sc_hd__xnor2_2
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12684_ _12689_/B _12684_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[11] sky130_fd_sc_hd__and2_4
XFILLER_0_37_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11635_ hold263/A _11635_/B vssd1 vssd1 vccd1 vccd1 _11724_/B sky130_fd_sc_hd__or2_1
XFILLER_0_71_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07246__A2 _10589_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11566_ _11758_/A _11566_/B vssd1 vssd1 vccd1 vccd1 _11568_/B sky130_fd_sc_hd__xor2_1
X_13305_ _13307_/CLK hold227/X vssd1 vssd1 vccd1 vccd1 hold225/A sky130_fd_sc_hd__dfxtp_1
X_10517_ _10513_/Y _10516_/Y _11886_/A vssd1 vssd1 vccd1 vccd1 _10517_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_52_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13236_ hold63/X _13236_/B vssd1 vssd1 vccd1 vccd1 _13236_/Y sky130_fd_sc_hd__nand2_1
X_11497_ _11497_/A _11497_/B vssd1 vssd1 vccd1 vccd1 _11499_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10448_ _10448_/A _10448_/B _10448_/C vssd1 vssd1 vccd1 vccd1 _10449_/C sky130_fd_sc_hd__nand3_1
X_13167_ hold292/X _12789_/B _13166_/X _13246_/B2 vssd1 vssd1 vccd1 vccd1 _13168_/B
+ sky130_fd_sc_hd__a22o_1
X_10379_ _10378_/A _10378_/B _10378_/Y _11624_/A vssd1 vssd1 vccd1 vccd1 _10379_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__07954__B1 _07752_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11847__A _11847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13098_ hold244/A _13097_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13098_/X sky130_fd_sc_hd__mux2_1
X_12118_ _12394_/A _10113_/B _12116_/Y _12117_/X vssd1 vssd1 vccd1 vccd1 _12118_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08221__A _08745_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12049_ _11973_/B _09158_/Y _12049_/S vssd1 vssd1 vccd1 vccd1 _12049_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10491__A_N _10493_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09171__A2 _09167_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06610_ _06612_/B vssd1 vssd1 vccd1 vccd1 _07345_/A sky130_fd_sc_hd__inv_2
X_07590_ _07590_/A _07590_/B vssd1 vssd1 vccd1 vccd1 _07593_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_75_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09260_ _09260_/A _09260_/B _09260_/C vssd1 vssd1 vccd1 vccd1 _09262_/A sky130_fd_sc_hd__or3_1
XFILLER_0_75_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08211_ _08211_/A _08211_/B vssd1 vssd1 vccd1 vccd1 _08213_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_117_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09191_ _07598_/A _07598_/B _07596_/X vssd1 vssd1 vccd1 vccd1 _09302_/A sky130_fd_sc_hd__a21oi_4
XFILLER_0_62_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07237__A2 _08436_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08142_ _08731_/A _08142_/B vssd1 vssd1 vccd1 vccd1 _08169_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_126_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08073_ _08073_/A _08073_/B _08073_/C vssd1 vssd1 vccd1 vccd1 _08075_/A sky130_fd_sc_hd__and3_1
X_07024_ _07050_/A _07050_/C _07223_/B _06960_/C vssd1 vssd1 vccd1 vccd1 _07026_/A
+ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout114_A _12824_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10544__A2 fanout59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11757__A _12073_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09227__A _10707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08975_ _08954_/A _08954_/B _08974_/X vssd1 vssd1 vccd1 vccd1 _08975_/Y sky130_fd_sc_hd__o21ai_1
Xhold26 hold26/A vssd1 vssd1 vccd1 vccd1 hold26/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold15 hold15/A vssd1 vssd1 vccd1 vccd1 hold15/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 hold37/A vssd1 vssd1 vccd1 vccd1 hold37/X sky130_fd_sc_hd__dlygate4sd3_1
X_07926_ _08029_/B vssd1 vssd1 vccd1 vccd1 _07926_/Y sky130_fd_sc_hd__inv_2
Xhold48 hold48/A vssd1 vssd1 vccd1 vccd1 hold48/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 hold59/A vssd1 vssd1 vccd1 vccd1 hold59/X sky130_fd_sc_hd__buf_1
X_07857_ _10927_/A1 _08741_/A2 _08617_/B _11367_/A vssd1 vssd1 vccd1 vccd1 _07858_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__13246__B2 _13246_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06808_ _07149_/A _09351_/B vssd1 vssd1 vccd1 vccd1 _09350_/B sky130_fd_sc_hd__nand2_1
X_07788_ _08745_/A _07788_/B vssd1 vssd1 vccd1 vccd1 _07790_/B sky130_fd_sc_hd__xnor2_2
X_09527_ _09527_/A _09527_/B vssd1 vssd1 vccd1 vccd1 _09527_/X sky130_fd_sc_hd__or2_1
X_06739_ _06805_/A _06702_/A _12680_/B _06738_/X vssd1 vssd1 vccd1 vccd1 _07100_/A
+ sky130_fd_sc_hd__a31o_4
XFILLER_0_93_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09897__A _09897_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08122__B1 _12820_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09458_ _09459_/A _09459_/B vssd1 vssd1 vccd1 vccd1 _09458_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_66_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout27_A _07688_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09389_ _09389_/A _09389_/B vssd1 vssd1 vccd1 vccd1 _09391_/A sky130_fd_sc_hd__xnor2_4
X_08409_ _09433_/A _08409_/B vssd1 vssd1 vccd1 vccd1 _08443_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_46_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11420_ _11420_/A vssd1 vssd1 vccd1 vccd1 _11420_/Y sky130_fd_sc_hd__inv_2
X_11351_ _09172_/B _11338_/X _11345_/X _11350_/Y vssd1 vssd1 vccd1 vccd1 _11351_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__07210__A _07210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06987__A1 _06981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11980__A1 _11707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10302_ _10302_/A _10302_/B vssd1 vssd1 vccd1 vccd1 _10304_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_104_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11282_ _11402_/A _11282_/B vssd1 vssd1 vccd1 vccd1 _11286_/B sky130_fd_sc_hd__or2_1
X_13021_ _13214_/A hold216/X vssd1 vssd1 vccd1 vccd1 hold217/A sky130_fd_sc_hd__and2_1
X_10233_ _09947_/X _10094_/X _10095_/X vssd1 vssd1 vccd1 vccd1 _10233_/X sky130_fd_sc_hd__a21o_1
XANTENNA__10571__A _10571_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11732__A1 _06924_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10164_ _10710_/A _10164_/B _10164_/C vssd1 vssd1 vccd1 vccd1 _10165_/C sky130_fd_sc_hd__nand3_1
XANTENNA__08041__A _08731_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07936__B1 _11751_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10095_ _10096_/A _10096_/B vssd1 vssd1 vccd1 vccd1 _10095_/X sky130_fd_sc_hd__and2_1
XANTENNA__13093__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12498__A _12664_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08361__B1 _08673_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12805_ hold35/X _12818_/B _12804_/Y _13113_/A vssd1 vssd1 vccd1 vccd1 hold36/A sky130_fd_sc_hd__o211a_1
XFILLER_0_57_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10997_ _10909_/X _10996_/Y _12290_/A vssd1 vssd1 vccd1 vccd1 _10997_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_127_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12736_ reg1_val[22] _12741_/B vssd1 vssd1 vccd1 vccd1 _12737_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_127_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12667_ _12666_/A _12663_/Y _12665_/B vssd1 vssd1 vccd1 vccd1 _12671_/A sky130_fd_sc_hd__o21a_2
XFILLER_0_38_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07219__A2 _07220_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11618_ _11618_/A _11618_/B vssd1 vssd1 vccd1 vccd1 _11618_/Y sky130_fd_sc_hd__nor2_1
X_12598_ _12605_/B _12598_/B vssd1 vssd1 vccd1 vccd1 new_PC[22] sky130_fd_sc_hd__xnor2_4
XANTENNA__08216__A _08752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12961__A _13214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11549_ _11519_/Y _11520_/X _11523_/Y _09163_/X _11548_/X vssd1 vssd1 vccd1 vccd1
+ _11549_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_52_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12680__B _12680_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13219_ _13235_/A hold257/X vssd1 vssd1 vccd1 vccd1 _13374_/D sky130_fd_sc_hd__and2_1
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11577__A _12210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11988__A2_N fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_10_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13343_/CLK sky130_fd_sc_hd__clkbuf_8
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08760_ _08761_/A _08761_/B vssd1 vssd1 vccd1 vccd1 _08760_/Y sky130_fd_sc_hd__nor2_1
X_08691_ _08660_/Y _08989_/A _08690_/B vssd1 vssd1 vccd1 vccd1 _08991_/B sky130_fd_sc_hd__a21oi_1
X_07711_ _07712_/A _07712_/B vssd1 vssd1 vccd1 vccd1 _07713_/A sky130_fd_sc_hd__and2_1
XFILLER_0_79_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07155__B2 _12264_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08352__B1 _08564_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07642_ _07642_/A _07642_/B vssd1 vssd1 vccd1 vccd1 _07990_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_88_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09312_ _09088_/X _09096_/X _09351_/B vssd1 vssd1 vccd1 vccd1 _09312_/X sky130_fd_sc_hd__mux2_1
X_07573_ _07573_/A _07573_/B _07573_/C vssd1 vssd1 vccd1 vccd1 _07574_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_48_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout231_A _09669_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06666__B1 _06771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09243_ _09242_/B _09242_/C _09593_/A vssd1 vssd1 vccd1 vccd1 _09245_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_63_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09174_ _09669_/S _09181_/B _09173_/X vssd1 vssd1 vccd1 vccd1 _09176_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_90_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08125_ _08731_/A _08125_/B vssd1 vssd1 vccd1 vccd1 _08130_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_43_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07091__B1 _12810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08056_ _12818_/A _08744_/A2 _08564_/B _12820_/A vssd1 vssd1 vccd1 vccd1 _08057_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_101_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07007_ _07254_/B _07254_/C _07364_/B1 vssd1 vssd1 vccd1 vccd1 _07045_/B sky130_fd_sc_hd__o21ai_2
XFILLER_0_11_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07918__B1 _08617_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08958_ _08958_/A _08958_/B vssd1 vssd1 vccd1 vccd1 _08960_/A sky130_fd_sc_hd__xor2_2
XANTENNA__07146__A1 _09444_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07909_ _07910_/A _07910_/B vssd1 vssd1 vccd1 vccd1 _07981_/B sky130_fd_sc_hd__nand2b_1
X_08889_ _07974_/A _07973_/B _07973_/C vssd1 vssd1 vccd1 vccd1 _08890_/B sky130_fd_sc_hd__a21o_1
XANTENNA__07146__B2 _12848_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10920_ _11180_/A _10920_/B vssd1 vssd1 vccd1 vccd1 _10922_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__10150__B1 _07282_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10851_ _10852_/A _10852_/B vssd1 vssd1 vccd1 vccd1 _10987_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08646__B2 _08646_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08646__A1 _08671_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10782_ _10782_/A _10782_/B vssd1 vssd1 vccd1 vccd1 _10783_/B sky130_fd_sc_hd__and2_1
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12521_ _12530_/A _12521_/B vssd1 vssd1 vccd1 vccd1 _12523_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_93_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06763__B _06799_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12452_ _12453_/A _12453_/B vssd1 vssd1 vccd1 vccd1 _12460_/B sky130_fd_sc_hd__or2_1
XFILLER_0_47_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11403_ _11402_/A _11402_/B _11404_/A vssd1 vssd1 vccd1 vccd1 _11403_/Y sky130_fd_sc_hd__o21ai_1
X_12383_ _12383_/A _12383_/B vssd1 vssd1 vccd1 vccd1 _12383_/X sky130_fd_sc_hd__or2_1
XFILLER_0_34_274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11334_ reg1_val[16] curr_PC[16] vssd1 vssd1 vccd1 vccd1 _11334_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_104_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11265_ _11266_/A _11266_/B vssd1 vssd1 vccd1 vccd1 _11267_/A sky130_fd_sc_hd__nand2_1
X_13004_ hold236/A _13004_/A2 _13006_/B1 hold225/X vssd1 vssd1 vccd1 vccd1 hold226/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10216_ _10078_/A _10077_/B _10075_/Y vssd1 vssd1 vccd1 vccd1 _10221_/A sky130_fd_sc_hd__o21ai_4
XFILLER_0_118_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11196_ _11196_/A _11196_/B _11196_/C vssd1 vssd1 vccd1 vccd1 _11197_/B sky130_fd_sc_hd__or3_1
XFILLER_0_27_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10147_ _10147_/A _10147_/B vssd1 vssd1 vccd1 vccd1 _10149_/A sky130_fd_sc_hd__xor2_1
XANTENNA__07137__A1 _07169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10078_ _10078_/A _10078_/B vssd1 vssd1 vccd1 vccd1 _10079_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_89_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07115__A _09716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06954__A _10710_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12719_ _12725_/A _12725_/B _12741_/B _06997_/C vssd1 vssd1 vccd1 vccd1 _12720_/B
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_84_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12197__A1 _07140_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10747__A2 _10782_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07073__B1 _07074_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09930_ _09931_/A _09931_/B vssd1 vssd1 vccd1 vccd1 _09930_/X sky130_fd_sc_hd__and2_1
XFILLER_0_111_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11100__A _11100_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09861_ _12076_/A _09861_/B vssd1 vssd1 vccd1 vccd1 _09863_/B sky130_fd_sc_hd__xnor2_1
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09792_ _09630_/A _09630_/B _09629_/A vssd1 vssd1 vccd1 vccd1 _09802_/A sky130_fd_sc_hd__a21o_2
X_08812_ _08811_/A _08811_/C _08811_/B vssd1 vssd1 vccd1 vccd1 _08813_/C sky130_fd_sc_hd__a21o_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08743_ _08743_/A _08743_/B vssd1 vssd1 vccd1 vccd1 _08746_/B sky130_fd_sc_hd__xor2_1
XANTENNA_fanout279_A _12790_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout181_A _12798_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08674_ _09445_/A _08678_/B vssd1 vssd1 vccd1 vccd1 _08677_/B sky130_fd_sc_hd__or2_1
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07625_ _07627_/A _07625_/B vssd1 vssd1 vccd1 vccd1 _08917_/B sky130_fd_sc_hd__or2_1
XFILLER_0_119_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06864__A _07149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07556_ _07556_/A _07556_/B vssd1 vssd1 vccd1 vccd1 _07558_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07487_ _07487_/A _07487_/B vssd1 vssd1 vccd1 vccd1 _07491_/A sky130_fd_sc_hd__xor2_1
X_09226_ _10445_/A _12834_/A _12836_/A _10706_/B2 vssd1 vssd1 vccd1 vccd1 _09227_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_32_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09157_ _09163_/A _09157_/B vssd1 vssd1 vccd1 vccd1 _09157_/X sky130_fd_sc_hd__or2_1
XFILLER_0_32_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10199__B1 _10575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09088_ reg1_val[3] reg1_val[28] _09108_/S vssd1 vssd1 vccd1 vccd1 _09088_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_31_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08108_ _08108_/A _08108_/B vssd1 vssd1 vccd1 vccd1 _08110_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_101_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08039_ _07226_/A _07226_/B _07149_/A vssd1 vssd1 vccd1 vccd1 _08041_/C sky130_fd_sc_hd__a21o_2
XFILLER_0_4_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout94_A _08216_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11050_ _10570_/A _12213_/A fanout56/X _10571_/A vssd1 vssd1 vccd1 vccd1 _11051_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12360__B2 _09142_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10001_ _09946_/A _09946_/B _09944_/X vssd1 vssd1 vccd1 vccd1 _10096_/A sky130_fd_sc_hd__a21oi_4
X_11952_ _11874_/B _11875_/A _11874_/A vssd1 vssd1 vccd1 vccd1 _11953_/B sky130_fd_sc_hd__o21ai_1
X_10903_ _09152_/Y _10883_/Y _10889_/Y _09172_/B _10902_/X vssd1 vssd1 vccd1 vccd1
+ _10903_/X sky130_fd_sc_hd__a221o_1
X_11883_ _11883_/A _11883_/B vssd1 vssd1 vccd1 vccd1 _11885_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_39_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10834_ _10835_/A _10835_/B _10835_/C vssd1 vssd1 vccd1 vccd1 _10976_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_94_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10426__A1 _10574_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10426__B2 _10575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10765_ _11633_/B _10890_/B hold189/A vssd1 vssd1 vccd1 vccd1 _10765_/Y sky130_fd_sc_hd__a21oi_1
X_12504_ reg1_val[9] curr_PC[9] _12622_/S vssd1 vssd1 vccd1 vccd1 _12506_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_82_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10296__A _10448_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10696_ _10844_/A _10683_/Y _10695_/C vssd1 vssd1 vccd1 vccd1 _10702_/B sky130_fd_sc_hd__o21ba_1
X_12435_ hold118/A _12435_/B vssd1 vssd1 vccd1 vccd1 _12435_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_120_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12366_ fanout6/X _12366_/B vssd1 vssd1 vccd1 vccd1 _12366_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__11839__B _11839_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11317_ _11098_/A _11209_/X _11211_/B vssd1 vssd1 vccd1 vccd1 _11317_/Y sky130_fd_sc_hd__a21oi_1
X_12297_ _12243_/A _12240_/Y _12242_/B vssd1 vssd1 vccd1 vccd1 _12348_/C sky130_fd_sc_hd__o21ai_2
XFILLER_0_120_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11248_ _12254_/A1 _11234_/B _11247_/X _09111_/S vssd1 vssd1 vccd1 vccd1 _11249_/C
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__07358__A1 _12826_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08555__B1 _08673_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12351__A1 _12394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07358__B2 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11179_ _10574_/A _11989_/A _12067_/A _10575_/A vssd1 vssd1 vccd1 vccd1 _11180_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11154__A2 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06949__A _10710_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06668__B _07220_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08307__B1 _08656_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13064__C1 _13128_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08390_ _07067_/A _07067_/B _08038_/A vssd1 vssd1 vccd1 vccd1 _08393_/B sky130_fd_sc_hd__a21oi_1
X_07410_ _12826_/A fanout74/X _10948_/B2 _12828_/A vssd1 vssd1 vccd1 vccd1 _07411_/B
+ sky130_fd_sc_hd__o22a_1
X_07341_ _12846_/A _09440_/B1 _12844_/A _09238_/B vssd1 vssd1 vccd1 vccd1 _07342_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_85_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12811__C1 _13128_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08086__A2 _08741_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07272_ _07107_/A _07107_/B _07309_/B vssd1 vssd1 vccd1 vccd1 _07272_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_0_116_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09011_ _08542_/Y _08703_/B _08544_/B vssd1 vssd1 vccd1 vccd1 _09013_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_14_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold101 hold101/A vssd1 vssd1 vccd1 vccd1 hold101/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold112 hold112/A vssd1 vssd1 vccd1 vccd1 hold112/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold134 hold134/A vssd1 vssd1 vccd1 vccd1 hold134/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold123 hold123/A vssd1 vssd1 vccd1 vccd1 hold123/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08404__A _08722_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold167 hold167/A vssd1 vssd1 vccd1 vccd1 hold167/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold156 hold156/A vssd1 vssd1 vccd1 vccd1 hold156/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold145 hold145/A vssd1 vssd1 vccd1 vccd1 hold145/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold178 hold178/A vssd1 vssd1 vccd1 vccd1 hold178/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold189 hold189/A vssd1 vssd1 vccd1 vccd1 hold189/X sky130_fd_sc_hd__dlygate4sd3_1
X_09913_ _09913_/A _09913_/B vssd1 vssd1 vccd1 vccd1 _09927_/A sky130_fd_sc_hd__xnor2_1
X_09844_ _12394_/A _06924_/X _09843_/Y _12403_/A1 _06782_/Y vssd1 vssd1 vccd1 vccd1
+ _09844_/X sky130_fd_sc_hd__o32a_1
XFILLER_0_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06987_ _06981_/A _11020_/A _07074_/A _07074_/C _07074_/B vssd1 vssd1 vccd1 vccd1
+ _06988_/B sky130_fd_sc_hd__o41a_2
X_09775_ _09775_/A _09775_/B vssd1 vssd1 vccd1 vccd1 _09789_/A sky130_fd_sc_hd__xnor2_1
X_08726_ _08726_/A _08726_/B vssd1 vssd1 vccd1 vccd1 _08738_/A sky130_fd_sc_hd__xnor2_1
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08657_ _08666_/A _08666_/B vssd1 vssd1 vccd1 vccd1 _08657_/Y sky130_fd_sc_hd__nor2_1
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07521__B2 fanout30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07521__A1 _07688_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07608_ _11261_/A _07608_/B vssd1 vssd1 vccd1 vccd1 _07610_/B sky130_fd_sc_hd__xnor2_1
X_08588_ _08589_/B _08589_/C _08589_/A vssd1 vssd1 vccd1 vccd1 _09004_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_119_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07539_ _07540_/A _07540_/B _07540_/C _07540_/D vssd1 vssd1 vccd1 vccd1 _09212_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_36_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07285__B1 _08436_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10550_ _10551_/B _10551_/A vssd1 vssd1 vccd1 vccd1 _10720_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_107_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09209_ _09209_/A _09209_/B vssd1 vssd1 vccd1 vccd1 _09214_/A sky130_fd_sc_hd__nand2_2
X_10481_ _10342_/A _10342_/B _10340_/Y vssd1 vssd1 vccd1 vccd1 _10483_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_17_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12220_ _12146_/A _12147_/Y _12277_/A _12219_/Y vssd1 vssd1 vccd1 vccd1 _12277_/B
+ sky130_fd_sc_hd__a211oi_2
X_12151_ _12214_/C _12151_/B vssd1 vssd1 vccd1 vccd1 _12153_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_20_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11102_ _11102_/A _11102_/B _11320_/A vssd1 vssd1 vccd1 vccd1 _11102_/Y sky130_fd_sc_hd__nor3_1
X_12082_ _12156_/A _12082_/B vssd1 vssd1 vccd1 vccd1 _12084_/B sky130_fd_sc_hd__and2_1
XANTENNA__11136__A2 _11121_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11033_ _11033_/A _11033_/B _11033_/C _11033_/D vssd1 vssd1 vccd1 vccd1 _11034_/B
+ sky130_fd_sc_hd__or4_2
XANTENNA__11541__C1 _12307_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12984_ hold189/X _13004_/A2 _13006_/B1 _13295_/Q vssd1 vssd1 vccd1 vccd1 hold190/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11935_ _11936_/A _11936_/B vssd1 vssd1 vccd1 vccd1 _11935_/X sky130_fd_sc_hd__and2_1
XFILLER_0_86_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11866_ _11866_/A _12098_/A vssd1 vssd1 vccd1 vccd1 _12024_/B sky130_fd_sc_hd__nand2_1
XANTENNA__13061__A2 _13087_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11797_ _11797_/A _11797_/B vssd1 vssd1 vccd1 vccd1 _11797_/Y sky130_fd_sc_hd__xnor2_1
X_10817_ _10680_/A _10680_/B _10677_/A vssd1 vssd1 vccd1 vccd1 _10820_/A sky130_fd_sc_hd__a21o_1
X_10748_ _10748_/A _10748_/B _10748_/C vssd1 vssd1 vccd1 vccd1 _10748_/X sky130_fd_sc_hd__or3_1
XFILLER_0_54_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12418_ _12372_/A _12371_/Y _12418_/S vssd1 vssd1 vccd1 vccd1 _12419_/B sky130_fd_sc_hd__mux2_1
X_10679_ _11269_/A _10679_/B vssd1 vssd1 vccd1 vccd1 _10680_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_112_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08224__A _08742_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12349_ reg1_val[28] _12348_/C reg1_val[29] vssd1 vssd1 vccd1 vccd1 _12349_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_121_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06910_ instruction[14] _06884_/Y _06909_/X _06634_/B vssd1 vssd1 vccd1 vccd1 reg1_idx[3]
+ sky130_fd_sc_hd__o211a_4
XFILLER_0_49_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_32 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07890_ _07890_/A _07890_/B vssd1 vssd1 vccd1 vccd1 _07915_/A sky130_fd_sc_hd__nor2_1
XANTENNA__10335__B1 _11171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06841_ reg1_val[26] _07140_/B vssd1 vssd1 vccd1 vccd1 _06841_/X sky130_fd_sc_hd__and2_1
XANTENNA__07751__A1 _07033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06772_ reg2_val[5] _06720_/B _12429_/B vssd1 vssd1 vccd1 vccd1 _06774_/B sky130_fd_sc_hd__a21oi_4
X_09560_ _09560_/A _09560_/B vssd1 vssd1 vccd1 vccd1 _09630_/A sky130_fd_sc_hd__xor2_4
X_09491_ _09376_/X _09542_/C _09490_/Y vssd1 vssd1 vccd1 vccd1 _09491_/X sky130_fd_sc_hd__a21o_1
X_08511_ _08519_/A _08519_/B _08505_/X vssd1 vssd1 vccd1 vccd1 _08517_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_77_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08442_ _08442_/A _08442_/B _08442_/C vssd1 vssd1 vccd1 vccd1 _08474_/A sky130_fd_sc_hd__or3_2
XFILLER_0_93_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_450 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07261__B1_N _10928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08373_ _08373_/A _08373_/B vssd1 vssd1 vccd1 vccd1 _08428_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_128_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07324_ _07233_/A _07233_/B _07231_/Y vssd1 vssd1 vccd1 vccd1 _07398_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_46_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12260__B1 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11063__A1 _11294_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11063__B2 _11146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07255_ reg1_val[28] _07254_/B _07254_/C _12765_/B _07364_/B1 vssd1 vssd1 vccd1 vccd1
+ _07256_/B sky130_fd_sc_hd__o41a_1
XFILLER_0_121_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10664__A _10664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07186_ _09441_/A _07188_/B vssd1 vssd1 vccd1 vccd1 _07187_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_41_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09827_ _09680_/X _10880_/B _11118_/A vssd1 vssd1 vccd1 vccd1 _09827_/X sky130_fd_sc_hd__mux2_1
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09758_ _09758_/A fanout7/X vssd1 vssd1 vccd1 vccd1 _09758_/X sky130_fd_sc_hd__or2_1
XFILLER_0_69_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08709_ _08490_/Y _08707_/A _08707_/B _08708_/X _09018_/A vssd1 vssd1 vccd1 vccd1
+ _08711_/B sky130_fd_sc_hd__a311o_1
XANTENNA__11826__B1 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11720_ hold177/A _11720_/B vssd1 vssd1 vccd1 vccd1 _11805_/B sky130_fd_sc_hd__or2_1
X_09689_ _10391_/A2 _09688_/X hold234/A vssd1 vssd1 vccd1 vccd1 _09689_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__09495__A1 _11118_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout40 _07226_/X vssd1 vssd1 vccd1 vccd1 _12836_/A sky130_fd_sc_hd__buf_4
XFILLER_0_37_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11651_ _09613_/A _12316_/A fanout12/X _09614_/A vssd1 vssd1 vccd1 vccd1 _11652_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_76_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout73 _09400_/A vssd1 vssd1 vccd1 vccd1 _09614_/A sky130_fd_sc_hd__clkbuf_8
Xfanout62 _12846_/A vssd1 vssd1 vccd1 vccd1 _12214_/A sky130_fd_sc_hd__clkbuf_8
Xfanout51 _12844_/A vssd1 vssd1 vccd1 vccd1 fanout51/X sky130_fd_sc_hd__clkbuf_8
X_11582_ _11582_/A _11582_/B vssd1 vssd1 vccd1 vccd1 _11583_/B sky130_fd_sc_hd__nand2_1
X_10602_ _10603_/A _10603_/B _10603_/C vssd1 vssd1 vccd1 vccd1 _10604_/A sky130_fd_sc_hd__o21a_1
X_13321_ _13343_/CLK _13321_/D vssd1 vssd1 vccd1 vccd1 hold148/A sky130_fd_sc_hd__dfxtp_1
X_10533_ _10410_/Y _10500_/Y _11792_/A vssd1 vssd1 vccd1 vccd1 _10624_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_52_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout84 _12830_/A vssd1 vssd1 vccd1 vccd1 _11472_/A sky130_fd_sc_hd__buf_8
XFILLER_0_37_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout95 _07076_/Y vssd1 vssd1 vccd1 vccd1 _08216_/B sky130_fd_sc_hd__buf_8
XFILLER_0_122_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10574__A _10574_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13252_ _13383_/CLK _13252_/D vssd1 vssd1 vccd1 vccd1 hold132/A sky130_fd_sc_hd__dfxtp_1
X_10464_ _11269_/A _10464_/B vssd1 vssd1 vccd1 vccd1 _10465_/B sky130_fd_sc_hd__xor2_1
XANTENNA__08044__A _08598_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13183_ _13235_/A _13183_/B vssd1 vssd1 vccd1 vccd1 _13366_/D sky130_fd_sc_hd__and2_1
X_10395_ hold273/A _09835_/B _10393_/X _09837_/A vssd1 vssd1 vccd1 vccd1 _10395_/X
+ sky130_fd_sc_hd__a31o_1
X_12203_ _12455_/S _12204_/B _12202_/Y _12200_/X vssd1 vssd1 vccd1 vccd1 dest_val[26]
+ sky130_fd_sc_hd__o31ai_4
XFILLER_0_32_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07430__B1 _09568_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08979__A _12423_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12134_ curr_PC[25] _12201_/C _12133_/Y vssd1 vssd1 vccd1 vccd1 _12134_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__07883__A _08722_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12857__A2 _13087_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12065_ _12065_/A _12065_/B vssd1 vssd1 vccd1 vccd1 _12066_/B sky130_fd_sc_hd__or2_1
X_11016_ hold212/A _11633_/B _11127_/B _11968_/B1 vssd1 vssd1 vccd1 vccd1 _11016_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__07733__A1 _08304_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07733__B2 fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12967_ _13214_/A hold198/X vssd1 vssd1 vccd1 vccd1 hold199/A sky130_fd_sc_hd__and2_1
XFILLER_0_87_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12898_ hold273/X hold7/X vssd1 vssd1 vccd1 vccd1 _13129_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__07497__B1 _09442_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08219__A _08733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11918_ _11918_/A _11918_/B vssd1 vssd1 vccd1 vccd1 _11919_/B sky130_fd_sc_hd__or2_1
XANTENNA__13034__A2 _06572_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07123__A _09343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11849_ _11931_/B _11849_/B vssd1 vssd1 vccd1 vccd1 _11853_/A sky130_fd_sc_hd__and2_1
XFILLER_0_27_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12793__A1 _12264_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07040_ _07041_/A _07041_/B vssd1 vssd1 vccd1 vccd1 _07040_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_30_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07421__B1 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08991_ _08991_/A _08991_/B vssd1 vssd1 vccd1 vccd1 _10106_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__10308__B1 _07282_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07942_ _07964_/A _07964_/B vssd1 vssd1 vccd1 vccd1 _07942_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__09713__A2 fanout16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07873_ _08727_/A2 _11751_/A _11766_/A _08727_/B1 vssd1 vssd1 vccd1 vccd1 _07874_/B
+ sky130_fd_sc_hd__o22a_1
X_06824_ _11332_/A _06823_/X _06704_/Y vssd1 vssd1 vccd1 vccd1 _06824_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__11520__A2 _11649_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09612_ _09611_/B _09611_/C _09746_/A vssd1 vssd1 vccd1 vccd1 _09618_/B sky130_fd_sc_hd__a21oi_1
X_09543_ _09543_/A _10275_/A vssd1 vssd1 vccd1 vccd1 _09853_/A sky130_fd_sc_hd__nand2_1
X_06755_ reg1_val[8] _07089_/A vssd1 vssd1 vccd1 vccd1 _06756_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_92_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06686_ _06686_/A _12639_/B vssd1 vssd1 vccd1 vccd1 _06686_/Y sky130_fd_sc_hd__nor2_1
X_09474_ _09474_/A _09474_/B vssd1 vssd1 vccd1 vccd1 _09476_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_78_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07488__B1 _10948_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08425_ _08426_/A _08426_/B vssd1 vssd1 vccd1 vccd1 _08425_/X sky130_fd_sc_hd__or2_1
XANTENNA__07033__A _07033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09659__S _09666_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08356_ _12810_/A _09238_/B _09440_/B1 _08739_/A1 vssd1 vssd1 vccd1 vccd1 _08357_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_74_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07307_ _07674_/A _07674_/B vssd1 vssd1 vccd1 vccd1 _07308_/B sky130_fd_sc_hd__and2b_1
XANTENNA__11587__A2 _12214_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08287_ _08287_/A _08287_/B vssd1 vssd1 vccd1 vccd1 _08345_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_6_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07238_ _09442_/A _07238_/B vssd1 vssd1 vccd1 vccd1 _07241_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_61_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07169_ _07169_/A _07169_/B vssd1 vssd1 vccd1 vccd1 _07169_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_14_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08799__A _11758_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10011__A2 _10589_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10180_ _10070_/B _10073_/B _10070_/A vssd1 vssd1 vccd1 vccd1 _10194_/A sky130_fd_sc_hd__o21ba_1
Xfanout241 _09147_/S vssd1 vssd1 vccd1 vccd1 _10252_/S sky130_fd_sc_hd__clkbuf_4
Xfanout230 _09505_/S vssd1 vssd1 vccd1 vccd1 _09666_/S sky130_fd_sc_hd__buf_6
Xfanout274 _06572_/Y vssd1 vssd1 vccd1 vccd1 _12788_/A sky130_fd_sc_hd__buf_4
Xfanout263 _12455_/S vssd1 vssd1 vccd1 vccd1 _12448_/S sky130_fd_sc_hd__buf_4
Xfanout252 _12428_/A vssd1 vssd1 vccd1 vccd1 _11876_/A sky130_fd_sc_hd__buf_4
Xfanout296 _06578_/Y vssd1 vssd1 vccd1 vccd1 _13210_/A sky130_fd_sc_hd__buf_2
Xfanout285 _06587_/X vssd1 vssd1 vccd1 vccd1 _12741_/B sky130_fd_sc_hd__buf_8
X_12821_ hold43/X _12818_/B _12820_/Y _13245_/A vssd1 vssd1 vccd1 vccd1 hold44/A sky130_fd_sc_hd__o211a_1
XFILLER_0_88_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06766__B _07036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07479__B1 _10022_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12752_ _12752_/A _12754_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[25] sky130_fd_sc_hd__xnor2_4
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12683_ _12683_/A _12683_/B _12683_/C vssd1 vssd1 vccd1 vccd1 _12684_/B sky130_fd_sc_hd__nand3_1
X_11703_ _11323_/B _11702_/Y _12026_/B vssd1 vssd1 vccd1 vccd1 _11704_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_127_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11634_ _11633_/B _11720_/B hold177/A vssd1 vssd1 vccd1 vccd1 _11634_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__11027__A1 _09156_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11565_ _11653_/A fanout12/X fanout8/X _08752_/B vssd1 vssd1 vccd1 vccd1 _11566_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10786__B1 _10571_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13304_ _13307_/CLK _13304_/D vssd1 vssd1 vccd1 vccd1 hold236/A sky130_fd_sc_hd__dfxtp_1
X_10516_ _10516_/A vssd1 vssd1 vccd1 vccd1 _10516_/Y sky130_fd_sc_hd__inv_2
X_11496_ _11497_/A _11497_/B vssd1 vssd1 vccd1 vccd1 _11496_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13235_ _13235_/A hold110/X vssd1 vssd1 vccd1 vccd1 _13378_/D sky130_fd_sc_hd__and2_1
X_10447_ _10448_/B _10448_/C _10448_/A vssd1 vssd1 vccd1 vccd1 _10449_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_20_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13166_ hold271/X _13165_/Y fanout2/A vssd1 vssd1 vccd1 vccd1 _13166_/X sky130_fd_sc_hd__mux2_1
X_10378_ _10378_/A _10378_/B vssd1 vssd1 vccd1 vccd1 _10378_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__07954__A1 _07099_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11847__B _12214_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13097_ _13097_/A _13097_/B vssd1 vssd1 vccd1 vccd1 _13097_/Y sky130_fd_sc_hd__xnor2_1
X_12117_ _12112_/Y _12113_/Y _12115_/X _12244_/S vssd1 vssd1 vccd1 vccd1 _12117_/X
+ sky130_fd_sc_hd__o31a_1
X_12048_ hold254/A _11636_/B _12119_/B _12047_/Y _12247_/C1 vssd1 vssd1 vccd1 vccd1
+ _12048_/X sky130_fd_sc_hd__a311o_1
XFILLER_0_46_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06957__A _12341_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12215__A0 _12213_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08210_ _08210_/A _08210_/B vssd1 vssd1 vccd1 vccd1 _08211_/B sky130_fd_sc_hd__xor2_1
XANTENNA__07788__A _08745_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09190_ _09542_/A _12426_/B _12426_/C _12426_/A vssd1 vssd1 vccd1 vccd1 _09190_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_62_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08141_ _08730_/A1 _11367_/A _08038_/A _10927_/A1 vssd1 vssd1 vccd1 vccd1 _08142_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_102_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11974__C1 _12307_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08072_ _08072_/A _08072_/B vssd1 vssd1 vccd1 vccd1 _08073_/C sky130_fd_sc_hd__xor2_1
XFILLER_0_102_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07023_ _12341_/A _07064_/B _09147_/S vssd1 vssd1 vccd1 vccd1 _07023_/X sky130_fd_sc_hd__and3_1
XFILLER_0_3_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09395__B1 _11146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08974_ _08939_/A _08939_/B _08954_/A _08954_/B vssd1 vssd1 vccd1 vccd1 _08974_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold16 hold16/A vssd1 vssd1 vccd1 vccd1 hold16/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold38 hold38/A vssd1 vssd1 vccd1 vccd1 hold38/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold27 hold27/A vssd1 vssd1 vccd1 vccd1 hold27/X sky130_fd_sc_hd__dlygate4sd3_1
X_07925_ _08745_/A _07925_/B vssd1 vssd1 vccd1 vccd1 _08029_/B sky130_fd_sc_hd__xnor2_1
Xhold49 hold49/A vssd1 vssd1 vccd1 vccd1 hold49/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09698__B2 _09111_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09698__A1 _09152_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07856_ _07856_/A _07856_/B vssd1 vssd1 vccd1 vccd1 _07878_/A sky130_fd_sc_hd__xor2_1
XANTENNA__13246__A2 _06892_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06807_ reg2_val[0] _06720_/B _06702_/A _06805_/X vssd1 vssd1 vccd1 vccd1 _09311_/S
+ sky130_fd_sc_hd__a22o_1
X_07787_ _08732_/A1 _08744_/A2 _08564_/B _10927_/A1 vssd1 vssd1 vccd1 vccd1 _07788_/B
+ sky130_fd_sc_hd__o22a_1
X_09526_ _09527_/A _09525_/B _11624_/A vssd1 vssd1 vccd1 vccd1 _09526_/X sky130_fd_sc_hd__a21o_1
X_06738_ reg2_val[10] _06799_/B vssd1 vssd1 vccd1 vccd1 _06738_/X sky130_fd_sc_hd__and2_1
XFILLER_0_78_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09457_ _09459_/A _09459_/B vssd1 vssd1 vccd1 vccd1 _09457_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_39_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08122__A1 _08741_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08122__B2 _08732_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06669_ _11727_/A _06669_/B vssd1 vssd1 vccd1 vccd1 _06676_/C sky130_fd_sc_hd__nor2_2
X_08408_ _12804_/A _08741_/A2 _08617_/B _08723_/B1 vssd1 vssd1 vccd1 vccd1 _08409_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_19_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09388_ _11673_/A _09388_/B vssd1 vssd1 vccd1 vccd1 _09389_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__12206__B1 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08339_ _08342_/A _08342_/B vssd1 vssd1 vccd1 vccd1 _08343_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_117_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11350_ _10113_/A _11234_/B _11349_/X vssd1 vssd1 vccd1 vccd1 _11350_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_104_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06987__A2 _11020_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10301_ _10302_/A _10302_/B vssd1 vssd1 vccd1 vccd1 _10480_/A sky130_fd_sc_hd__nor2_1
X_13020_ _13312_/Q _13213_/B2 _13213_/A2 hold215/X vssd1 vssd1 vccd1 vccd1 hold216/A
+ sky130_fd_sc_hd__a22o_1
X_11281_ _11280_/B _11281_/B vssd1 vssd1 vccd1 vccd1 _11282_/B sky130_fd_sc_hd__and2b_1
XANTENNA__13182__B2 _12790_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10232_ _10232_/A _10368_/A _10496_/A _10617_/A vssd1 vssd1 vccd1 vccd1 _10232_/X
+ sky130_fd_sc_hd__or4_1
XANTENNA__10571__B _10571_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07936__A1 _08727_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10163_ _10164_/B _10164_/C _10710_/A vssd1 vssd1 vccd1 vccd1 _10165_/B sky130_fd_sc_hd__a21o_1
XANTENNA__07936__B2 _08727_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10094_ _10096_/A _10096_/B vssd1 vssd1 vccd1 vccd1 _10094_/X sky130_fd_sc_hd__or2_1
XFILLER_0_107_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08361__A1 _08436_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13237__A2 _13246_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09153__A _12174_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08361__B2 fanout99/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11248__B2 _09111_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12804_ _12804_/A _12818_/B vssd1 vssd1 vccd1 vccd1 _12804_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_97_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10996_ _10996_/A _10996_/B vssd1 vssd1 vccd1 vccd1 _10996_/Y sky130_fd_sc_hd__nand2_2
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12735_ reg1_val[22] _12741_/B vssd1 vssd1 vccd1 vccd1 _12737_/A sky130_fd_sc_hd__or2_1
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12666_ _12666_/A _12666_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[8] sky130_fd_sc_hd__xor2_4
X_12597_ _12584_/Y _12605_/C _12607_/B vssd1 vssd1 vccd1 vccd1 _12598_/B sky130_fd_sc_hd__o21ai_4
XFILLER_0_65_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11617_ _11874_/A _11616_/B _11616_/C vssd1 vssd1 vccd1 vccd1 _11618_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_37_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11548_ _11527_/Y _11528_/X _11535_/X _11547_/X vssd1 vssd1 vccd1 vccd1 _11548_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__08216__B _08216_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_275 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xmax_cap238 _07044_/A vssd1 vssd1 vccd1 vccd1 _11118_/A sky130_fd_sc_hd__buf_4
X_11479_ _11479_/A _11479_/B vssd1 vssd1 vccd1 vccd1 _11489_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13218_ hold256/X _12789_/B _13217_/X _12790_/A vssd1 vssd1 vccd1 vccd1 hold257/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13149_ _12889_/X _13149_/B vssd1 vssd1 vccd1 vccd1 _13150_/B sky130_fd_sc_hd__nand2b_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07047__C_N _11172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07710_ _11758_/A _07710_/B vssd1 vssd1 vccd1 vccd1 _07712_/B sky130_fd_sc_hd__xnor2_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08690_ _08690_/A _08690_/B vssd1 vssd1 vccd1 vccd1 _08989_/B sky130_fd_sc_hd__nor2_1
XANTENNA__08352__A1 _07955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08352__B2 _07896_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07641_ _11908_/A _07641_/B vssd1 vssd1 vccd1 vccd1 _07642_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__11239__A1 _08980_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07572_ _07573_/A _07573_/B _07573_/C vssd1 vssd1 vccd1 vccd1 _07574_/A sky130_fd_sc_hd__o21a_1
X_09311_ _09085_/X _09089_/X _09311_/S vssd1 vssd1 vccd1 vccd1 _09311_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_88_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09852__A1 _11142_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10937__A _12076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09242_ _09593_/A _09242_/B _09242_/C vssd1 vssd1 vccd1 vccd1 _09245_/A sky130_fd_sc_hd__and3_1
XANTENNA__07863__B1 _08564_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09173_ _09131_/X _09181_/B _09351_/B vssd1 vssd1 vccd1 vccd1 _09173_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_28_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07615__B1 _08507_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08124_ _11367_/A _08038_/A _11472_/A _08730_/A1 vssd1 vssd1 vccd1 vccd1 _08125_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_114_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07091__B2 _08752_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07091__A1 _12808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10672__A _11470_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08055_ _08055_/A _08055_/B vssd1 vssd1 vccd1 vccd1 _08058_/B sky130_fd_sc_hd__xor2_1
XANTENNA__09238__A _10941_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07006_ _09666_/S _07006_/B vssd1 vssd1 vccd1 vccd1 _07006_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_12_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08142__A _08731_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07918__A1 _08732_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07918__B2 _10927_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08040__B1 _08731_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13194__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08957_ _08946_/A _08946_/B _08947_/Y vssd1 vssd1 vccd1 vccd1 _08962_/A sky130_fd_sc_hd__o21ai_2
X_07908_ _07908_/A _07908_/B vssd1 vssd1 vccd1 vccd1 _07910_/B sky130_fd_sc_hd__xnor2_1
X_08888_ _08876_/A _08876_/B _08877_/Y vssd1 vssd1 vccd1 vccd1 _08895_/A sky130_fd_sc_hd__o21ai_2
XANTENNA__07146__A2 _12846_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07839_ _07818_/B _07818_/C _07818_/A vssd1 vssd1 vccd1 vccd1 _07840_/C sky130_fd_sc_hd__o21ai_1
XANTENNA__10150__A1 _10567_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10150__B2 _10664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10850_ _10850_/A _10850_/B vssd1 vssd1 vccd1 vccd1 _10852_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_94_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09509_ _09365_/X _09508_/X _09974_/A vssd1 vssd1 vccd1 vccd1 _09509_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_93_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08646__A2 _08661_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10781_ _10780_/A _10777_/X _10778_/X _10780_/Y vssd1 vssd1 vccd1 vccd1 dest_val[11]
+ sky130_fd_sc_hd__a22o_4
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12520_ _12680_/B _12520_/B vssd1 vssd1 vccd1 vccd1 _12521_/B sky130_fd_sc_hd__or2_1
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12451_ _12460_/A _12451_/B vssd1 vssd1 vccd1 vccd1 _12453_/B sky130_fd_sc_hd__nand2_1
XANTENNA__07221__A _08038_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11402_ _11402_/A _11402_/B vssd1 vssd1 vccd1 vccd1 _11404_/B sky130_fd_sc_hd__nor2_1
X_12382_ _12413_/B _12382_/B vssd1 vssd1 vccd1 vccd1 _12382_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_0_34_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11333_ _11226_/Y _11230_/B _11228_/B vssd1 vssd1 vccd1 vccd1 _11337_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_50_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10582__A _11261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09148__A _12626_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11264_ _11394_/A _11264_/B vssd1 vssd1 vccd1 vccd1 _11266_/B sky130_fd_sc_hd__nor2_1
XANTENNA__08052__A _08742_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13003_ _13009_/A hold237/X vssd1 vssd1 vccd1 vccd1 _13304_/D sky130_fd_sc_hd__and2_1
XANTENNA__12363__C1 _12455_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10215_ _10079_/A _10079_/B _10062_/A vssd1 vssd1 vccd1 vccd1 _10225_/A sky130_fd_sc_hd__a21o_2
X_11195_ _11196_/A _11196_/B _11196_/C vssd1 vssd1 vccd1 vccd1 _11197_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_118_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10146_ _10147_/A _10147_/B vssd1 vssd1 vccd1 vccd1 _10146_/Y sky130_fd_sc_hd__nand2b_1
X_10077_ _10077_/A _10077_/B vssd1 vssd1 vccd1 vccd1 _10078_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_69_172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06954__B _06954_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10979_ _10979_/A _10979_/B vssd1 vssd1 vccd1 vccd1 _10981_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__11641__B2 _12254_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12718_ _12718_/A _12718_/B vssd1 vssd1 vccd1 vccd1 _12725_/C sky130_fd_sc_hd__nand2_2
XANTENNA__07131__A _07210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12197__A2 _11343_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12649_ reg1_val[5] _12649_/B vssd1 vssd1 vccd1 vccd1 _12650_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_5_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12691__B _12692_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09860_ _07017_/X _10664_/A _10567_/A fanout30/X vssd1 vssd1 vccd1 vccd1 _09861_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_110_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09791_ _09791_/A _09791_/B vssd1 vssd1 vccd1 vccd1 _09804_/A sky130_fd_sc_hd__xor2_4
X_08811_ _08811_/A _08811_/B _08811_/C vssd1 vssd1 vccd1 vccd1 _08813_/B sky130_fd_sc_hd__nand3_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08742_ _08742_/A _08742_/B vssd1 vssd1 vccd1 vccd1 _08743_/B sky130_fd_sc_hd__xnor2_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09522__B1 _09351_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08673_ _08673_/A _08673_/B vssd1 vssd1 vccd1 vccd1 _08678_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_95_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout174_A _09236_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07624_ _07624_/A _07624_/B _07993_/A vssd1 vssd1 vccd1 vccd1 _07625_/B sky130_fd_sc_hd__and3_1
XFILLER_0_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09825__A1 _11118_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13082__B1 _06892_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07555_ _07555_/A _07555_/B vssd1 vssd1 vccd1 vccd1 _07556_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_48_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10667__A _10959_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07486_ _07487_/A _07487_/B vssd1 vssd1 vccd1 vccd1 _09209_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_8_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09225_ _09415_/B _09225_/B vssd1 vssd1 vccd1 vccd1 _09249_/A sky130_fd_sc_hd__nor2_1
XANTENNA__08137__A _11564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09667__S _09669_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09156_ _09163_/A _09157_/B vssd1 vssd1 vccd1 vccd1 _09156_/Y sky130_fd_sc_hd__nor2_8
XANTENNA__10199__A1 _11294_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10199__B2 _10418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09087_ _09085_/X _09086_/X _09336_/S vssd1 vssd1 vccd1 vccd1 _09087_/X sky130_fd_sc_hd__mux2_1
XANTENNA__08261__B1 _08656_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08107_ _08108_/A _08108_/B vssd1 vssd1 vccd1 vccd1 _08765_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_16_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13137__B2 _12790_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08038_ _08038_/A _08038_/B _08038_/C vssd1 vssd1 vccd1 vccd1 _08041_/B sky130_fd_sc_hd__or3_1
X_10000_ _09854_/B _09958_/B _10748_/A vssd1 vssd1 vccd1 vccd1 _10000_/X sky130_fd_sc_hd__a21o_1
XANTENNA_fanout87_A _07204_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09989_ reg1_val[5] curr_PC[5] vssd1 vssd1 vccd1 vccd1 _09990_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08600__A _09897_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07216__A _10165_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11951_ _11985_/B _11951_/B vssd1 vssd1 vccd1 vccd1 _11951_/Y sky130_fd_sc_hd__nand2b_1
X_10902_ _10891_/X _10892_/Y _11630_/B _09111_/S _10899_/X vssd1 vssd1 vccd1 vccd1
+ _10902_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_98_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11882_ reg1_val[22] curr_PC[22] vssd1 vssd1 vccd1 vccd1 _11883_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_67_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09431__A _09431_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10833_ _10833_/A _10833_/B vssd1 vssd1 vccd1 vccd1 _10835_/C sky130_fd_sc_hd__or2_1
X_10764_ hold203/A _10764_/B vssd1 vssd1 vccd1 vccd1 _10890_/B sky130_fd_sc_hd__or2_1
XFILLER_0_94_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10426__A2 _11472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12503_ _12509_/B _12503_/B vssd1 vssd1 vccd1 vccd1 new_PC[8] sky130_fd_sc_hd__and2_4
XFILLER_0_66_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10695_ _10844_/A _10695_/B _10695_/C vssd1 vssd1 vccd1 vccd1 _10844_/B sky130_fd_sc_hd__and3b_1
X_12434_ hold215/A _12399_/X _12434_/B1 vssd1 vssd1 vccd1 vccd1 _12435_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_81_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07886__A _11385_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12365_ _10928_/A _07508_/B fanout6/X _12316_/B vssd1 vssd1 vccd1 vccd1 _12365_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_22_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11316_ _11316_/A _11316_/B vssd1 vssd1 vccd1 vccd1 _11421_/B sky130_fd_sc_hd__and2_2
XANTENNA__06716__A_N _06981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12296_ _09653_/A _09061_/A _09061_/B _09163_/X vssd1 vssd1 vccd1 vccd1 _12296_/X
+ sky130_fd_sc_hd__a31o_1
X_11247_ _10119_/S _09146_/X _09181_/X vssd1 vssd1 vccd1 vccd1 _11247_/X sky130_fd_sc_hd__o21a_1
XANTENNA__08555__A1 _12804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07358__A2 _10948_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08555__B2 _09768_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11178_ _11176_/Y _11178_/B vssd1 vssd1 vccd1 vccd1 _11181_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__13128__A _13128_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10251__S _11118_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10129_ _09991_/A _09988_/Y _09990_/B vssd1 vssd1 vccd1 vccd1 _10133_/A sky130_fd_sc_hd__o21a_1
XANTENNA__07126__A _09442_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08307__B2 _08436_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08307__A1 _08739_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12967__A _13214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06965__A _06988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12686__B _12686_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07340_ _09594_/A _07340_/B vssd1 vssd1 vccd1 vccd1 _07350_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_18_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09010_ _09010_/A _09010_/B vssd1 vssd1 vccd1 vccd1 _09015_/A sky130_fd_sc_hd__xnor2_1
X_07271_ _07672_/A _07672_/B _07234_/X vssd1 vssd1 vccd1 vccd1 _07309_/B sky130_fd_sc_hd__o21a_2
XFILLER_0_60_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold102 hold102/A vssd1 vssd1 vccd1 vccd1 hold102/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold113 hold128/X vssd1 vssd1 vccd1 vccd1 hold113/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold135 hold135/A vssd1 vssd1 vccd1 vccd1 hold135/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold124 hold124/A vssd1 vssd1 vccd1 vccd1 hold124/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12207__A _12317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold157 hold157/A vssd1 vssd1 vccd1 vccd1 hold157/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 hold168/A vssd1 vssd1 vccd1 vccd1 hold168/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold146 hold146/A vssd1 vssd1 vccd1 vccd1 hold146/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold179 hold179/A vssd1 vssd1 vccd1 vccd1 hold179/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09912_ _09912_/A _09912_/B vssd1 vssd1 vccd1 vccd1 _09913_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_1_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09843_ _09843_/A _09843_/B vssd1 vssd1 vccd1 vccd1 _09843_/Y sky130_fd_sc_hd__xnor2_2
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07036__A _07036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09774_ _09774_/A _09774_/B vssd1 vssd1 vccd1 vccd1 _09775_/B sky130_fd_sc_hd__xnor2_1
X_06986_ _10707_/A _06986_/B vssd1 vssd1 vccd1 vccd1 _06986_/Y sky130_fd_sc_hd__xnor2_2
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08725_ _08726_/A _08726_/B vssd1 vssd1 vccd1 vccd1 _08793_/A sky130_fd_sc_hd__nor2_1
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08656_ _08673_/A _08656_/B vssd1 vssd1 vccd1 vccd1 _08666_/B sky130_fd_sc_hd__or2_1
XFILLER_0_49_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09251__A _09251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08587_ _08609_/A _08609_/B vssd1 vssd1 vccd1 vccd1 _08589_/C sky130_fd_sc_hd__nand2_1
XANTENNA__07521__A2 _12804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07607_ _09768_/A1 _07087_/A _07087_/B fanout66/X _12808_/A vssd1 vssd1 vccd1 vccd1
+ _07608_/B sky130_fd_sc_hd__o32a_1
X_07538_ _07537_/B _07537_/C _11987_/A vssd1 vssd1 vccd1 vccd1 _07540_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_119_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07469_ _07470_/A _07470_/B vssd1 vssd1 vccd1 vccd1 _09205_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_64_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07285__A1 _07149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07285__B2 _12214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09208_ _09208_/A _09208_/B vssd1 vssd1 vccd1 vccd1 _09285_/A sky130_fd_sc_hd__xnor2_4
X_10480_ _10480_/A _10480_/B vssd1 vssd1 vccd1 vccd1 _10483_/A sky130_fd_sc_hd__or2_1
X_09139_ reg1_val[5] reg1_val[26] _09142_/S vssd1 vssd1 vccd1 vccd1 _09139_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_115_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12150_ _12150_/A _12261_/A vssd1 vssd1 vccd1 vccd1 _12151_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_20_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11101_ _10866_/Y _11320_/A _11319_/A vssd1 vssd1 vccd1 vccd1 _11515_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_32_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12081_ _12081_/A _12081_/B _12081_/C vssd1 vssd1 vccd1 vccd1 _12082_/B sky130_fd_sc_hd__or3_1
X_11032_ _10871_/A _10871_/B _10996_/A _10996_/B vssd1 vssd1 vccd1 vccd1 _11033_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09734__B1 _08507_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12983_ _13013_/A hold204/X vssd1 vssd1 vccd1 vccd1 _13294_/D sky130_fd_sc_hd__and2_1
X_11934_ _11934_/A _11934_/B vssd1 vssd1 vccd1 vccd1 _11936_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_115_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11865_ _11698_/A _11781_/A _11783_/B vssd1 vssd1 vccd1 vccd1 _11865_/Y sky130_fd_sc_hd__a21oi_1
X_11796_ _11794_/X _11795_/X _12423_/A vssd1 vssd1 vccd1 vccd1 _11797_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_82_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10816_ _10444_/A _10710_/B _10711_/Y vssd1 vssd1 vccd1 vccd1 _10821_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_125_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10747_ _10660_/X _10782_/B _10746_/Y vssd1 vssd1 vccd1 vccd1 _10747_/X sky130_fd_sc_hd__o21a_1
XANTENNA_clkbuf_4_11_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10678_ _10570_/A _10571_/B _12067_/A _10571_/A vssd1 vssd1 vccd1 vccd1 _10679_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_112_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09100__S _09108_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12417_ _12417_/A _12417_/B vssd1 vssd1 vccd1 vccd1 _12419_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06787__B1 _06785_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12348_ reg1_val[28] reg1_val[29] _12348_/C vssd1 vssd1 vccd1 vccd1 _12429_/C sky130_fd_sc_hd__and3_1
XFILLER_0_50_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12279_ _12414_/B vssd1 vssd1 vccd1 vccd1 _12380_/B sky130_fd_sc_hd__inv_2
X_06840_ reg1_val[27] _07144_/A vssd1 vssd1 vccd1 vccd1 _06840_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__10335__A1 _11146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_58 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10335__B2 _11294_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07751__A2 _07033_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06771_ _06771_/A _06771_/B _12654_/B vssd1 vssd1 vccd1 vccd1 _06771_/X sky130_fd_sc_hd__or3b_1
X_08510_ _08740_/A _08546_/A _08547_/A vssd1 vssd1 vccd1 vccd1 _08519_/B sky130_fd_sc_hd__a21oi_1
X_09490_ _09376_/X _09542_/C _11707_/A vssd1 vssd1 vccd1 vccd1 _09490_/Y sky130_fd_sc_hd__o21ai_1
X_08441_ _09445_/A _08441_/B vssd1 vssd1 vccd1 vccd1 _08442_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_105_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08372_ _08372_/A _08372_/B vssd1 vssd1 vccd1 vccd1 _08428_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_85_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07323_ _07573_/B _07323_/B vssd1 vssd1 vccd1 vccd1 _07325_/B sky130_fd_sc_hd__nor2_1
XANTENNA__12260__A1 fanout12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12260__B2 _12316_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11063__A2 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout137_A _12812_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07254_ reg1_val[28] _07254_/B _07254_/C _12765_/B vssd1 vssd1 vccd1 vccd1 _07503_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_0_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10664__B _12316_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07185_ reg1_val[6] _07185_/B vssd1 vssd1 vccd1 vccd1 _07188_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_14_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06793__A3 _12639_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09826_ _09122_/X _09144_/X _10250_/S vssd1 vssd1 vccd1 vccd1 _10880_/B sky130_fd_sc_hd__mux2_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06969_ _06961_/Y _06966_/Y _11343_/A vssd1 vssd1 vccd1 vccd1 _06969_/Y sky130_fd_sc_hd__a21oi_1
X_09757_ _10165_/A _09757_/B vssd1 vssd1 vccd1 vccd1 _09761_/A sky130_fd_sc_hd__xor2_1
XANTENNA__06950__B1 _07200_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08708_ _08710_/A _08710_/B vssd1 vssd1 vccd1 vccd1 _08708_/X sky130_fd_sc_hd__and2_1
XANTENNA__11826__A1 _12067_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09688_ hold238/A hold248/A hold290/A vssd1 vssd1 vccd1 vccd1 _09688_/X sky130_fd_sc_hd__or3_1
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11826__B2 _12150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08639_ _08622_/B _08626_/Y _08629_/X _08638_/Y vssd1 vssd1 vccd1 vccd1 _08695_/A
+ sky130_fd_sc_hd__a211oi_1
XFILLER_0_49_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11650_ _11034_/B _11650_/B _11650_/C _11650_/D vssd1 vssd1 vccd1 vccd1 _12169_/A
+ sky130_fd_sc_hd__nand4b_4
Xfanout30 _07014_/Y vssd1 vssd1 vccd1 vccd1 fanout30/X sky130_fd_sc_hd__buf_6
XFILLER_0_92_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout63 _07138_/Y vssd1 vssd1 vccd1 vccd1 _12846_/A sky130_fd_sc_hd__clkbuf_8
Xfanout52 _07169_/Y vssd1 vssd1 vccd1 vccd1 _12844_/A sky130_fd_sc_hd__buf_4
XFILLER_0_64_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout41 _12834_/A vssd1 vssd1 vccd1 vccd1 _11751_/A sky130_fd_sc_hd__buf_6
Xfanout74 fanout75/X vssd1 vssd1 vccd1 vccd1 fanout74/X sky130_fd_sc_hd__buf_6
X_11581_ _11582_/A _11582_/B vssd1 vssd1 vccd1 vccd1 _11583_/A sky130_fd_sc_hd__or2_1
X_10601_ _10601_/A _10601_/B vssd1 vssd1 vccd1 vccd1 _10603_/C sky130_fd_sc_hd__xor2_1
X_13320_ _13343_/CLK hold6/X vssd1 vssd1 vccd1 vccd1 hold5/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10532_ _10780_/A _10409_/X _10502_/X _10531_/X vssd1 vssd1 vccd1 vccd1 dest_val[9]
+ sky130_fd_sc_hd__o22a_4
XFILLER_0_52_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout85 _12830_/A vssd1 vssd1 vccd1 vccd1 _09745_/B sky130_fd_sc_hd__buf_4
Xfanout96 _12818_/A vssd1 vssd1 vccd1 vccd1 _10818_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_107_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10574__B _10574_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13251_ _13380_/CLK hold60/X vssd1 vssd1 vccd1 vccd1 hold59/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10463_ _10570_/A fanout48/X _10570_/B _10571_/A vssd1 vssd1 vccd1 vccd1 _10464_/B
+ sky130_fd_sc_hd__o22a_1
X_13182_ hold293/X _12789_/B _13181_/X _12790_/A vssd1 vssd1 vccd1 vccd1 _13183_/B
+ sky130_fd_sc_hd__a22o_1
X_10394_ _09835_/B _10393_/X hold273/A vssd1 vssd1 vccd1 vccd1 _10394_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_103_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12202_ curr_PC[25] _12201_/C curr_PC[26] vssd1 vssd1 vccd1 vccd1 _12202_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_20_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07430__A1 _12842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07430__B2 _12844_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12133_ curr_PC[25] _12201_/C _12455_/S vssd1 vssd1 vccd1 vccd1 _12133_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__10590__A _10710_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12064_ _12065_/A _12065_/B vssd1 vssd1 vccd1 vccd1 _12066_/A sky130_fd_sc_hd__nand2_1
X_11015_ _11633_/B _11127_/B hold212/A vssd1 vssd1 vccd1 vccd1 _11015_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__09183__A1 _09108_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07733__A2 fanout99/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12966_ hold238/A _13213_/B2 _13213_/A2 hold197/X vssd1 vssd1 vccd1 vccd1 hold198/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11817__B2 _09163_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12897_ hold7/X hold273/X vssd1 vssd1 vccd1 vccd1 _12897_/X sky130_fd_sc_hd__and2b_1
XANTENNA__07497__A1 _07149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11917_ _11918_/A _11918_/B vssd1 vssd1 vccd1 vccd1 _12012_/B sky130_fd_sc_hd__nand2_1
XTAP_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11848_ _11847_/A _12214_/B _11847_/C vssd1 vssd1 vccd1 vccd1 _11849_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_28_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12793__A2 _13087_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11779_ _11779_/A _11779_/B vssd1 vssd1 vccd1 vccd1 _11782_/C sky130_fd_sc_hd__xor2_1
XFILLER_0_27_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07421__B2 _07149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07421__A1 _08436_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08990_ _09960_/B _09961_/A vssd1 vssd1 vccd1 vccd1 _10105_/B sky130_fd_sc_hd__and2_1
XFILLER_0_11_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09174__A1 _09669_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10308__A1 _10664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10308__B2 _10818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07941_ _08072_/A _08072_/B _07930_/X vssd1 vssd1 vccd1 vccd1 _07964_/B sky130_fd_sc_hd__a21oi_2
X_07872_ _07876_/A _07876_/B vssd1 vssd1 vccd1 vccd1 _07872_/X sky130_fd_sc_hd__or2_1
X_06823_ _11224_/A _06822_/X _06710_/X vssd1 vssd1 vccd1 vccd1 _06823_/X sky130_fd_sc_hd__o21ba_1
X_09611_ _09746_/A _09611_/B _09611_/C vssd1 vssd1 vccd1 vccd1 _09618_/A sky130_fd_sc_hd__and3_1
X_06754_ reg1_val[8] _07089_/A vssd1 vssd1 vccd1 vccd1 _06754_/Y sky130_fd_sc_hd__nor2_1
X_09542_ _09542_/A _09542_/B _09542_/C vssd1 vssd1 vccd1 vccd1 _10275_/A sky130_fd_sc_hd__and3_1
X_06685_ instruction[28] _06694_/B vssd1 vssd1 vccd1 vccd1 _12639_/B sky130_fd_sc_hd__and2_4
XFILLER_0_93_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09473_ _09473_/A _09473_/B vssd1 vssd1 vccd1 vccd1 _09474_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_66_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07488__B2 _12830_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07488__A1 _12828_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08424_ _08424_/A _08424_/B vssd1 vssd1 vccd1 vccd1 _08426_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__07033__B _07033_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08437__B1 _08730_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08355_ _10949_/A _08414_/A vssd1 vssd1 vccd1 vccd1 _08368_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_18_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07306_ _07308_/A _07306_/B vssd1 vssd1 vccd1 vccd1 _07674_/B sky130_fd_sc_hd__nor2_2
XANTENNA__11587__A3 _11557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08286_ _08288_/B _08288_/A vssd1 vssd1 vccd1 vccd1 _08290_/A sky130_fd_sc_hd__nand2b_1
X_07237_ _12848_/A _08436_/B _10941_/B _07149_/A vssd1 vssd1 vccd1 vccd1 _07238_/B
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_61_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07168_ _07140_/C _07142_/B _07142_/C _07223_/B vssd1 vssd1 vccd1 vccd1 _07169_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_112_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07099_ _07099_/A _07099_/B vssd1 vssd1 vccd1 vccd1 _07099_/X sky130_fd_sc_hd__and2_1
Xfanout220 _13213_/A2 vssd1 vssd1 vccd1 vccd1 _13016_/B1 sky130_fd_sc_hd__buf_2
XFILLER_0_100_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout231 _09669_/S vssd1 vssd1 vccd1 vccd1 _09663_/S sky130_fd_sc_hd__clkbuf_8
Xfanout264 _12455_/S vssd1 vssd1 vccd1 vccd1 _12622_/S sky130_fd_sc_hd__clkbuf_8
Xfanout253 _09159_/X vssd1 vssd1 vccd1 vccd1 _09527_/B sky130_fd_sc_hd__buf_4
Xfanout242 _06779_/X vssd1 vssd1 vccd1 vccd1 _09147_/S sky130_fd_sc_hd__buf_2
Xfanout297 _13242_/A vssd1 vssd1 vccd1 vccd1 _13128_/A sky130_fd_sc_hd__buf_4
Xfanout275 _13213_/B2 vssd1 vssd1 vccd1 vccd1 _13004_/A2 sky130_fd_sc_hd__buf_4
X_09809_ _09810_/A _09810_/B _10368_/A vssd1 vssd1 vccd1 vccd1 _09811_/A sky130_fd_sc_hd__a21o_1
Xfanout286 _06587_/X vssd1 vssd1 vccd1 vccd1 _12782_/A sky130_fd_sc_hd__buf_8
X_12820_ _12820_/A _12830_/B vssd1 vssd1 vccd1 vccd1 _12820_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_69_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07479__B2 _12842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07479__A1 _12840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12751_ reg1_val[25] _12782_/A vssd1 vssd1 vccd1 vccd1 _12754_/B sky130_fd_sc_hd__xnor2_4
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12682_ _12683_/A _12683_/B _12683_/C vssd1 vssd1 vccd1 vccd1 _12689_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_37_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11702_ _11702_/A _11868_/A vssd1 vssd1 vccd1 vccd1 _11702_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_127_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11633_ hold177/A _11633_/B _11720_/B vssd1 vssd1 vccd1 vccd1 _11633_/X sky130_fd_sc_hd__and3_1
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11564_ _11564_/A _11564_/B vssd1 vssd1 vccd1 vccd1 _11568_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__10786__A1 _07087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10786__B2 fanout66/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13303_ _13307_/CLK _13303_/D vssd1 vssd1 vccd1 vccd1 hold210/A sky130_fd_sc_hd__dfxtp_1
X_10515_ _10111_/X _10514_/X _11233_/S vssd1 vssd1 vccd1 vccd1 _10516_/A sky130_fd_sc_hd__mux2_1
X_11495_ _11495_/A _11495_/B vssd1 vssd1 vccd1 vccd1 _11497_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_122_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13234_ hold298/X _12790_/A _13233_/Y _12789_/B hold109/X vssd1 vssd1 vccd1 vccd1
+ hold110/A sky130_fd_sc_hd__a32o_1
XFILLER_0_33_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10446_ _07154_/A _07154_/B _10706_/B2 vssd1 vssd1 vccd1 vccd1 _10448_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_60_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13165_ _13165_/A _13165_/B vssd1 vssd1 vccd1 vccd1 _13165_/Y sky130_fd_sc_hd__xnor2_1
X_10377_ _06815_/X _10376_/X _12388_/S vssd1 vssd1 vccd1 vccd1 _10378_/B sky130_fd_sc_hd__mux2_1
XANTENNA__07954__A2 _07099_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13096_ _12913_/X _13096_/B vssd1 vssd1 vccd1 vccd1 _13097_/B sky130_fd_sc_hd__nand2b_1
X_12116_ _12113_/Y _12115_/X _12112_/Y vssd1 vssd1 vccd1 vccd1 _12116_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__07260__B1_N _10928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12047_ _11636_/B _12119_/B hold254/A vssd1 vssd1 vccd1 vccd1 _12047_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__09614__A _09614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06957__B _07064_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12949_ _13206_/B _13207_/A _12869_/X vssd1 vssd1 vccd1 vccd1 _13211_/B sky130_fd_sc_hd__a21o_1
XANTENNA__07134__A _07223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06973__A _07130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12186__S _12429_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08140_ _08140_/A _08140_/B vssd1 vssd1 vccd1 vccd1 _08150_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__10777__A1 _11876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08071_ _07916_/A _07916_/B _07916_/C vssd1 vssd1 vccd1 vccd1 _08073_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_113_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07022_ reg1_val[23] _07022_/B vssd1 vssd1 vccd1 vccd1 _07524_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_3_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09919__B1 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11726__B1 _12247_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13191__A2 _13213_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10529__A1 _12254_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09395__A1 _07099_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08973_ _08971_/A _08971_/B _08963_/X vssd1 vssd1 vccd1 vccd1 _09487_/C sky130_fd_sc_hd__a21boi_1
Xhold17 hold17/A vssd1 vssd1 vccd1 vccd1 hold17/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold28 hold28/A vssd1 vssd1 vccd1 vccd1 hold28/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07924_ _12820_/A _08744_/A2 _08564_/B _08741_/B2 vssd1 vssd1 vccd1 vccd1 _07925_/B
+ sky130_fd_sc_hd__o22a_1
Xhold39 hold39/A vssd1 vssd1 vccd1 vccd1 hold39/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09698__A2 _09672_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07855_ _07854_/B _07854_/C _07850_/X vssd1 vssd1 vccd1 vccd1 _07905_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_127_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06806_ reg2_val[0] _06720_/B _06702_/A _06805_/X vssd1 vssd1 vccd1 vccd1 _06806_/Y
+ sky130_fd_sc_hd__a22oi_1
X_07786_ _08733_/A _07786_/B vssd1 vssd1 vccd1 vccd1 _07790_/A sky130_fd_sc_hd__xnor2_2
X_06737_ _10767_/S _06737_/B vssd1 vssd1 vccd1 vccd1 _10752_/A sky130_fd_sc_hd__nor2_1
X_09525_ _09527_/A _09525_/B vssd1 vssd1 vccd1 vccd1 _09525_/Y sky130_fd_sc_hd__nor2_1
X_06668_ reg1_val[20] _07220_/A vssd1 vssd1 vccd1 vccd1 _06669_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_78_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09456_ _09456_/A _09456_/B vssd1 vssd1 vccd1 vccd1 _09459_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__08122__A2 _08656_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07330__B1 _12840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08407_ _08419_/B _08419_/A vssd1 vssd1 vccd1 vccd1 _08421_/A sky130_fd_sc_hd__and2b_1
XANTENNA__12206__A1 fanout16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06599_ reg1_val[31] _07064_/B vssd1 vssd1 vccd1 vccd1 _08980_/B sky130_fd_sc_hd__xor2_4
X_09387_ fanout30/X _12808_/A _07089_/Y _07688_/B vssd1 vssd1 vccd1 vccd1 _09388_/B
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_47_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12206__B2 _07282_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10768__A1 _12307_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08338_ _08381_/B _08381_/A vssd1 vssd1 vccd1 vccd1 _08342_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_19_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08269_ _08329_/A _08329_/B _08265_/X vssd1 vssd1 vccd1 vccd1 _08280_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_22_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06987__A3 _07074_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11280_ _11281_/B _11280_/B vssd1 vssd1 vccd1 vccd1 _11402_/A sky130_fd_sc_hd__and2b_1
X_10300_ _10159_/A _10158_/Y _10154_/Y vssd1 vssd1 vccd1 vccd1 _10302_/B sky130_fd_sc_hd__o21a_1
XANTENNA__08603__A _09433_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10231_ _10231_/A _10231_/B vssd1 vssd1 vccd1 vccd1 _10741_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_14_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13182__A2 _12789_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12390__B1 _09156_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06739__A3 _12680_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10162_ _07154_/A _07154_/B _08507_/B vssd1 vssd1 vccd1 vccd1 _10164_/C sky130_fd_sc_hd__a21o_1
XANTENNA__07936__A2 _11558_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10093_ _10093_/A _10093_/B vssd1 vssd1 vccd1 vccd1 _10096_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__08041__C _08041_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08361__A2 _08727_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12803_ hold49/X _12818_/B _12802_/Y _13113_/A vssd1 vssd1 vccd1 vccd1 hold50/A sky130_fd_sc_hd__o211a_1
XFILLER_0_84_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10995_ _11100_/B _11424_/A _10995_/C vssd1 vssd1 vccd1 vccd1 _10996_/B sky130_fd_sc_hd__nand3_1
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12734_ _12746_/B _12734_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[21] sky130_fd_sc_hd__xor2_4
XFILLER_0_123_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12665_ _12663_/Y _12665_/B vssd1 vssd1 vccd1 vccd1 _12666_/B sky130_fd_sc_hd__nand2b_2
XFILLER_0_37_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12596_ _12596_/A vssd1 vssd1 vccd1 vccd1 _12605_/C sky130_fd_sc_hd__inv_2
XFILLER_0_65_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11616_ _11874_/A _11616_/B _11616_/C vssd1 vssd1 vccd1 vccd1 _11618_/A sky130_fd_sc_hd__and3_1
X_11547_ _11545_/Y _11546_/X _11539_/X _11543_/X vssd1 vssd1 vccd1 vccd1 _11547_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_114_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09609__A _11294_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11478_ _11478_/A _11478_/B vssd1 vssd1 vccd1 vccd1 _11479_/B sky130_fd_sc_hd__or2_1
XFILLER_0_0_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13217_ hold281/A _13216_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13217_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_0_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10429_ _10430_/A _10430_/B vssd1 vssd1 vccd1 vccd1 _10429_/X sky130_fd_sc_hd__and2_1
X_13148_ _13245_/A _13148_/B vssd1 vssd1 vccd1 vccd1 _13359_/D sky130_fd_sc_hd__and2_1
XANTENNA__07129__A _07130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13079_ _07522_/A _13087_/B2 hold114/X vssd1 vssd1 vccd1 vccd1 hold115/A sky130_fd_sc_hd__o21a_1
XANTENNA__12133__B1 _12455_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08352__A2 _08744_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07640_ _12804_/A _09614_/A _12802_/A _09613_/A vssd1 vssd1 vccd1 vccd1 _07641_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_88_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07571_ _07571_/A _07571_/B vssd1 vssd1 vccd1 vccd1 _07573_/C sky130_fd_sc_hd__xor2_1
XFILLER_0_87_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09310_ _09190_/X _09542_/B _09309_/Y vssd1 vssd1 vccd1 vccd1 _09371_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__07799__A _08304_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10447__B1 _10448_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07312__B1 _12802_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09241_ _09441_/A _09241_/B _09241_/C vssd1 vssd1 vccd1 vccd1 _09242_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_75_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07863__A1 _08741_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07863__B2 _08732_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09172_ reg1_val[31] _09172_/B vssd1 vssd1 vccd1 vccd1 _09181_/B sky130_fd_sc_hd__and2_2
XFILLER_0_90_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07615__A1 _11294_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08123_ _08733_/A _08123_/B vssd1 vssd1 vccd1 vccd1 _08130_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_126_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07615__B2 _10418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08054_ _08740_/A _08054_/B vssd1 vssd1 vccd1 vccd1 _08055_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_114_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09368__A1 _11118_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07005_ _09669_/S _07006_/B vssd1 vssd1 vccd1 vccd1 _09251_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__07091__A2 _11653_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09238__B _09238_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07039__A _11987_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07918__A2 _08741_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09254__A _12412_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08956_ _08951_/A _08951_/B _08949_/X vssd1 vssd1 vccd1 vccd1 _08965_/A sky130_fd_sc_hd__a21oi_2
X_07907_ _07908_/A _07908_/B vssd1 vssd1 vccd1 vccd1 _07981_/A sky130_fd_sc_hd__nand2b_1
X_08887_ _09043_/B _08840_/Y _09042_/B _09049_/A vssd1 vssd1 vccd1 vccd1 _08887_/X
+ sky130_fd_sc_hd__and4bb_1
X_07838_ _07838_/A _07838_/B vssd1 vssd1 vccd1 vccd1 _07840_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__10686__B1 _10930_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10150__A2 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09508_ _09136_/X _09140_/X _09663_/S vssd1 vssd1 vccd1 vccd1 _09508_/X sky130_fd_sc_hd__mux2_1
X_07769_ _07769_/A _07769_/B vssd1 vssd1 vccd1 vccd1 _07770_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout32_A _12412_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10780_ _10780_/A _10906_/B vssd1 vssd1 vccd1 vccd1 _10780_/Y sky130_fd_sc_hd__nor2_1
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09439_ _09439_/A _09439_/B vssd1 vssd1 vccd1 vccd1 _09460_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_54_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12450_ _12629_/B _12450_/B vssd1 vssd1 vccd1 vccd1 _12451_/B sky130_fd_sc_hd__or2_1
XANTENNA__07221__B _08038_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11401_ _11275_/A _11275_/B _11267_/A vssd1 vssd1 vccd1 vccd1 _11404_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_105_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12381_ _11870_/B _12380_/Y _12379_/X vssd1 vssd1 vccd1 vccd1 _12382_/B sky130_fd_sc_hd__o21ba_1
XFILLER_0_105_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11332_ _11332_/A _11332_/B vssd1 vssd1 vccd1 vccd1 _11332_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_62_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09359__B2 _12394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11263_ _11263_/A _11263_/B vssd1 vssd1 vccd1 vccd1 _11264_/B sky130_fd_sc_hd__and2_1
X_13002_ hold210/X _13004_/A2 _13006_/B1 hold236/X vssd1 vssd1 vccd1 vccd1 hold237/A
+ sky130_fd_sc_hd__a22o_1
X_10214_ _10214_/A _10214_/B vssd1 vssd1 vccd1 vccd1 _10227_/A sky130_fd_sc_hd__xnor2_4
X_11194_ _11070_/A _11070_/B _11068_/X vssd1 vssd1 vccd1 vccd1 _11196_/C sky130_fd_sc_hd__a21o_1
X_10145_ _10959_/A _10145_/B vssd1 vssd1 vccd1 vccd1 _10147_/B sky130_fd_sc_hd__xnor2_1
X_10076_ _10076_/A _10076_/B _10076_/C vssd1 vssd1 vccd1 vccd1 _10077_/B sky130_fd_sc_hd__nor3_2
XFILLER_0_89_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07542__B1 fanout66/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10978_ _10846_/A _10845_/B _10843_/X vssd1 vssd1 vccd1 vccd1 _10979_/B sky130_fd_sc_hd__a21oi_1
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09103__S _09108_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12717_ reg1_val[18] _12741_/B vssd1 vssd1 vccd1 vccd1 _12718_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_128_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07131__B _07131_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12648_ reg1_val[5] _12649_/B vssd1 vssd1 vccd1 vccd1 _12648_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_26_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12579_ _12611_/A _12579_/B vssd1 vssd1 vccd1 vccd1 _12580_/B sky130_fd_sc_hd__or2_1
XFILLER_0_80_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10492__B _10493_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10904__A1 _09156_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08810_ _08046_/A _08046_/C _08046_/B vssd1 vssd1 vccd1 vccd1 _08811_/C sky130_fd_sc_hd__a21o_1
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09790_ _09788_/Y _09790_/B vssd1 vssd1 vccd1 vccd1 _09791_/B sky130_fd_sc_hd__and2b_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08741_ _12820_/A _08741_/A2 _08617_/B _08741_/B2 vssd1 vssd1 vccd1 vccd1 _08742_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09522__A1 _09343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09522__B2 _12626_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08672_ _08681_/A _08672_/B vssd1 vssd1 vccd1 vccd1 _08678_/A sky130_fd_sc_hd__xnor2_1
X_07623_ _07621_/A _07621_/B _07984_/A vssd1 vssd1 vccd1 vccd1 _07626_/B sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout167_A _08584_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07554_ _07555_/B _07555_/A vssd1 vssd1 vccd1 vccd1 _07554_/X sky130_fd_sc_hd__and2b_1
X_07485_ _07485_/A _07485_/B vssd1 vssd1 vccd1 vccd1 _07487_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_36_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09224_ _09223_/B _09224_/B vssd1 vssd1 vccd1 vccd1 _09225_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_8_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09155_ _09170_/B _09159_/B vssd1 vssd1 vccd1 vccd1 _09155_/X sky130_fd_sc_hd__or2_1
XANTENNA__10199__A2 _10574_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09086_ _12626_/A reg1_val[31] _09108_/S vssd1 vssd1 vccd1 vccd1 _09086_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_71_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08261__A1 _08436_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08261__B2 fanout99/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08106_ _08106_/A _08106_/B vssd1 vssd1 vccd1 vccd1 _08108_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_4_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13137__A2 _12789_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08037_ _08733_/A _08037_/B vssd1 vssd1 vccd1 vccd1 _08042_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_31_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09988_ reg1_val[5] curr_PC[5] vssd1 vssd1 vccd1 vccd1 _09988_/Y sky130_fd_sc_hd__nor2_1
X_08939_ _08939_/A _08939_/B vssd1 vssd1 vccd1 vccd1 _09065_/B sky130_fd_sc_hd__xnor2_4
X_11950_ _11951_/B _11985_/B vssd1 vssd1 vccd1 vccd1 _11950_/Y sky130_fd_sc_hd__nand2b_1
X_10901_ _11630_/B vssd1 vssd1 vccd1 vccd1 _10901_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_98_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11881_ reg1_val[22] curr_PC[22] vssd1 vssd1 vccd1 vccd1 _11883_/A sky130_fd_sc_hd__or2_1
XANTENNA__13073__A1 _11987_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10832_ _10961_/A _10961_/B vssd1 vssd1 vccd1 vccd1 _10833_/B sky130_fd_sc_hd__and2_1
X_10763_ _12244_/S _10762_/X _10759_/X vssd1 vssd1 vccd1 vccd1 _10763_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_13_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10259__A1_N _07080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12502_ _12502_/A _12502_/B _12502_/C vssd1 vssd1 vccd1 vccd1 _12503_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_125_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10694_ _10835_/B _10694_/B vssd1 vssd1 vccd1 vccd1 _10695_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_120_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12433_ hold109/A _12431_/X _12432_/Y vssd1 vssd1 vccd1 vccd1 _12433_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_35_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07886__B _07886_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09159__A _09168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12364_ _12317_/A _12317_/B _12320_/A vssd1 vssd1 vccd1 vccd1 _12372_/A sky130_fd_sc_hd__a21o_1
XANTENNA__08063__A _08722_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11315_ _11315_/A _11315_/B _11315_/C vssd1 vssd1 vccd1 vccd1 _11316_/B sky130_fd_sc_hd__nand3_1
X_12295_ _09653_/A _09061_/A _09061_/B vssd1 vssd1 vccd1 vccd1 _12295_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_31_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11246_ _06988_/A _12404_/A _11243_/Y _11245_/Y vssd1 vssd1 vccd1 vccd1 _11249_/B
+ sky130_fd_sc_hd__a211o_1
XANTENNA__09201__B1 _12808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08555__A2 _08661_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11177_ _11177_/A _11177_/B _11177_/C vssd1 vssd1 vccd1 vccd1 _11178_/B sky130_fd_sc_hd__nand3_1
X_10128_ _06767_/X _09154_/Y _09158_/Y _10109_/A _10127_/X vssd1 vssd1 vccd1 vccd1
+ _10128_/X sky130_fd_sc_hd__a221o_1
XANTENNA__07407__A _07485_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07763__B1 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08307__A2 _08732_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10059_ _10059_/A _10059_/B vssd1 vssd1 vccd1 vccd1 _10061_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__06965__B _06981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07142__A _07144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07270_ _07270_/A _07270_/B vssd1 vssd1 vccd1 vccd1 _07672_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_58_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06981__A _06981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09440__B1 _09440_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold103 hold103/A vssd1 vssd1 vccd1 vccd1 hold103/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_51 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold114 hold114/A vssd1 vssd1 vccd1 vccd1 hold114/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold125 hold125/A vssd1 vssd1 vccd1 vccd1 hold125/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold158 hold158/A vssd1 vssd1 vccd1 vccd1 hold158/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold136 hold136/A vssd1 vssd1 vccd1 vccd1 hold136/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold147 hold147/A vssd1 vssd1 vccd1 vccd1 hold147/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09911_ _09911_/A _09911_/B vssd1 vssd1 vccd1 vccd1 _09912_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_1_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold169 hold169/A vssd1 vssd1 vccd1 vccd1 hold169/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_95_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09842_ _09840_/Y _09842_/B vssd1 vssd1 vccd1 vccd1 _09843_/B sky130_fd_sc_hd__nand2b_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07155__A2_N _12852_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09773_ _09774_/A _09774_/B vssd1 vssd1 vccd1 vccd1 _09773_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__07754__B1 _11908_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout284_A _06587_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06985_ _06985_/A _06985_/B vssd1 vssd1 vccd1 vccd1 _06985_/X sky130_fd_sc_hd__and2_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08724_ _08724_/A _08724_/B vssd1 vssd1 vccd1 vccd1 _08726_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__09532__A _12423_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08655_ _08655_/A _08655_/B vssd1 vssd1 vccd1 vccd1 _08666_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_68_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13055__A1 _11164_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09251__B _12264_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08586_ _08586_/A _08586_/B vssd1 vssd1 vccd1 vccd1 _08609_/B sky130_fd_sc_hd__xor2_1
X_07606_ _11470_/A _07606_/B vssd1 vssd1 vccd1 vccd1 _07610_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_88_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07537_ _11987_/A _07537_/B _07537_/C vssd1 vssd1 vccd1 vccd1 _07540_/C sky130_fd_sc_hd__and3_1
XANTENNA__07052__A _11987_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11066__B1 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06891__A _12788_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07468_ _07569_/A _07468_/B vssd1 vssd1 vccd1 vccd1 _07470_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_64_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07285__A2 fanout59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09207_ _09208_/B _09208_/A vssd1 vssd1 vccd1 vccd1 _09469_/B sky130_fd_sc_hd__and2b_1
X_07399_ _07399_/A _07399_/B vssd1 vssd1 vccd1 vccd1 _08958_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_106_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09138_ reg1_val[4] reg1_val[27] _09142_/S vssd1 vssd1 vccd1 vccd1 _09138_/X sky130_fd_sc_hd__mux2_1
X_09069_ _09485_/B _09069_/B vssd1 vssd1 vccd1 vccd1 _12392_/A sky130_fd_sc_hd__xnor2_2
X_11100_ _11100_/A _11100_/B vssd1 vssd1 vccd1 vccd1 _11320_/A sky130_fd_sc_hd__or2_1
X_12080_ _12081_/A _12081_/B _12081_/C vssd1 vssd1 vccd1 vccd1 _12156_/A sky130_fd_sc_hd__o21ai_1
X_11031_ _12448_/S _11028_/X _11029_/X _11030_/Y vssd1 vssd1 vccd1 vccd1 dest_val[13]
+ sky130_fd_sc_hd__a22o_4
XANTENNA__09734__A1 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09734__B2 _12214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12982_ hold203/X _13004_/A2 _13006_/B1 hold189/X vssd1 vssd1 vccd1 vccd1 hold204/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_86_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09442__A _09442_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11933_ _11934_/A _11934_/B vssd1 vssd1 vccd1 vccd1 _11933_/X sky130_fd_sc_hd__and2b_1
XANTENNA__06785__B _06799_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11864_ _12165_/A vssd1 vssd1 vccd1 vccd1 _12098_/B sky130_fd_sc_hd__inv_2
XANTENNA__08170__B1 _08216_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10815_ _10971_/A _10804_/Y _10814_/C vssd1 vssd1 vccd1 vccd1 _10822_/B sky130_fd_sc_hd__o21ba_1
XANTENNA__11057__B1 _12067_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11795_ _06676_/C _06827_/Y _06831_/B vssd1 vssd1 vccd1 vccd1 _11795_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_67_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10746_ _10660_/X _10782_/B _12290_/A vssd1 vssd1 vccd1 vccd1 _10746_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_55_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07897__A _11564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10677_ _10677_/A _10677_/B vssd1 vssd1 vccd1 vccd1 _10680_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_125_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12416_ _12333_/Y _12414_/C _12414_/X _12230_/B _12415_/Y vssd1 vssd1 vccd1 vccd1
+ _12417_/B sky130_fd_sc_hd__o221a_1
XFILLER_0_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12347_ _12426_/A _09077_/A _09077_/B _12428_/A _12346_/Y vssd1 vssd1 vccd1 vccd1
+ _12362_/B sky130_fd_sc_hd__o311a_1
XFILLER_0_50_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12278_ _12276_/X _12278_/B vssd1 vssd1 vccd1 vccd1 _12414_/B sky130_fd_sc_hd__nand2b_1
X_11229_ _11117_/A _11117_/B _11115_/B vssd1 vssd1 vccd1 vccd1 _11230_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_4_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07736__B1 _12820_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10335__A2 fanout23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06770_ _06575_/Y _06589_/X _06592_/Y _12654_/B _06596_/A vssd1 vssd1 vccd1 vccd1
+ _06770_/X sky130_fd_sc_hd__o2111a_2
XANTENNA__12697__B _12698_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06695__B _12634_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08440_ _08721_/B1 _08661_/A2 _08727_/B1 _08739_/A1 vssd1 vssd1 vccd1 vccd1 _08441_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_86_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08371_ _08371_/A _08371_/B vssd1 vssd1 vccd1 vccd1 _08372_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_128_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09498__S _09666_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07322_ _07322_/A _07322_/B vssd1 vssd1 vccd1 vccd1 _07323_/B sky130_fd_sc_hd__and2_1
XFILLER_0_45_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12260__A2 fanout9/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07253_ reg1_val[24] reg1_val[25] reg1_val[26] reg1_val[27] vssd1 vssd1 vccd1 vccd1
+ _12765_/B sky130_fd_sc_hd__or4_2
XFILLER_0_116_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07184_ reg1_val[4] reg1_val[5] _07160_/B _07200_/A vssd1 vssd1 vccd1 vccd1 _07185_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_6_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08431__A _08740_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09825_ _11118_/A _09823_/X _09824_/X _11233_/S vssd1 vssd1 vccd1 vccd1 _09825_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07047__A _11180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06968_ _06961_/Y _06966_/Y _07223_/B vssd1 vssd1 vccd1 vccd1 _06968_/X sky130_fd_sc_hd__a21o_1
X_09756_ _09568_/A _09567_/B _09568_/B fanout13/X vssd1 vssd1 vccd1 vccd1 _09757_/B
+ sky130_fd_sc_hd__o22a_1
X_09687_ _09686_/B _09687_/B vssd1 vssd1 vccd1 vccd1 _09687_/Y sky130_fd_sc_hd__nand2b_1
X_08707_ _08707_/A _08707_/B vssd1 vssd1 vccd1 vccd1 _09017_/B sky130_fd_sc_hd__nand2_1
XANTENNA__11826__A2 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06899_ instruction[12] _06902_/B vssd1 vssd1 vccd1 vccd1 dest_idx[1] sky130_fd_sc_hd__and2_4
XFILLER_0_96_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08638_ _08652_/A _08652_/B vssd1 vssd1 vccd1 vccd1 _08638_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_96_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08569_ _08572_/A _08572_/B vssd1 vssd1 vccd1 vccd1 _08571_/B sky130_fd_sc_hd__nor2_1
Xfanout20 _09609_/B vssd1 vssd1 vccd1 vccd1 _10570_/A sky130_fd_sc_hd__buf_6
XFILLER_0_37_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout31 _12412_/B vssd1 vssd1 vccd1 vccd1 _12214_/B sky130_fd_sc_hd__buf_4
XFILLER_0_107_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout42 _12834_/A vssd1 vssd1 vccd1 vccd1 _10575_/B sky130_fd_sc_hd__buf_4
Xfanout64 _09396_/B vssd1 vssd1 vccd1 vccd1 _10571_/A sky130_fd_sc_hd__clkbuf_8
Xfanout53 _12842_/A vssd1 vssd1 vccd1 vccd1 _11989_/A sky130_fd_sc_hd__clkbuf_8
X_10600_ _10455_/A _10455_/C _10455_/B vssd1 vssd1 vccd1 vccd1 _10601_/B sky130_fd_sc_hd__a21bo_1
X_11580_ _11580_/A _11580_/B vssd1 vssd1 vccd1 vccd1 _11582_/B sky130_fd_sc_hd__or2_1
XFILLER_0_92_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout86 _07207_/X vssd1 vssd1 vccd1 vccd1 _12830_/A sky130_fd_sc_hd__buf_4
X_10531_ _11876_/A _10503_/X _10504_/Y _10530_/Y vssd1 vssd1 vccd1 vccd1 _10531_/X
+ sky130_fd_sc_hd__a31o_1
Xfanout97 _07075_/Y vssd1 vssd1 vccd1 vccd1 _12818_/A sky130_fd_sc_hd__buf_8
XANTENNA_fanout9_A fanout9/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout75 _06985_/X vssd1 vssd1 vccd1 vccd1 fanout75/X sky130_fd_sc_hd__buf_8
XFILLER_0_9_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13250_ _13355_/CLK _13250_/D vssd1 vssd1 vccd1 vccd1 hold61/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12201_ curr_PC[25] curr_PC[26] _12201_/C vssd1 vssd1 vccd1 vccd1 _12204_/B sky130_fd_sc_hd__and3_1
X_10462_ _11163_/A _10462_/B vssd1 vssd1 vccd1 vccd1 _10465_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13181_ hold263/X _13180_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13181_/X sky130_fd_sc_hd__mux2_1
X_10393_ hold294/A _10522_/C vssd1 vssd1 vccd1 vccd1 _10393_/X sky130_fd_sc_hd__or2_1
XFILLER_0_60_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07430__A2 _09567_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09437__A _10449_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12132_ _12103_/Y _12104_/X _12107_/X _12131_/X vssd1 vssd1 vccd1 vccd1 _12132_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_32_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12063_ _12261_/A _12063_/B vssd1 vssd1 vccd1 vccd1 _12065_/B sky130_fd_sc_hd__xnor2_1
X_11014_ _13295_/Q _11014_/B vssd1 vssd1 vccd1 vccd1 _11127_/B sky130_fd_sc_hd__or2_1
XANTENNA__12798__A _12798_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12965_ _13214_/A hold239/X vssd1 vssd1 vccd1 vccd1 _13285_/D sky130_fd_sc_hd__and2_1
XANTENNA__11278__B1 _11923_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08143__B1 _08727_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11916_ _12012_/A _11916_/B vssd1 vssd1 vccd1 vccd1 _11918_/B sky130_fd_sc_hd__and2_1
X_12896_ hold288/A hold33/X vssd1 vssd1 vccd1 vccd1 _13134_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__07497__A2 _12412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11847_ _11847_/A _12214_/B _11847_/C vssd1 vssd1 vccd1 vccd1 _11931_/B sky130_fd_sc_hd__or3_1
XTAP_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11778_ _11779_/B _11779_/A vssd1 vssd1 vccd1 vccd1 _11861_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09111__S _09111_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10729_ _10729_/A _10729_/B vssd1 vssd1 vccd1 vccd1 _10731_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_27_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13379_ _13380_/CLK hold66/X vssd1 vssd1 vccd1 vccd1 hold63/A sky130_fd_sc_hd__dfxtp_1
Xclkbuf_4_7_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13314_/CLK sky130_fd_sc_hd__clkbuf_8
XANTENNA__07421__A2 _12854_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07957__B1 _11564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07940_ _07940_/A _07940_/B vssd1 vssd1 vccd1 vccd1 _08072_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_76_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07709__B1 _08752_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10308__A2 fanout16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07871_ _08731_/A _07871_/B vssd1 vssd1 vccd1 vccd1 _07876_/B sky130_fd_sc_hd__xnor2_1
X_06822_ _11111_/A _06821_/X _06716_/Y vssd1 vssd1 vccd1 vccd1 _06822_/X sky130_fd_sc_hd__o21a_1
X_09610_ _10418_/A _09745_/A vssd1 vssd1 vccd1 vccd1 _09611_/C sky130_fd_sc_hd__or2_1
X_06753_ _07089_/A reg1_val[8] vssd1 vssd1 vccd1 vccd1 _06753_/X sky130_fd_sc_hd__and2b_1
X_09541_ _10780_/A _09701_/B _09540_/Y _09538_/X vssd1 vssd1 vccd1 vccd1 dest_val[2]
+ sky130_fd_sc_hd__o31ai_4
XFILLER_0_116_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06684_ _06866_/A vssd1 vssd1 vccd1 vccd1 _11623_/A sky130_fd_sc_hd__inv_2
X_09472_ _09473_/A _09473_/B vssd1 vssd1 vccd1 vccd1 _09472_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__07488__A2 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08423_ _08454_/A _08454_/B _08386_/Y vssd1 vssd1 vccd1 vccd1 _08426_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_74_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08354_ _08413_/A _08413_/B vssd1 vssd1 vccd1 vccd1 _08414_/A sky130_fd_sc_hd__nor2_1
X_07305_ _07633_/A _07294_/C _07294_/A vssd1 vssd1 vccd1 vccd1 _07306_/B sky130_fd_sc_hd__a21oi_1
X_08285_ _08285_/A _08285_/B vssd1 vssd1 vccd1 vccd1 _08288_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_116_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07236_ _09441_/A _07236_/B vssd1 vssd1 vccd1 vccd1 _07241_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_33_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07167_ _07167_/A _09758_/A vssd1 vssd1 vccd1 vccd1 _07167_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__10691__A _11172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07098_ _11470_/A _11470_/B _09746_/A vssd1 vssd1 vccd1 vccd1 _07099_/B sky130_fd_sc_hd__or3b_4
Xfanout221 _06890_/Y vssd1 vssd1 vccd1 vccd1 _13213_/A2 sky130_fd_sc_hd__buf_4
XFILLER_0_100_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout232 _06800_/Y vssd1 vssd1 vccd1 vccd1 _09669_/S sky130_fd_sc_hd__clkbuf_8
Xfanout210 _09441_/A vssd1 vssd1 vccd1 vccd1 _08733_/A sky130_fd_sc_hd__buf_12
Xfanout265 _12455_/S vssd1 vssd1 vccd1 vccd1 _12586_/S sky130_fd_sc_hd__clkbuf_4
Xfanout243 _12394_/A vssd1 vssd1 vccd1 vccd1 _11886_/A sky130_fd_sc_hd__buf_4
Xfanout254 _09159_/X vssd1 vssd1 vccd1 vccd1 _12402_/A0 sky130_fd_sc_hd__clkbuf_4
Xfanout287 _06586_/X vssd1 vssd1 vccd1 vccd1 _06694_/B sky130_fd_sc_hd__clkbuf_8
Xfanout276 _13213_/B2 vssd1 vssd1 vccd1 vccd1 _13016_/A2 sky130_fd_sc_hd__buf_2
Xfanout298 _13242_/A vssd1 vssd1 vccd1 vccd1 _13235_/A sky130_fd_sc_hd__buf_4
X_09808_ _09808_/A _09808_/B vssd1 vssd1 vccd1 vccd1 _10368_/A sky130_fd_sc_hd__xnor2_4
XANTENNA_fanout62_A _12846_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09739_ _10449_/A _09739_/B vssd1 vssd1 vccd1 vccd1 _09741_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_69_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07479__A2 _10167_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09873__B1 _11766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12750_ _12750_/A _12754_/A vssd1 vssd1 vccd1 vccd1 _12752_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_96_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12681_ _12681_/A _12689_/A vssd1 vssd1 vccd1 vccd1 _12683_/C sky130_fd_sc_hd__nand2_1
X_11701_ _11510_/X _11868_/A _11699_/Y vssd1 vssd1 vccd1 vccd1 _12026_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_127_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11632_ hold200/A _11632_/B vssd1 vssd1 vccd1 vccd1 _11720_/B sky130_fd_sc_hd__or2_1
XANTENNA__13242__A _13242_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11248__A2_N _11234_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07240__A _09445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11432__B1 _11876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13302_ _13307_/CLK hold179/X vssd1 vssd1 vccd1 vccd1 hold177/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11563_ _11908_/A _11563_/B vssd1 vssd1 vccd1 vccd1 _11564_/B sky130_fd_sc_hd__xor2_1
XANTENNA__10786__A2 _07087_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10514_ _09324_/X _09332_/X _11010_/S vssd1 vssd1 vccd1 vccd1 _10514_/X sky130_fd_sc_hd__mux2_1
X_11494_ _11394_/A _11393_/B _11391_/Y vssd1 vssd1 vccd1 vccd1 _11495_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_18_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13233_ _12959_/B _13233_/B vssd1 vssd1 vccd1 vccd1 _13233_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__12292__S _12388_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10445_ _10445_/A _10941_/B vssd1 vssd1 vccd1 vccd1 _10448_/B sky130_fd_sc_hd__or2_1
X_13164_ _12883_/X _13164_/B vssd1 vssd1 vccd1 vccd1 _13165_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__09167__A _09168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10376_ _06760_/Y _10241_/Y _06762_/B vssd1 vssd1 vccd1 vccd1 _10376_/X sky130_fd_sc_hd__o21a_1
X_12115_ reg1_val[25] curr_PC[25] vssd1 vssd1 vccd1 vccd1 _12115_/X sky130_fd_sc_hd__and2_1
X_13095_ _13245_/A hold245/X vssd1 vssd1 vccd1 vccd1 _13348_/D sky130_fd_sc_hd__and2_1
X_12046_ hold265/A _12046_/B vssd1 vssd1 vccd1 vccd1 _12119_/B sky130_fd_sc_hd__or2_1
XANTENNA__09614__B _10963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08116__B1 _07955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12948_ _13202_/A _12947_/B _12871_/X vssd1 vssd1 vccd1 vccd1 _13207_/A sky130_fd_sc_hd__a21o_1
XANTENNA__07134__B _07135_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12879_ hold263/X hold21/X vssd1 vssd1 vccd1 vccd1 _13179_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_75_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07150__A _07343_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09616__B1 _11987_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08070_ _08874_/A _08874_/B _08050_/Y vssd1 vssd1 vccd1 vccd1 _08078_/B sky130_fd_sc_hd__a21boi_1
XFILLER_0_102_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09919__A1 _12810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09919__B2 _10413_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07021_ _07254_/B _06998_/B _12726_/B _07364_/B1 vssd1 vssd1 vccd1 vccd1 _07022_/B
+ sky130_fd_sc_hd__o31a_2
XFILLER_0_30_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09395__A2 _07099_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08972_ _09060_/A _08972_/B _09072_/B _09075_/A vssd1 vssd1 vccd1 vccd1 _08977_/A
+ sky130_fd_sc_hd__nand4_2
Xhold18 hold18/A vssd1 vssd1 vccd1 vccd1 hold18/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 hold29/A vssd1 vssd1 vccd1 vccd1 hold29/X sky130_fd_sc_hd__dlygate4sd3_1
X_07923_ _07923_/A _07923_/B vssd1 vssd1 vccd1 vccd1 _08029_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07854_ _07854_/A _07854_/B _07854_/C vssd1 vssd1 vccd1 vccd1 _07969_/A sky130_fd_sc_hd__and3_1
X_06805_ _06805_/A _12629_/B vssd1 vssd1 vccd1 vccd1 _06805_/X sky130_fd_sc_hd__and2_1
XANTENNA__10162__B1 _08507_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07785_ _08656_/B _08038_/B _08038_/C _11558_/A _08732_/A2 vssd1 vssd1 vccd1 vccd1
+ _07786_/B sky130_fd_sc_hd__o32a_1
X_06736_ reg1_val[11] _06963_/A vssd1 vssd1 vccd1 vccd1 _06737_/B sky130_fd_sc_hd__nor2_1
X_09524_ _06809_/X _09523_/Y _12388_/S vssd1 vssd1 vccd1 vccd1 _09525_/B sky130_fd_sc_hd__mux2_1
XANTENNA__08658__A1 _08733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06667_ reg1_val[20] _07220_/A vssd1 vssd1 vccd1 vccd1 _11727_/A sky130_fd_sc_hd__and2_1
X_09455_ _09906_/A _09455_/B vssd1 vssd1 vccd1 vccd1 _09456_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__07330__B2 _09567_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07330__A1 _12842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08406_ _08434_/A _08434_/B _08402_/Y vssd1 vssd1 vccd1 vccd1 _08419_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_47_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06598_ instruction[41] _06596_/A _06596_/B _06585_/X vssd1 vssd1 vccd1 vccd1 _07064_/B
+ sky130_fd_sc_hd__a31o_4
X_09386_ _09386_/A _09386_/B vssd1 vssd1 vccd1 vccd1 _09389_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_46_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12206__A2 fanout12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08156__A _08724_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08337_ _08335_/A _08335_/B _08336_/X vssd1 vssd1 vccd1 vccd1 _08381_/B sky130_fd_sc_hd__o21ba_1
X_08268_ _08728_/A _08268_/B vssd1 vssd1 vccd1 vccd1 _08329_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_116_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07219_ _07220_/B _07220_/C _07220_/A vssd1 vssd1 vccd1 vccd1 _08038_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_21_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10230_ _10231_/A _10231_/B vssd1 vssd1 vccd1 vccd1 _10230_/X sky130_fd_sc_hd__and2_1
XFILLER_0_30_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08199_ _08197_/A _08197_/B _08246_/A vssd1 vssd1 vccd1 vccd1 _08214_/A sky130_fd_sc_hd__o21ai_2
X_10161_ _10941_/B _10589_/A vssd1 vssd1 vccd1 vccd1 _10164_/B sky130_fd_sc_hd__or2_1
X_10092_ _10092_/A _10092_/B vssd1 vssd1 vccd1 vccd1 _10093_/B sky130_fd_sc_hd__xor2_4
X_12802_ _12802_/A _12818_/B vssd1 vssd1 vccd1 vccd1 _12802_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_97_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10994_ _11424_/A _10995_/C _11100_/B vssd1 vssd1 vccd1 vccd1 _10996_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_96_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09450__A _11384_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12733_ reg1_val[20] _12741_/B _12729_/A vssd1 vssd1 vccd1 vccd1 _12734_/B sky130_fd_sc_hd__a21oi_4
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12664_ reg1_val[8] _12664_/B vssd1 vssd1 vccd1 vccd1 _12665_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_38_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12595_ _12595_/A _12595_/B vssd1 vssd1 vccd1 vccd1 _12596_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_53_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11615_ _11614_/A _11614_/B _12290_/A vssd1 vssd1 vccd1 vccd1 _11615_/Y sky130_fd_sc_hd__a21oi_1
X_11546_ hold200/A _11450_/B _11632_/B _11968_/B1 vssd1 vssd1 vccd1 vccd1 _11546_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_107_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07085__B1 _11261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08821__A1 _11758_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13216_ _13216_/A _13216_/B vssd1 vssd1 vccd1 vccd1 _13216_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__09609__B _09609_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12316__A _12316_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11477_ _11478_/A _11478_/B vssd1 vssd1 vccd1 vccd1 _11479_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_12_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10428_ _10428_/A _10428_/B vssd1 vssd1 vccd1 vccd1 _10430_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13147_ hold287/X _06890_/Y _13146_/X _13246_/B2 vssd1 vssd1 vccd1 vccd1 _13148_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__07129__B _11343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10359_ _10360_/A _10360_/B vssd1 vssd1 vccd1 vccd1 _10359_/X sky130_fd_sc_hd__and2_1
X_13078_ _13341_/Q _12791_/A _13080_/B1 hold113/X _13113_/A vssd1 vssd1 vccd1 vccd1
+ hold114/A sky130_fd_sc_hd__o221a_1
XFILLER_0_57_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09534__C1 _06924_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12029_ _12170_/A _12030_/B _12030_/C vssd1 vssd1 vccd1 vccd1 _12029_/X sky130_fd_sc_hd__a21o_1
XANTENNA__10144__B1 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10396__A2_N _12404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12436__A2 _07064_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_78 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07570_ _07504_/Y _07370_/Y _07570_/S vssd1 vssd1 vccd1 vccd1 _07571_/B sky130_fd_sc_hd__mux2_2
XANTENNA__06984__A _10448_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07799__B _08436_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09240_ _09241_/B _09241_/C _09441_/A vssd1 vssd1 vccd1 vccd1 _09242_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_75_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10998__A2 _10996_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07312__A1 fanout30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07312__B2 _07688_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07863__A2 _08744_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09171_ hold260/A _09167_/Y _09169_/Y hold290/A _09166_/X vssd1 vssd1 vccd1 vccd1
+ _09171_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_90_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07615__A2 _10589_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08122_ _08741_/B2 _08656_/B _12820_/A _08732_/A2 vssd1 vssd1 vccd1 vccd1 _08123_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_31_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08053_ _08436_/A fanout87/X fanout82/X fanout99/X vssd1 vssd1 vccd1 vccd1 _08054_/B
+ sky130_fd_sc_hd__o22a_1
X_07004_ _12341_/A _07064_/B _09351_/B vssd1 vssd1 vccd1 vccd1 _07006_/B sky130_fd_sc_hd__and3_2
XFILLER_0_3_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout112_A _07522_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08040__A2 _08041_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08955_ _09065_/B _09073_/B vssd1 vssd1 vccd1 vccd1 _08972_/B sky130_fd_sc_hd__nor2_1
X_07906_ _07966_/A _07966_/B _07880_/X vssd1 vssd1 vccd1 vccd1 _07908_/B sky130_fd_sc_hd__a21o_1
X_08886_ _09042_/B _09049_/A vssd1 vssd1 vccd1 vccd1 _08886_/X sky130_fd_sc_hd__and2_1
X_07837_ _07838_/A _07838_/B vssd1 vssd1 vccd1 vccd1 _07837_/X sky130_fd_sc_hd__and2b_1
XANTENNA__10686__B2 _10575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10686__A1 _10574_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07768_ _07768_/A _07768_/B vssd1 vssd1 vccd1 vccd1 _07769_/B sky130_fd_sc_hd__nand2_1
X_06719_ _11130_/S _06719_/B vssd1 vssd1 vccd1 vccd1 _11111_/A sky130_fd_sc_hd__nor2_1
X_09507_ _09505_/X _09506_/X _09974_/A vssd1 vssd1 vccd1 vccd1 _09507_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_78_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09270__A _11987_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07699_ _08731_/A _07699_/B vssd1 vssd1 vccd1 vccd1 _07794_/A sky130_fd_sc_hd__xnor2_1
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09438_ _09439_/B vssd1 vssd1 vccd1 vccd1 _09438_/Y sky130_fd_sc_hd__inv_2
XANTENNA_fanout25_A _09613_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09369_ _10119_/S _09368_/Y _09181_/X vssd1 vssd1 vccd1 vccd1 _12394_/B sky130_fd_sc_hd__o21ai_2
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12380_ _12380_/A _12380_/B _12380_/C _12413_/A vssd1 vssd1 vccd1 vccd1 _12380_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_35_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11400_ _11293_/B _11295_/B _11293_/A vssd1 vssd1 vccd1 vccd1 _11405_/A sky130_fd_sc_hd__o21bai_2
X_11331_ _11332_/A _11332_/B vssd1 vssd1 vccd1 vccd1 _11331_/X sky130_fd_sc_hd__or2_1
XFILLER_0_62_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11262_ _11263_/A _11263_/B vssd1 vssd1 vccd1 vccd1 _11394_/A sky130_fd_sc_hd__nor2_1
X_13001_ _13013_/A hold211/X vssd1 vssd1 vccd1 vccd1 _13303_/D sky130_fd_sc_hd__and2_1
XANTENNA__12363__A1 _06838_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10213_ _10213_/A _10213_/B vssd1 vssd1 vccd1 vccd1 _10214_/B sky130_fd_sc_hd__xnor2_4
X_11193_ _11078_/A _11077_/B _11075_/X vssd1 vssd1 vccd1 vccd1 _11198_/A sky130_fd_sc_hd__a21o_1
XANTENNA__09445__A _09445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10144_ _10413_/A _10797_/B fanout5/X _12810_/A vssd1 vssd1 vccd1 vccd1 _10145_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_118_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06788__B _11118_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10075_ _10076_/A _10076_/B _10076_/C vssd1 vssd1 vccd1 vccd1 _10075_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__09531__A2 _11343_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07542__B2 _07075_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07542__A1 _10664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10977_ _11088_/B _10977_/B vssd1 vssd1 vccd1 vccd1 _10979_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_128_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12716_ reg1_val[18] _12741_/B vssd1 vssd1 vccd1 vccd1 _12718_/A sky130_fd_sc_hd__or2_1
XFILLER_0_128_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12647_ _12646_/A _12643_/Y _12645_/B vssd1 vssd1 vccd1 vccd1 _12651_/A sky130_fd_sc_hd__o21a_2
XFILLER_0_26_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12051__B1 _09152_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07058__B1 _07200_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12578_ _12611_/A _12579_/B vssd1 vssd1 vccd1 vccd1 _12580_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_53_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11529_ reg1_val[18] curr_PC[18] vssd1 vssd1 vccd1 vccd1 _11532_/A sky130_fd_sc_hd__or2_1
XFILLER_0_41_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_45 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08740_ _08740_/A _08740_/B vssd1 vssd1 vccd1 vccd1 _08743_/A sky130_fd_sc_hd__xnor2_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09522__A2 _09505_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08671_ _08730_/A1 _07821_/A _08436_/B _08671_/B2 vssd1 vssd1 vccd1 vccd1 _08672_/B
+ sky130_fd_sc_hd__o22a_1
X_07622_ _07983_/A _07983_/B vssd1 vssd1 vccd1 vccd1 _07984_/A sky130_fd_sc_hd__or2_1
XANTENNA__08730__B1 _08038_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13082__A2 _06572_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07553_ _07564_/A _07564_/B _07549_/X vssd1 vssd1 vccd1 vccd1 _07555_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_124_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07484_ _12824_/A _10941_/A _07076_/Y _12826_/A vssd1 vssd1 vccd1 vccd1 _07485_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07297__B1 _10022_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09223_ _09224_/B _09223_/B vssd1 vssd1 vccd1 vccd1 _09415_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_91_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09154_ _09170_/B _09159_/B vssd1 vssd1 vccd1 vccd1 _09154_/Y sky130_fd_sc_hd__nor2_4
XFILLER_0_90_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07049__B1 _09147_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08105_ _08106_/A _08106_/B vssd1 vssd1 vccd1 vccd1 _08765_/A sky130_fd_sc_hd__or2_1
X_09085_ reg1_val[1] reg1_val[30] _09108_/S vssd1 vssd1 vccd1 vccd1 _09085_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_71_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08261__A2 _08732_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08036_ _10927_/A1 _08732_/A2 _08656_/B _11367_/A vssd1 vssd1 vccd1 vccd1 _08037_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_3_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09265__A _11146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09987_ _09843_/A _09840_/Y _09842_/B vssd1 vssd1 vccd1 vccd1 _09991_/A sky130_fd_sc_hd__o21a_1
X_08938_ _08939_/A _08939_/B vssd1 vssd1 vccd1 vccd1 _09073_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_98_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08869_ _08869_/A _08869_/B vssd1 vssd1 vccd1 vccd1 _09042_/B sky130_fd_sc_hd__xor2_4
X_10900_ _10119_/S _09671_/X _09181_/X vssd1 vssd1 vccd1 vccd1 _11630_/B sky130_fd_sc_hd__o21a_1
XANTENNA__08721__B1 _08721_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13058__C1 _13128_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11880_ _11880_/A _11880_/B vssd1 vssd1 vccd1 vccd1 _11880_/Y sky130_fd_sc_hd__xnor2_1
X_10831_ _10961_/A _10961_/B vssd1 vssd1 vccd1 vccd1 _10833_/A sky130_fd_sc_hd__nor2_1
X_10762_ _09820_/Y _10761_/Y _11233_/S vssd1 vssd1 vccd1 vccd1 _10762_/X sky130_fd_sc_hd__mux2_1
XANTENNA__07288__B1 _12067_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12501_ _12502_/A _12502_/B _12502_/C vssd1 vssd1 vccd1 vccd1 _12509_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_82_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12432_ hold109/A _12431_/X _09167_/Y vssd1 vssd1 vccd1 vccd1 _12432_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_109_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10693_ _10693_/A _10693_/B vssd1 vssd1 vccd1 vccd1 _10694_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_105_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12363_ _06838_/B _11343_/B _12339_/Y _12362_/X _12455_/S vssd1 vssd1 vccd1 vccd1
+ dest_val[29] sky130_fd_sc_hd__o221a_4
XFILLER_0_23_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12294_ _12293_/A _12293_/B _12293_/Y _09156_/Y vssd1 vssd1 vccd1 vccd1 _12312_/A
+ sky130_fd_sc_hd__o211a_1
X_11314_ _11315_/A _11315_/B _11315_/C vssd1 vssd1 vccd1 vccd1 _11316_/A sky130_fd_sc_hd__a21o_1
X_11245_ _12307_/B1 _11244_/X _06713_/B vssd1 vssd1 vccd1 vccd1 _11245_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__09201__B2 _07688_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09201__A1 fanout30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10898__A1 _12307_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07763__A1 _08732_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11176_ _11177_/A _11177_/B _11177_/C vssd1 vssd1 vccd1 vccd1 _11176_/Y sky130_fd_sc_hd__a21oi_1
X_10127_ _07036_/A _12404_/A _11973_/B _06769_/B _10126_/Y vssd1 vssd1 vccd1 vccd1
+ _10127_/X sky130_fd_sc_hd__a221o_1
XANTENNA__07763__B2 _10927_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10058_ _10059_/A _10059_/B vssd1 vssd1 vccd1 vccd1 _10218_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_89_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07279__B1 _10571_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09440__A1 _12852_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold104 hold111/X vssd1 vssd1 vccd1 vccd1 hold104/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold115 hold115/A vssd1 vssd1 vccd1 vccd1 hold115/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold126 hold126/A vssd1 vssd1 vccd1 vccd1 hold126/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09440__B2 _12854_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold159 hold159/A vssd1 vssd1 vccd1 vccd1 hold159/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold148 hold148/A vssd1 vssd1 vccd1 vccd1 hold148/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold137 hold137/A vssd1 vssd1 vccd1 vccd1 hold137/X sky130_fd_sc_hd__dlygate4sd3_1
X_09910_ _09910_/A _09910_/B vssd1 vssd1 vccd1 vccd1 _09911_/B sky130_fd_sc_hd__and2_1
XFILLER_0_0_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11535__C1 _06924_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10889__A1 _12244_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09841_ reg1_val[4] curr_PC[4] vssd1 vssd1 vccd1 vccd1 _09842_/B sky130_fd_sc_hd__nand2_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09772_ _09772_/A _09772_/B vssd1 vssd1 vccd1 vccd1 _09774_/B sky130_fd_sc_hd__xnor2_2
X_06984_ _10448_/A _10949_/A _06986_/B vssd1 vssd1 vccd1 vccd1 _06985_/B sky130_fd_sc_hd__nand3_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08723_ fanout75/X _07896_/A _08723_/B1 _08304_/B vssd1 vssd1 vccd1 vccd1 _08724_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout277_A hold65/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10959__A _10959_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08654_ _08650_/A _08650_/C _08650_/B vssd1 vssd1 vccd1 vccd1 _08689_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__13055__A2 _13087_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08585_ _08613_/A _08592_/B _08578_/X vssd1 vssd1 vccd1 vccd1 _08609_/A sky130_fd_sc_hd__a21o_1
X_07605_ _10664_/A fanout94/X _10567_/A fanout69/X vssd1 vssd1 vccd1 vccd1 _07606_/B
+ sky130_fd_sc_hd__o22a_1
X_07536_ _09400_/A _10567_/A vssd1 vssd1 vccd1 vccd1 _07537_/C sky130_fd_sc_hd__or2_1
XANTENNA__07052__B _11987_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11066__B2 _09745_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11066__A1 _10418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09206_ _09469_/A _09206_/B vssd1 vssd1 vccd1 vccd1 _09208_/B sky130_fd_sc_hd__or2_2
X_07467_ _07468_/B _07569_/A vssd1 vssd1 vccd1 vccd1 _09205_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_76_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07398_ _07398_/A _07398_/B vssd1 vssd1 vccd1 vccd1 _08958_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_63_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08164__A _11385_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09137_ _09133_/X _09136_/X _09663_/S vssd1 vssd1 vccd1 vccd1 _09137_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_44_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07442__B1 _12810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09068_ _09060_/A _08972_/B _08975_/Y vssd1 vssd1 vccd1 vccd1 _09069_/B sky130_fd_sc_hd__a21boi_2
XFILLER_0_44_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10577__B1 _11180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08019_ _08019_/A _08019_/B vssd1 vssd1 vccd1 vccd1 _08021_/B sky130_fd_sc_hd__xnor2_2
XANTENNA_fanout92_A _07833_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10329__B1 _10575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11030_ curr_PC[13] _11139_/C _10780_/A vssd1 vssd1 vccd1 vccd1 _11030_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__09734__A2 _10589_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07508__A _10928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11541__A2 _09527_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12981_ _13013_/A hold231/X vssd1 vssd1 vccd1 vccd1 _13293_/D sky130_fd_sc_hd__and2_1
XFILLER_0_99_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10501__B1 _10500_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11932_ _11932_/A _11932_/B vssd1 vssd1 vccd1 vccd1 _11934_/B sky130_fd_sc_hd__nor2_1
XANTENNA__08170__A1 _08752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13046__A2 _12788_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08170__B2 _08798_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11863_ _11863_/A _11863_/B vssd1 vssd1 vccd1 vccd1 _12165_/A sky130_fd_sc_hd__nand2_2
X_10814_ _10971_/A _10814_/B _10814_/C vssd1 vssd1 vccd1 vccd1 _10971_/B sky130_fd_sc_hd__and3b_1
XANTENNA__11057__A1 fanout66/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11057__B2 _07087_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11794_ _06676_/C _11710_/Y _11727_/A vssd1 vssd1 vccd1 vccd1 _11794_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_67_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10745_ _10782_/B vssd1 vssd1 vccd1 vccd1 _11033_/C sky130_fd_sc_hd__inv_2
XFILLER_0_55_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10676_ _10676_/A _10676_/B vssd1 vssd1 vccd1 vccd1 _10677_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_125_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13395_ instruction[4] vssd1 vssd1 vccd1 vccd1 sign_extend sky130_fd_sc_hd__buf_12
XFILLER_0_63_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12415_ _12330_/B _12374_/A _12376_/B vssd1 vssd1 vccd1 vccd1 _12415_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_105_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12346_ _12426_/A _09077_/A _09077_/B vssd1 vssd1 vccd1 vccd1 _12346_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_50_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12309__A1 _09111_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12309__B2 _09152_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12277_ _12277_/A _12277_/B _12277_/C vssd1 vssd1 vccd1 vccd1 _12278_/B sky130_fd_sc_hd__or3_1
XFILLER_0_10_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11228_ _11226_/Y _11228_/B vssd1 vssd1 vccd1 vccd1 _11230_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_65_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07736__B2 _08432_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07736__A1 _10537_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11159_ _11160_/A _11160_/B vssd1 vssd1 vccd1 vccd1 _11159_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08370_ _08370_/A _08370_/B vssd1 vssd1 vccd1 vccd1 _08372_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_85_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07321_ _07322_/A _07322_/B vssd1 vssd1 vccd1 vccd1 _07573_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_58_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07252_ _07300_/B _07300_/A vssd1 vssd1 vccd1 vccd1 _07267_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_61_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07183_ reg1_val[7] _07183_/B vssd1 vssd1 vccd1 vccd1 _07183_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_53_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09808__A _09808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09527__B _09527_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09824_ _11231_/S _09824_/B vssd1 vssd1 vccd1 vccd1 _09824_/X sky130_fd_sc_hd__or2_1
XANTENNA__07047__B _11987_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06967_ _11020_/A _07074_/A _06967_/C _06967_/D vssd1 vssd1 vccd1 vccd1 _07133_/B
+ sky130_fd_sc_hd__or4_2
X_09755_ _09755_/A _09755_/B vssd1 vssd1 vccd1 vccd1 _09764_/A sky130_fd_sc_hd__xor2_2
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06898_ instruction[11] _06902_/B vssd1 vssd1 vccd1 vccd1 dest_idx[0] sky130_fd_sc_hd__and2_4
X_09686_ _09687_/B _09686_/B vssd1 vssd1 vccd1 vccd1 _09686_/Y sky130_fd_sc_hd__nand2b_1
X_08706_ _09008_/A _09008_/B _09018_/B _08542_/Y vssd1 vssd1 vccd1 vccd1 _08707_/B
+ sky130_fd_sc_hd__a211o_1
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08637_ _08637_/A _08637_/B vssd1 vssd1 vccd1 vccd1 _08652_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_69_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13028__A2 _12788_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08568_ _08575_/A _08575_/B _08561_/X vssd1 vssd1 vccd1 vccd1 _08572_/B sky130_fd_sc_hd__a21oi_1
Xfanout21 _07099_/X vssd1 vssd1 vccd1 vccd1 _09609_/B sky130_fd_sc_hd__clkbuf_8
Xfanout10 fanout9/A vssd1 vssd1 vccd1 vccd1 _10797_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_0_119_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10628__S _12174_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07519_ _07519_/A _07519_/B vssd1 vssd1 vccd1 vccd1 _07520_/B sky130_fd_sc_hd__or2_1
X_08499_ _08584_/A _08499_/B vssd1 vssd1 vccd1 vccd1 _08501_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_76_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout32 _12412_/B vssd1 vssd1 vccd1 vccd1 _12316_/B sky130_fd_sc_hd__clkbuf_8
Xfanout43 _07221_/X vssd1 vssd1 vccd1 vccd1 _12834_/A sky130_fd_sc_hd__clkbuf_8
Xfanout54 _12842_/A vssd1 vssd1 vccd1 vccd1 _10571_/B sky130_fd_sc_hd__buf_4
Xfanout65 _09745_/A vssd1 vssd1 vccd1 vccd1 _09396_/B sky130_fd_sc_hd__buf_6
XFILLER_0_49_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10798__B1 _10959_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10530_ _06924_/X _10517_/X _10529_/X _10508_/X vssd1 vssd1 vccd1 vccd1 _10530_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_92_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout87 _07204_/X vssd1 vssd1 vccd1 vccd1 fanout87/X sky130_fd_sc_hd__buf_6
Xfanout98 fanout99/X vssd1 vssd1 vccd1 vccd1 _10664_/A sky130_fd_sc_hd__clkbuf_8
Xfanout76 _09548_/A vssd1 vssd1 vccd1 vccd1 _12317_/A sky130_fd_sc_hd__buf_8
XFILLER_0_107_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10461_ fanout74/X _12214_/A fanout59/X _10948_/B2 vssd1 vssd1 vccd1 vccd1 _10462_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__13200__A2 _13213_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12200_ _12172_/X _12177_/X _12180_/X _12199_/X _06881_/X vssd1 vssd1 vccd1 vccd1
+ _12200_/X sky130_fd_sc_hd__a41o_1
XFILLER_0_44_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11907__A_N _11908_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13180_ _13180_/A _13180_/B vssd1 vssd1 vccd1 vccd1 _13180_/Y sky130_fd_sc_hd__xnor2_1
X_10392_ _06756_/B _09158_/Y _09154_/Y vssd1 vssd1 vccd1 vccd1 _10392_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__07415__B1 _12852_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12131_ _06924_/X _12118_/X _12130_/X _12111_/X vssd1 vssd1 vccd1 vccd1 _12131_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07238__A _09442_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12062_ _12213_/A fanout9/X fanout4/X _12150_/A vssd1 vssd1 vccd1 vccd1 _12063_/B
+ sky130_fd_sc_hd__o22a_1
X_11013_ _11886_/A _11009_/X _11012_/Y _09172_/B vssd1 vssd1 vccd1 vccd1 _11013_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_126_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12964_ hold248/A _13213_/B2 _13213_/A2 hold238/X vssd1 vssd1 vccd1 vccd1 hold239/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09172__B _09172_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11278__A1 _07819_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11278__B2 fanout24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08143__A1 _08741_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08143__B2 _08732_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11915_ _11915_/A _11915_/B vssd1 vssd1 vccd1 vccd1 _11916_/B sky130_fd_sc_hd__nand2_1
X_12895_ hold33/X hold288/A vssd1 vssd1 vccd1 vccd1 _12895_/X sky130_fd_sc_hd__and2b_1
XTAP_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11846_ _11846_/A _11846_/B vssd1 vssd1 vccd1 vccd1 _11847_/C sky130_fd_sc_hd__xnor2_1
XTAP_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07701__A _08728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11777_ _11777_/A _11777_/B vssd1 vssd1 vccd1 vccd1 _11779_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_125_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10728_ _10729_/A _10729_/B vssd1 vssd1 vccd1 vccd1 _10854_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_27_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10659_ _11033_/A _11033_/B vssd1 vssd1 vccd1 vccd1 _10782_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_51_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13378_ _13378_/CLK _13378_/D vssd1 vssd1 vccd1 vccd1 hold109/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07406__B1 _08216_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12329_ _12327_/A _12327_/B _12327_/C vssd1 vssd1 vccd1 vccd1 _12330_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_11_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07148__A _07149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07709__B2 _09768_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07709__A1 _12804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07870_ _08038_/A _11847_/A _11923_/A _08730_/A1 vssd1 vssd1 vccd1 vccd1 _07871_/B
+ sky130_fd_sc_hd__o22a_1
X_06821_ _11004_/A _06820_/X _06722_/Y vssd1 vssd1 vccd1 vccd1 _06821_/X sky130_fd_sc_hd__o21a_1
XANTENNA__06932__A2 _12341_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06752_ _06805_/A _06702_/A _12669_/B _06751_/X vssd1 vssd1 vccd1 vccd1 _07089_/A
+ sky130_fd_sc_hd__a31o_4
X_09540_ curr_PC[0] curr_PC[1] curr_PC[2] vssd1 vssd1 vccd1 vccd1 _09540_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_92_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09471_ _09281_/A _09281_/B _09279_/Y vssd1 vssd1 vccd1 vccd1 _09473_/B sky130_fd_sc_hd__a21bo_2
X_06683_ _11638_/A _06683_/B vssd1 vssd1 vccd1 vccd1 _06866_/A sky130_fd_sc_hd__nor2_1
XANTENNA__09882__A1 _08632_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08422_ _08422_/A _08422_/B vssd1 vssd1 vccd1 vccd1 _08454_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_86_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout142_A _10148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08353_ _08745_/A _08353_/B vssd1 vssd1 vccd1 vccd1 _08413_/B sky130_fd_sc_hd__xnor2_1
X_07304_ _07628_/A _07628_/B _07301_/X vssd1 vssd1 vccd1 vccd1 _07674_/A sky130_fd_sc_hd__a21oi_4
X_08284_ _08284_/A _08284_/B vssd1 vssd1 vccd1 vccd1 _08288_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_6_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07235_ _12842_/A _09440_/B1 _12840_/A _09238_/B vssd1 vssd1 vccd1 vccd1 _07236_/B
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_61_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07166_ _07166_/A _07166_/B vssd1 vssd1 vccd1 vccd1 _07166_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_14_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07097_ _11384_/A _09746_/A _11470_/B vssd1 vssd1 vccd1 vccd1 _07099_/A sky130_fd_sc_hd__or3b_4
XFILLER_0_2_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout200 _12790_/Y vssd1 vssd1 vccd1 vccd1 _12856_/B sky130_fd_sc_hd__buf_4
Xfanout222 _12789_/B vssd1 vssd1 vccd1 vccd1 _06892_/B sky130_fd_sc_hd__clkbuf_8
Xfanout211 _09898_/A vssd1 vssd1 vccd1 vccd1 _09441_/A sky130_fd_sc_hd__buf_12
Xfanout244 _06771_/X vssd1 vssd1 vccd1 vccd1 _12394_/A sky130_fd_sc_hd__buf_4
Xfanout233 _06794_/X vssd1 vssd1 vccd1 vccd1 _10250_/S sky130_fd_sc_hd__clkbuf_8
Xfanout255 _09157_/X vssd1 vssd1 vccd1 vccd1 _11624_/A sky130_fd_sc_hd__buf_4
XFILLER_0_5_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout288 _06586_/X vssd1 vssd1 vccd1 vccd1 _06634_/B sky130_fd_sc_hd__clkbuf_4
Xfanout277 hold65/X vssd1 vssd1 vccd1 vccd1 _13213_/B2 sky130_fd_sc_hd__buf_4
Xfanout266 _06882_/Y vssd1 vssd1 vccd1 vccd1 _12455_/S sky130_fd_sc_hd__clkbuf_16
Xfanout299 _13109_/A vssd1 vssd1 vccd1 vccd1 _13113_/A sky130_fd_sc_hd__buf_4
X_09807_ _09808_/A _09808_/B vssd1 vssd1 vccd1 vccd1 _09807_/X sky130_fd_sc_hd__and2_1
X_07999_ _07999_/A _07999_/B vssd1 vssd1 vccd1 vccd1 _08000_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_5_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09738_ fanout59/X _10167_/A1 _10022_/B1 _10941_/B vssd1 vssd1 vccd1 vccd1 _09739_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_96_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09669_ _09333_/X _09335_/X _09669_/S vssd1 vssd1 vccd1 vccd1 _09669_/X sky130_fd_sc_hd__mux2_1
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09873__B2 fanout94/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09873__A1 _10941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08617__A _08673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12680_ reg1_val[11] _12680_/B vssd1 vssd1 vccd1 vccd1 _12689_/A sky130_fd_sc_hd__nand2_1
X_11700_ _11700_/A _11700_/B _11700_/C vssd1 vssd1 vccd1 vccd1 _11868_/A sky130_fd_sc_hd__or3_1
XANTENNA__11680__A1 _11564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07884__B1 _09768_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11631_ _12394_/A _11629_/Y _11630_/X _09172_/B vssd1 vssd1 vccd1 vccd1 _11644_/B
+ sky130_fd_sc_hd__o211a_1
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11562_ _09613_/A fanout56/X _12316_/A _09614_/A vssd1 vssd1 vccd1 vccd1 _11563_/B
+ sky130_fd_sc_hd__o22a_1
X_13301_ _13307_/CLK hold202/X vssd1 vssd1 vccd1 vccd1 hold200/A sky130_fd_sc_hd__dfxtp_1
X_10513_ _10513_/A _10513_/B vssd1 vssd1 vccd1 vccd1 _10513_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_80_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10786__A3 _10570_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10640__C1 _09172_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11493_ _11381_/A _11381_/B _11378_/A vssd1 vssd1 vccd1 vccd1 _11495_/A sky130_fd_sc_hd__a21o_1
X_13232_ _13235_/A hold251/X vssd1 vssd1 vccd1 vccd1 _13377_/D sky130_fd_sc_hd__and2_1
XANTENNA__09448__A _10707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10444_ _10444_/A _10444_/B vssd1 vssd1 vccd1 vccd1 _10452_/A sky130_fd_sc_hd__xnor2_1
X_13163_ _13245_/A hold272/X vssd1 vssd1 vccd1 vccd1 _13362_/D sky130_fd_sc_hd__and2_1
XANTENNA__09167__B _09170_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10375_ _09653_/A _08996_/A _08996_/B _09163_/X vssd1 vssd1 vccd1 vccd1 _10375_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_32_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12114_ reg1_val[25] curr_PC[25] vssd1 vssd1 vccd1 vccd1 _12114_/X sky130_fd_sc_hd__or2_1
XFILLER_0_32_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13094_ hold244/X _06892_/B _13093_/X _06572_/A vssd1 vssd1 vccd1 vccd1 hold245/A
+ sky130_fd_sc_hd__a22o_1
X_12045_ hold218/A _12434_/B1 _12123_/B _12401_/B1 vssd1 vssd1 vccd1 vccd1 _12045_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_46_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12448__A0 _09343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08116__A1 _08304_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08116__B2 fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12947_ _12871_/X _12947_/B vssd1 vssd1 vccd1 vccd1 _13202_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_99_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12878_ hold21/X hold263/X vssd1 vssd1 vccd1 vccd1 _12878_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_87_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07431__A _10165_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11829_ _12210_/A _11829_/B vssd1 vssd1 vccd1 vccd1 _11830_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_127_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11974__A2 _09527_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07020_ _07254_/B _12726_/B _07364_/B1 vssd1 vssd1 vccd1 vccd1 _07084_/B sky130_fd_sc_hd__o21ai_2
XANTENNA__08262__A _08733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08971_ _08971_/A _08971_/B vssd1 vssd1 vccd1 vccd1 _09649_/B sky130_fd_sc_hd__xnor2_2
Xhold19 hold19/A vssd1 vssd1 vccd1 vccd1 hold19/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12512__A _12673_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07922_ _07923_/A _07923_/B vssd1 vssd1 vccd1 vccd1 _07922_/Y sky130_fd_sc_hd__nor2_1
X_07853_ _07853_/A _07853_/B vssd1 vssd1 vccd1 vccd1 _07854_/C sky130_fd_sc_hd__xor2_1
XANTENNA__07606__A _11470_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10162__A1 _07154_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06804_ _09343_/A _09666_/S vssd1 vssd1 vccd1 vccd1 _09350_/A sky130_fd_sc_hd__xnor2_2
X_07784_ _07784_/A _07784_/B vssd1 vssd1 vccd1 vccd1 _07978_/A sky130_fd_sc_hd__xor2_1
X_06735_ reg1_val[11] _06963_/A vssd1 vssd1 vccd1 vccd1 _10767_/S sky130_fd_sc_hd__and2_1
X_09523_ _09523_/A _09523_/B vssd1 vssd1 vccd1 vccd1 _09523_/Y sky130_fd_sc_hd__nand2_1
X_06666_ _06664_/Y _06703_/B1 _06771_/A reg2_val[20] vssd1 vssd1 vccd1 vccd1 _07220_/A
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_66_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09454_ fanout75/X _10574_/B _10575_/B _06986_/Y vssd1 vssd1 vccd1 vccd1 _09455_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_93_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07330__A2 _09568_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09385_ _09385_/A _09385_/B vssd1 vssd1 vccd1 vccd1 _09386_/B sky130_fd_sc_hd__nand2_1
X_08405_ _08405_/A _08405_/B vssd1 vssd1 vccd1 vccd1 _08434_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06597_ _06575_/Y _06596_/Y _06585_/X vssd1 vssd1 vccd1 vccd1 _07420_/A sky130_fd_sc_hd__o21ba_2
XFILLER_0_47_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08336_ _08347_/B _08347_/A vssd1 vssd1 vccd1 vccd1 _08336_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_74_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07094__A1 _07089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08267_ _12818_/A _08727_/A2 _08727_/B1 _12820_/A vssd1 vssd1 vccd1 vccd1 _08268_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_15_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13167__B2 _13246_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07218_ _10320_/A _10321_/A _08584_/A vssd1 vssd1 vccd1 vccd1 _07218_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09268__A _10574_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08198_ _08245_/A _08245_/B vssd1 vssd1 vccd1 vccd1 _08246_/A sky130_fd_sc_hd__or2_1
X_07149_ _07149_/A _09343_/A vssd1 vssd1 vccd1 vccd1 _07149_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_42_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08043__B1 _11558_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10160_ _10019_/A _10019_/B _10015_/X vssd1 vssd1 vccd1 vccd1 _10172_/A sky130_fd_sc_hd__o21ai_1
X_10091_ _10092_/A _10092_/B vssd1 vssd1 vccd1 vccd1 _10091_/X sky130_fd_sc_hd__and2_1
XANTENNA__11038__A _12073_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12801_ _09598_/A _13077_/A2 hold89/X _13113_/A vssd1 vssd1 vccd1 vccd1 _13254_/D
+ sky130_fd_sc_hd__o211a_1
X_10993_ _10499_/A _10499_/B _10499_/C _10992_/X vssd1 vssd1 vccd1 vccd1 _10995_/C
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_96_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07857__B1 _08617_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12732_ _12730_/Y _12732_/B vssd1 vssd1 vccd1 vccd1 _12746_/B sky130_fd_sc_hd__nand2b_2
XFILLER_0_127_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07251__A _08584_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12663_ reg1_val[8] _12664_/B vssd1 vssd1 vccd1 vccd1 _12663_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_38_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12594_ _12579_/B _12587_/B _12611_/A vssd1 vssd1 vccd1 vccd1 _12607_/B sky130_fd_sc_hd__o21ai_2
X_11614_ _11614_/A _11614_/B vssd1 vssd1 vccd1 vccd1 _11614_/X sky130_fd_sc_hd__or2_1
X_11545_ _11450_/B _11632_/B hold200/A vssd1 vssd1 vccd1 vccd1 _11545_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_92_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07085__A1 _11269_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09178__A _11118_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11476_ _11476_/A _11476_/B vssd1 vssd1 vccd1 vccd1 _11478_/B sky130_fd_sc_hd__and2_1
XFILLER_0_122_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13215_ _12864_/X _13215_/B vssd1 vssd1 vccd1 vccd1 _13216_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__12316__B _12316_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10427_ _11180_/A _10427_/B vssd1 vssd1 vccd1 vccd1 _10428_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_110_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13146_ hold285/X _13145_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13146_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_103_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09906__A _09906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10358_ _10358_/A _10358_/B vssd1 vssd1 vccd1 vccd1 _10360_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_0_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13077_ _07013_/B _13077_/A2 hold68/X vssd1 vssd1 vccd1 vccd1 hold69/A sky130_fd_sc_hd__o21a_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10289_ _10149_/A _10149_/B _10146_/Y vssd1 vssd1 vccd1 vccd1 _10290_/B sky130_fd_sc_hd__o21a_1
XANTENNA__09117__S _09142_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12028_ _12162_/A _12028_/B vssd1 vssd1 vccd1 vccd1 _12030_/C sky130_fd_sc_hd__xor2_2
XANTENNA__10144__A1 _10413_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10144__B2 _12810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10787__A _11261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06984__B _10949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07312__A2 _09423_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08257__A _08722_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09170_ _09170_/A _09170_/B vssd1 vssd1 vccd1 vccd1 _09170_/X sky130_fd_sc_hd__or2_1
XFILLER_0_56_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08273__B1 _08617_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08121_ _08121_/A _08121_/B vssd1 vssd1 vccd1 vccd1 _08139_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_114_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08052_ _08742_/A _08052_/B vssd1 vssd1 vccd1 vccd1 _08055_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_114_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07003_ _12210_/A vssd1 vssd1 vccd1 vccd1 _11673_/A sky130_fd_sc_hd__inv_8
XANTENNA__10907__B1 _11142_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout105_A _11987_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08954_ _08954_/A _08954_/B vssd1 vssd1 vccd1 vccd1 _09073_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07336__A _08584_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07905_ _07905_/A _07905_/B vssd1 vssd1 vccd1 vccd1 _07966_/B sky130_fd_sc_hd__xnor2_2
X_08885_ _08885_/A _08885_/B vssd1 vssd1 vccd1 vccd1 _09049_/A sky130_fd_sc_hd__xnor2_2
X_07836_ _07836_/A _07836_/B vssd1 vssd1 vccd1 vccd1 _07838_/B sky130_fd_sc_hd__xor2_1
XANTENNA__10686__A2 _10575_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09828__A1 _09147_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12388__S _12388_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07767_ _07768_/A _07768_/B vssd1 vssd1 vccd1 vccd1 _07769_/A sky130_fd_sc_hd__or2_1
X_06718_ reg1_val[14] _06981_/A vssd1 vssd1 vccd1 vccd1 _06719_/B sky130_fd_sc_hd__nor2_1
X_09506_ _09121_/X _09125_/X _09669_/S vssd1 vssd1 vccd1 vccd1 _09506_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_79_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06894__B _06896_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07698_ _08436_/B _11989_/A fanout51/X _07149_/A vssd1 vssd1 vccd1 vccd1 _07699_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07071__A _11163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06649_ _06647_/X _06649_/B _06846_/A vssd1 vssd1 vccd1 vccd1 _06874_/A sky130_fd_sc_hd__nand3b_1
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09437_ _10449_/A _09437_/B vssd1 vssd1 vccd1 vccd1 _09439_/B sky130_fd_sc_hd__xnor2_1
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09368_ _11118_/A _09367_/A _09177_/Y vssd1 vssd1 vccd1 vccd1 _09368_/Y sky130_fd_sc_hd__a21oi_2
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09299_ _09299_/A _09299_/B vssd1 vssd1 vccd1 vccd1 _09302_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__12060__A1 _12455_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout18_A _12852_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08319_ _08742_/A _08319_/B vssd1 vssd1 vccd1 vccd1 _08322_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_19_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_60 instruction[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11330_ _06823_/X _11329_/X _12174_/S vssd1 vssd1 vccd1 vccd1 _11332_/B sky130_fd_sc_hd__mux2_1
XANTENNA__10071__B1 _10575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11261_ _11261_/A _11261_/B vssd1 vssd1 vccd1 vccd1 _11263_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_15_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13000_ hold177/X _13004_/A2 _13006_/B1 hold210/X vssd1 vssd1 vccd1 vccd1 hold211/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12363__A2 _11343_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10212_ _10210_/X _10212_/B vssd1 vssd1 vccd1 vccd1 _10213_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_30_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11192_ _11079_/A _11079_/B _11073_/A vssd1 vssd1 vccd1 vccd1 _11203_/A sky130_fd_sc_hd__a21oi_1
X_10143_ _10088_/A _10088_/B _10089_/X vssd1 vssd1 vccd1 vccd1 _10228_/A sky130_fd_sc_hd__o21bai_4
XANTENNA__11571__B1 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10074_ _10076_/A _10076_/B _10076_/C vssd1 vssd1 vccd1 vccd1 _10077_/A sky130_fd_sc_hd__o21a_1
XANTENNA__07542__A2 _11653_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10976_ _10976_/A _10976_/B _10976_/C vssd1 vssd1 vccd1 vccd1 _10977_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_84_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12715_ _12715_/A _12725_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[17] sky130_fd_sc_hd__xnor2_4
XFILLER_0_127_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12646_ _12646_/A _12646_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[4] sky130_fd_sc_hd__xnor2_4
XANTENNA__12051__A1 _07166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12577_ reg1_val[20] curr_PC[20] _12586_/S vssd1 vssd1 vccd1 vccd1 _12579_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_25_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11528_ _06693_/X _11524_/X _11526_/Y _11624_/A vssd1 vssd1 vccd1 vccd1 _11528_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_53_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11459_ _11360_/A _11649_/A _11649_/B _12031_/A vssd1 vssd1 vccd1 vccd1 _11519_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_7_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13158__A _13242_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13129_ _12897_/X _13129_/B vssd1 vssd1 vccd1 vccd1 _13130_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__09355__B _12341_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11562__B1 _12316_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07156__A _08645_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08670_ _08670_/A _08670_/B vssd1 vssd1 vccd1 vccd1 _08987_/A sky130_fd_sc_hd__nor2_1
X_07621_ _07621_/A _07621_/B vssd1 vssd1 vccd1 vccd1 _07983_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__08730__B2 _11558_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08730__A1 _08730_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07552_ _07552_/A _07552_/B vssd1 vssd1 vccd1 vccd1 _07564_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_88_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10310__A _12810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07483_ _10707_/A _07483_/B vssd1 vssd1 vccd1 vccd1 _07487_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__07297__A1 _11472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07297__B2 _11558_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09222_ _10449_/A _09222_/B vssd1 vssd1 vccd1 vccd1 _09224_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09153_ _12174_/S _09153_/B vssd1 vssd1 vccd1 vccd1 _09153_/Y sky130_fd_sc_hd__nand2_1
XANTENNA_fanout222_A _12789_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08104_ _08731_/A _08104_/B vssd1 vssd1 vccd1 vccd1 _08106_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_126_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09084_ _12423_/A _09153_/B vssd1 vssd1 vccd1 vccd1 _09127_/S sky130_fd_sc_hd__nand2_4
XFILLER_0_4_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08035_ _08034_/B _08034_/C _08034_/A vssd1 vssd1 vccd1 vccd1 _08069_/A sky130_fd_sc_hd__o21ba_1
XFILLER_0_3_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09986_ _09964_/A _12402_/A0 _09985_/X vssd1 vssd1 vccd1 vccd1 _09986_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__09265__B _09396_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08937_ _08937_/A _08937_/B vssd1 vssd1 vccd1 vccd1 _08939_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_98_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08868_ _08869_/A _08869_/B vssd1 vssd1 vccd1 vccd1 _08868_/X sky130_fd_sc_hd__and2_1
XFILLER_0_99_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07819_ _08752_/A _07819_/B vssd1 vssd1 vccd1 vccd1 _07824_/A sky130_fd_sc_hd__nor2_1
XANTENNA__08721__A1 _10537_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08721__B2 _08432_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08799_ _11758_/A _08799_/B vssd1 vssd1 vccd1 vccd1 _08801_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_67_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10830_ _10707_/A _06952_/Y _12412_/A _10829_/X vssd1 vssd1 vccd1 vccd1 _10961_/B
+ sky130_fd_sc_hd__a31o_1
X_10761_ _10761_/A vssd1 vssd1 vccd1 vccd1 _10761_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_94_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07288__B2 _09236_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07288__A1 _09444_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12500_ _12509_/A _12500_/B vssd1 vssd1 vccd1 vccd1 _12502_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_66_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10692_ _10693_/A _10693_/B vssd1 vssd1 vccd1 vccd1 _10835_/B sky130_fd_sc_hd__and2_1
XFILLER_0_125_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12431_ hold298/A _12396_/X _09835_/B vssd1 vssd1 vccd1 vccd1 _12431_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_82_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11051__A _11269_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12362_ _12362_/A _12362_/B _12362_/C _12361_/X vssd1 vssd1 vccd1 vccd1 _12362_/X
+ sky130_fd_sc_hd__or4b_1
X_12293_ _12293_/A _12293_/B vssd1 vssd1 vccd1 vccd1 _12293_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_50_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11313_ _11313_/A _11313_/B vssd1 vssd1 vccd1 vccd1 _11315_/C sky130_fd_sc_hd__xnor2_1
X_11244_ _09527_/B _09354_/B _11244_/S vssd1 vssd1 vccd1 vccd1 _11244_/X sky130_fd_sc_hd__mux2_1
XANTENNA__06799__B _06799_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09201__A2 _09768_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11175_ _11261_/A _11175_/B vssd1 vssd1 vccd1 vccd1 _11177_/C sky130_fd_sc_hd__xor2_1
X_10126_ hold242/A _11452_/B1 _10256_/B _10125_/Y _09837_/A vssd1 vssd1 vccd1 vccd1
+ _10126_/Y sky130_fd_sc_hd__a311oi_4
XFILLER_0_100_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07763__A2 fanout87/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10057_ _10218_/A _10057_/B vssd1 vssd1 vccd1 vccd1 _10059_/B sky130_fd_sc_hd__and2_1
XANTENNA__07704__A _12210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10568__A_N _10567_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07279__B2 _10664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07279__A1 _10570_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10959_ _10959_/A _10959_/B vssd1 vssd1 vccd1 vccd1 _10961_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_128_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12629_ reg1_val[1] _12629_/B vssd1 vssd1 vccd1 vccd1 _12630_/B sky130_fd_sc_hd__or2_1
XFILLER_0_14_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10035__B1 _10959_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08228__B1 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09440__A2 _09238_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold105 hold105/A vssd1 vssd1 vccd1 vccd1 hold105/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold116 hold126/X vssd1 vssd1 vccd1 vccd1 hold116/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold149 hold149/A vssd1 vssd1 vccd1 vccd1 hold149/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 hold138/A vssd1 vssd1 vccd1 vccd1 hold138/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold127 hold127/A vssd1 vssd1 vccd1 vccd1 hold127/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09840_ reg1_val[4] curr_PC[4] vssd1 vssd1 vccd1 vccd1 _09840_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__08400__B1 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10024__B fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09771_ _09771_/A _09771_/B vssd1 vssd1 vccd1 vccd1 _09772_/B sky130_fd_sc_hd__xnor2_2
X_06983_ _10448_/A _10949_/A _06986_/B vssd1 vssd1 vccd1 vccd1 _06985_/A sky130_fd_sc_hd__or3_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08722_ _08722_/A _08722_/B vssd1 vssd1 vccd1 vccd1 _08726_/A sky130_fd_sc_hd__xnor2_2
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12520__A _12680_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08653_ _08653_/A _08653_/B vssd1 vssd1 vccd1 vccd1 _08991_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08584_ _08584_/A _08584_/B vssd1 vssd1 vccd1 vccd1 _08592_/B sky130_fd_sc_hd__xnor2_2
X_07604_ _07604_/A _07604_/B vssd1 vssd1 vccd1 vccd1 _07624_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_76_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07535_ _07033_/A _07033_/B _10413_/A vssd1 vssd1 vccd1 vccd1 _07537_/B sky130_fd_sc_hd__a21o_1
XANTENNA__11066__A2 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07466_ _07434_/B _07437_/B _07434_/A vssd1 vssd1 vccd1 vccd1 _07468_/B sky130_fd_sc_hd__o21ba_1
X_09205_ _09205_/A _09205_/B _09205_/C vssd1 vssd1 vccd1 vccd1 _09206_/B sky130_fd_sc_hd__and3_1
XFILLER_0_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07397_ _07399_/A _07399_/B vssd1 vssd1 vccd1 vccd1 _07397_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_44_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09136_ _09134_/X _09135_/X _09336_/S vssd1 vssd1 vccd1 vccd1 _09136_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_115_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07442__B2 _11171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07442__A1 fanout23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09067_ _09072_/A _09067_/B vssd1 vssd1 vccd1 vccd1 _09077_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__09276__A _10422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08018_ _08019_/B _08019_/A vssd1 vssd1 vccd1 vccd1 _08018_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_4_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10329__A1 _10418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10329__B2 _11472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07508__B _07508_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09969_ _09316_/X _09323_/X _10250_/S vssd1 vssd1 vccd1 vccd1 _09969_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout85_A _12830_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12980_ hold230/X _13004_/A2 _13006_/B1 hold203/X vssd1 vssd1 vccd1 vccd1 hold231/A
+ sky130_fd_sc_hd__a22o_1
X_11931_ _11931_/A _11931_/B _11931_/C vssd1 vssd1 vccd1 vccd1 _11932_/B sky130_fd_sc_hd__and3_1
XANTENNA__08170__A2 fanout69/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11862_ _11862_/A vssd1 vssd1 vccd1 vccd1 _11863_/B sky130_fd_sc_hd__inv_2
XANTENNA__12254__A1 _12254_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10813_ _10813_/A _10813_/B vssd1 vssd1 vccd1 vccd1 _10814_/C sky130_fd_sc_hd__xor2_1
XANTENNA__11057__A2 _12150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11793_ _11793_/A _11793_/B vssd1 vssd1 vccd1 vccd1 _11793_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_67_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08355__A _10949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10744_ _11102_/B _10744_/B vssd1 vssd1 vccd1 vccd1 _10782_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_70_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10675_ _10676_/A _10676_/B vssd1 vssd1 vccd1 vccd1 _10677_/A sky130_fd_sc_hd__and2_1
X_13394_ instruction[10] vssd1 vssd1 vccd1 vccd1 pred_idx[2] sky130_fd_sc_hd__buf_12
X_12414_ _12414_/A _12414_/B _12414_/C vssd1 vssd1 vccd1 vccd1 _12414_/X sky130_fd_sc_hd__or3_1
XFILLER_0_35_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12345_ _12345_/A _12345_/B vssd1 vssd1 vccd1 vccd1 _12362_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_62_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06787__A3 _12644_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12309__A2 _09672_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08630__B1 _08673_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12276_ _12277_/A _12277_/B _12277_/C vssd1 vssd1 vccd1 vccd1 _12276_/X sky130_fd_sc_hd__o21a_1
X_11227_ reg1_val[15] curr_PC[15] vssd1 vssd1 vccd1 vccd1 _11228_/B sky130_fd_sc_hd__nand2_1
XANTENNA__07197__B1 _07200_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07736__A2 _12818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11158_ _11158_/A _11158_/B vssd1 vssd1 vccd1 vccd1 _11160_/B sky130_fd_sc_hd__xor2_1
X_10109_ _10109_/A _10109_/B vssd1 vssd1 vccd1 vccd1 _10109_/Y sky130_fd_sc_hd__nand2_1
X_11089_ _11089_/A _11089_/B vssd1 vssd1 vccd1 vccd1 _11090_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_77_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07320_ _09716_/A _07320_/B vssd1 vssd1 vccd1 vccd1 _07322_/B sky130_fd_sc_hd__xor2_1
XANTENNA__10795__A _10928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07251_ _08584_/A _07251_/B vssd1 vssd1 vccd1 vccd1 _07300_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_6_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07182_ _07200_/A _07182_/B vssd1 vssd1 vccd1 vccd1 _07183_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_5_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10008__B1 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11756__B1 _12316_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09808__B _09808_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09823_ _09106_/X _09129_/X _10248_/S vssd1 vssd1 vccd1 vccd1 _09823_/X sky130_fd_sc_hd__mux2_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06966_ _11020_/A _07074_/A _06967_/C _06967_/D vssd1 vssd1 vccd1 vccd1 _06966_/Y
+ sky130_fd_sc_hd__nor4_2
X_09754_ _11470_/A _09754_/B vssd1 vssd1 vccd1 vccd1 _09755_/B sky130_fd_sc_hd__xnor2_2
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06897_ _06897_/A _06897_/B vssd1 vssd1 vccd1 vccd1 _06902_/B sky130_fd_sc_hd__or2_2
X_09685_ _12388_/S _06810_/X _09684_/X vssd1 vssd1 vccd1 vccd1 _09687_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_69_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08705_ _09010_/A _09010_/B vssd1 vssd1 vccd1 vccd1 _09018_/B sky130_fd_sc_hd__and2_1
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08636_ _08636_/A _08636_/B _08636_/C vssd1 vssd1 vccd1 vccd1 _08652_/A sky130_fd_sc_hd__or3_4
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08567_ _08567_/A _08567_/B vssd1 vssd1 vccd1 vccd1 _08575_/B sky130_fd_sc_hd__xnor2_1
Xfanout11 _07366_/Y vssd1 vssd1 vccd1 vccd1 fanout9/A sky130_fd_sc_hd__buf_4
XFILLER_0_77_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout22 _07087_/X vssd1 vssd1 vccd1 vccd1 _11653_/A sky130_fd_sc_hd__buf_8
XANTENNA__11444__C1 _09172_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07518_ _07519_/A _07519_/B vssd1 vssd1 vccd1 vccd1 _07520_/A sky130_fd_sc_hd__nand2_1
Xfanout55 _07166_/Y vssd1 vssd1 vccd1 vccd1 _12842_/A sky130_fd_sc_hd__clkbuf_8
X_08498_ _08798_/B2 _08744_/A2 _08564_/B _08646_/B2 vssd1 vssd1 vccd1 vccd1 _08499_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_76_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout44 _12840_/A vssd1 vssd1 vccd1 vccd1 _11923_/A sky130_fd_sc_hd__buf_6
Xfanout33 _12261_/A vssd1 vssd1 vccd1 vccd1 _10959_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_37_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout88 _07204_/X vssd1 vssd1 vccd1 vccd1 _10589_/A sky130_fd_sc_hd__buf_6
XFILLER_0_91_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07449_ _07449_/A _07449_/B vssd1 vssd1 vccd1 vccd1 _07456_/A sky130_fd_sc_hd__xnor2_1
Xfanout99 _12816_/A vssd1 vssd1 vccd1 vccd1 fanout99/X sky130_fd_sc_hd__buf_8
Xfanout66 _08752_/B vssd1 vssd1 vccd1 vccd1 fanout66/X sky130_fd_sc_hd__buf_6
Xfanout77 _09548_/A vssd1 vssd1 vccd1 vccd1 _10928_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_36_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11995__B1 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10460_ _10458_/Y _10460_/B vssd1 vssd1 vccd1 vccd1 _10476_/A sky130_fd_sc_hd__nand2b_2
XFILLER_0_17_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_507 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07415__A1 _09444_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09119_ reg1_val[10] reg1_val[21] _09142_/S vssd1 vssd1 vccd1 vccd1 _09119_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_72_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10391_ hold220/A _10391_/A2 _10518_/B _11968_/B1 vssd1 vssd1 vccd1 vccd1 _10391_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__07415__B2 _09236_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12130_ _12124_/Y _12125_/X _12129_/Y _12122_/X vssd1 vssd1 vccd1 vccd1 _12130_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_103_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12061_ _12030_/B _12030_/C _12170_/A vssd1 vssd1 vccd1 vccd1 _12103_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_3_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11012_ _12394_/A _11012_/B vssd1 vssd1 vccd1 vccd1 _11012_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__07179__B1 _10963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12963_ _13214_/A hold249/X vssd1 vssd1 vccd1 vccd1 _13284_/D sky130_fd_sc_hd__and2_1
XFILLER_0_99_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11278__A2 _11989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08143__A2 _08727_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11914_ _11915_/A _11915_/B vssd1 vssd1 vccd1 vccd1 _12012_/A sky130_fd_sc_hd__or2_1
X_12894_ hold269/X hold37/X vssd1 vssd1 vccd1 vccd1 _13139_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__07351__B1 _12830_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11845_ _11846_/A _11846_/B vssd1 vssd1 vccd1 vccd1 _11931_/A sky130_fd_sc_hd__nand2_1
XTAP_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11776_ _11777_/A _11777_/B vssd1 vssd1 vccd1 vccd1 _11861_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_27_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10727_ _10727_/A _10727_/B vssd1 vssd1 vccd1 vccd1 _10729_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_82_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10658_ _10658_/A _10658_/B _10500_/Y _10624_/B vssd1 vssd1 vccd1 vccd1 _11033_/B
+ sky130_fd_sc_hd__or4bb_1
XANTENNA__07406__A1 _12822_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13377_ _13378_/CLK _13377_/D vssd1 vssd1 vccd1 vccd1 hold298/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07406__B2 _12824_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10589_ _10589_/A fanout6/X vssd1 vssd1 vccd1 vccd1 _10590_/B sky130_fd_sc_hd__nor2_1
XANTENNA__07429__A _10710_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12328_ _12328_/A vssd1 vssd1 vccd1 vccd1 _12330_/A sky130_fd_sc_hd__inv_2
XANTENNA__07148__B _09343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12259_ _11673_/A _12210_/B _12211_/X vssd1 vssd1 vccd1 vccd1 _12263_/A sky130_fd_sc_hd__a21o_1
XANTENNA__07709__A2 _07087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06820_ _10879_/A _06819_/X _06728_/Y vssd1 vssd1 vccd1 vccd1 _06820_/X sky130_fd_sc_hd__o21a_1
XANTENNA__07164__A _09445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06751_ reg2_val[8] _06799_/B vssd1 vssd1 vccd1 vccd1 _06751_/X sky130_fd_sc_hd__and2_1
XFILLER_0_116_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06682_ reg1_val[19] _07210_/A vssd1 vssd1 vccd1 vccd1 _06683_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_92_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09470_ _09260_/A _09260_/C _09260_/B vssd1 vssd1 vccd1 vccd1 _09473_/A sky130_fd_sc_hd__o21bai_4
XFILLER_0_116_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08421_ _08421_/A _08421_/B vssd1 vssd1 vccd1 vccd1 _08454_/A sky130_fd_sc_hd__or2_1
XFILLER_0_58_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06625__A_N _07343_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08352_ _07955_/A _08744_/A2 _08564_/B _07896_/A vssd1 vssd1 vccd1 vccd1 _08353_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_18_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07303_ _08000_/A _07303_/B vssd1 vssd1 vccd1 vccd1 _07628_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_73_254 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08283_ _08291_/A _08291_/B vssd1 vssd1 vccd1 vccd1 _08283_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_73_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07234_ _07270_/A _07270_/B vssd1 vssd1 vccd1 vccd1 _07234_/X sky130_fd_sc_hd__or2_1
XANTENNA_fanout135_A _12814_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_82 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout302_A _06578_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07165_ _09441_/A _09758_/A _07163_/X vssd1 vssd1 vccd1 vccd1 _07165_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_42_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07096_ reg1_val[18] _07096_/B vssd1 vssd1 vccd1 vccd1 _11470_/B sky130_fd_sc_hd__xnor2_4
Xfanout223 _06890_/Y vssd1 vssd1 vccd1 vccd1 _12789_/B sky130_fd_sc_hd__clkbuf_8
Xfanout201 _12830_/B vssd1 vssd1 vccd1 vccd1 _12818_/B sky130_fd_sc_hd__buf_4
XFILLER_0_100_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout212 _09445_/A vssd1 vssd1 vccd1 vccd1 _08728_/A sky130_fd_sc_hd__buf_12
XFILLER_0_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout234 _06794_/X vssd1 vssd1 vccd1 vccd1 _10248_/S sky130_fd_sc_hd__clkbuf_4
Xfanout245 _06596_/Y vssd1 vssd1 vccd1 vccd1 _06703_/B1 sky130_fd_sc_hd__buf_4
Xfanout256 _08436_/B vssd1 vssd1 vccd1 vccd1 _08038_/A sky130_fd_sc_hd__clkbuf_8
Xfanout278 _13246_/B2 vssd1 vssd1 vccd1 vccd1 _06572_/A sky130_fd_sc_hd__buf_4
Xfanout289 _06771_/A vssd1 vssd1 vccd1 vccd1 _06720_/B sky130_fd_sc_hd__buf_4
Xfanout267 _06881_/X vssd1 vssd1 vccd1 vccd1 _11142_/S sky130_fd_sc_hd__clkbuf_16
X_09806_ _09808_/A _09808_/B vssd1 vssd1 vccd1 vccd1 _09806_/X sky130_fd_sc_hd__or2_1
X_07998_ _07770_/A _07770_/B _07769_/A vssd1 vssd1 vccd1 vccd1 _08004_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__07074__A _07074_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06949_ _10710_/A vssd1 vssd1 vccd1 vccd1 _10444_/A sky130_fd_sc_hd__inv_6
X_09737_ _10448_/A _09737_/B vssd1 vssd1 vccd1 vccd1 _09741_/A sky130_fd_sc_hd__xnor2_1
X_09668_ _09666_/X _09667_/X _09974_/A vssd1 vssd1 vccd1 vccd1 _09668_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_96_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout48_A _12838_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09873__A2 _11751_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09599_ _09446_/A _09446_/B _09442_/Y vssd1 vssd1 vccd1 vccd1 _09603_/A sky130_fd_sc_hd__a21oi_2
X_08619_ _08733_/A _08619_/B vssd1 vssd1 vccd1 vccd1 _08628_/B sky130_fd_sc_hd__xnor2_2
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11630_ _12244_/S _11630_/B vssd1 vssd1 vccd1 vccd1 _11630_/X sky130_fd_sc_hd__or2_1
XANTENNA__09086__A0 _12626_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08617__B _08617_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11561_ _11570_/A vssd1 vssd1 vccd1 vccd1 _11561_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_21_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12139__B _12412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13300_ _13307_/CLK hold176/X vssd1 vssd1 vccd1 vccd1 _13300_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_119_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10512_ _10510_/Y _10512_/B vssd1 vssd1 vccd1 vccd1 _10513_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_92_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_438 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11492_ _11371_/A _11371_/B _11370_/A vssd1 vssd1 vccd1 vccd1 _11497_/A sky130_fd_sc_hd__a21o_1
X_13231_ hold250/X _12789_/B _13230_/X _12790_/A vssd1 vssd1 vccd1 vccd1 hold251/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10443_ _10589_/A fanout13/X fanout6/X _07208_/Y vssd1 vssd1 vccd1 vccd1 _10444_/B
+ sky130_fd_sc_hd__o22a_1
X_13162_ hold271/X _06890_/Y _13161_/X _13246_/B2 vssd1 vssd1 vccd1 vccd1 hold272/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10374_ _09653_/A _08996_/A _08996_/B vssd1 vssd1 vccd1 vccd1 _10374_/Y sky130_fd_sc_hd__a21oi_1
X_12113_ reg1_val[25] curr_PC[25] vssd1 vssd1 vccd1 vccd1 _12113_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_20_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13093_ hold260/A _13092_/X fanout1/X vssd1 vssd1 vccd1 vccd1 _13093_/X sky130_fd_sc_hd__mux2_1
X_12044_ _12434_/B1 _12123_/B hold218/A vssd1 vssd1 vccd1 vccd1 _12044_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__11218__B _11650_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08116__A2 _07896_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12946_ hold265/A hold19/X vssd1 vssd1 vccd1 vccd1 _12947_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_99_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12877_ hold15/X hold293/A vssd1 vssd1 vccd1 vccd1 _12877_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_87_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11234__A _11886_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11828_ fanout29/X _12213_/A fanout56/X fanout27/X vssd1 vssd1 vccd1 vccd1 _11829_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_28_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11759_ _09613_/A fanout12/X fanout8/X _09614_/A vssd1 vssd1 vccd1 vccd1 _11760_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_70_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08970_ _08971_/A _08971_/B vssd1 vssd1 vccd1 vccd1 _09075_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_53_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07921_ _08740_/A _07921_/B vssd1 vssd1 vccd1 vccd1 _07923_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__11895__C1 _12307_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07852_ _07807_/B _07848_/X _07849_/Y _07824_/X vssd1 vssd1 vccd1 vccd1 _07854_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_127_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12439__A1 _09108_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06803_ _09343_/A _09666_/S vssd1 vssd1 vccd1 vccd1 _09523_/A sky130_fd_sc_hd__or2_1
XANTENNA__10162__A2 _07154_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09522_ _09343_/A _09505_/S _09351_/B _12626_/A vssd1 vssd1 vccd1 vccd1 _09523_/B
+ sky130_fd_sc_hd__a22o_1
X_07783_ _07783_/A _07783_/B vssd1 vssd1 vccd1 vccd1 _07784_/B sky130_fd_sc_hd__xnor2_1
X_06734_ _06963_/A reg1_val[11] vssd1 vssd1 vccd1 vccd1 _06734_/X sky130_fd_sc_hd__and2b_1
XANTENNA__09313__S _09666_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06665_ reg2_val[20] _06771_/A _06703_/B1 _06664_/Y vssd1 vssd1 vccd1 vccd1 _07223_/A
+ sky130_fd_sc_hd__o2bb2a_2
X_09453_ _09453_/A _09453_/B vssd1 vssd1 vccd1 vccd1 _09456_/A sky130_fd_sc_hd__nand2_1
X_09384_ _09385_/A _09385_/B vssd1 vssd1 vccd1 vccd1 _09386_/A sky130_fd_sc_hd__or2_1
XFILLER_0_59_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08404_ _08722_/A _08404_/B vssd1 vssd1 vccd1 vccd1 _08434_/A sky130_fd_sc_hd__xnor2_1
X_06596_ _06596_/A _06596_/B vssd1 vssd1 vccd1 vccd1 _06596_/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_52_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08335_ _08335_/A _08335_/B vssd1 vssd1 vccd1 vccd1 _08347_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_117_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08266_ _08266_/A _08266_/B vssd1 vssd1 vccd1 vccd1 _08329_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_6_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13167__A2 _12789_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07217_ _10165_/A _07217_/B vssd1 vssd1 vccd1 vccd1 _10320_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_61_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09268__B _10567_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08197_ _08197_/A _08197_/B vssd1 vssd1 vccd1 vccd1 _08245_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_104_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07148_ _07149_/A _09343_/A vssd1 vssd1 vccd1 vccd1 _08632_/C sky130_fd_sc_hd__and2_1
XFILLER_0_15_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08043__A1 _08727_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09240__B1 _09441_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08043__B2 _08727_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07079_ _07036_/A _06960_/C _09147_/S _06964_/A _07074_/B vssd1 vssd1 vccd1 vccd1
+ _07080_/B sky130_fd_sc_hd__o41a_2
X_10090_ _10090_/A _10090_/B vssd1 vssd1 vccd1 vccd1 _10092_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_10_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12800_ hold88/X _12818_/B vssd1 vssd1 vccd1 vccd1 hold89/A sky130_fd_sc_hd__or2_1
X_10992_ _10992_/A _11215_/A vssd1 vssd1 vccd1 vccd1 _10992_/X sky130_fd_sc_hd__or2_1
XFILLER_0_69_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07532__A _11065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07857__A1 _10927_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07857__B2 _11367_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12731_ reg1_val[21] _12741_/B vssd1 vssd1 vccd1 vccd1 _12732_/B sky130_fd_sc_hd__nand2_2
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12662_ _12661_/A _12658_/Y _12660_/B vssd1 vssd1 vccd1 vccd1 _12666_/A sky130_fd_sc_hd__o21a_2
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11613_ _11785_/A _11613_/B vssd1 vssd1 vccd1 vccd1 _11649_/D sky130_fd_sc_hd__xor2_1
XANTENNA__11989__A _11989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12593_ _12591_/X _12593_/B vssd1 vssd1 vccd1 vccd1 _12605_/B sky130_fd_sc_hd__nand2b_2
XFILLER_0_92_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11810__C1 _12247_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11544_ _13300_/Q _11544_/B vssd1 vssd1 vccd1 vccd1 _11632_/B sky130_fd_sc_hd__or2_1
XFILLER_0_108_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07085__A2 _07090_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11475_ _11475_/A _11475_/B _11475_/C vssd1 vssd1 vccd1 vccd1 _11476_/B sky130_fd_sc_hd__or3_1
XFILLER_0_123_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13214_ _13214_/A _13214_/B vssd1 vssd1 vccd1 vccd1 _13373_/D sky130_fd_sc_hd__and2_1
X_10426_ _10574_/A _11472_/A _10574_/B _10575_/A vssd1 vssd1 vccd1 vccd1 _10427_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_0_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13145_ _13145_/A _13145_/B vssd1 vssd1 vccd1 vccd1 _13145_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_103_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10357_ _10358_/A _10358_/B vssd1 vssd1 vccd1 vccd1 _10412_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_21_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13076_ hold67/X _12791_/A _13080_/B1 _13341_/Q _13113_/A vssd1 vssd1 vccd1 vccd1
+ hold68/A sky130_fd_sc_hd__o221a_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10288_ _10288_/A _10288_/B vssd1 vssd1 vccd1 vccd1 _10290_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__09534__A1 _12394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12027_ _11323_/B _11702_/Y _12025_/Y _12026_/X _12023_/X vssd1 vssd1 vccd1 vccd1
+ _12028_/B sky130_fd_sc_hd__a311oi_4
XANTENNA__10144__A2 _10797_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13094__B2 _06572_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12929_ _13144_/B _13145_/A _12891_/X vssd1 vssd1 vccd1 vccd1 _13150_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_88_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06984__C _06986_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08273__A1 _08721_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08273__B2 _08739_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08120_ _08120_/A _08120_/B vssd1 vssd1 vccd1 vccd1 _08121_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_114_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08051_ _08741_/B2 _08741_/A2 _08617_/B _08732_/A1 vssd1 vssd1 vccd1 vccd1 _08052_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_114_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07002_ reg1_val[27] _07002_/B vssd1 vssd1 vccd1 vccd1 _07522_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_3_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10027__B _10027_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08953_ _08954_/A _08954_/B vssd1 vssd1 vccd1 vccd1 _09072_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07904_ _07903_/A _07972_/A vssd1 vssd1 vccd1 vccd1 _07966_/A sky130_fd_sc_hd__nand2b_1
X_08884_ _08885_/B _08885_/A vssd1 vssd1 vccd1 vccd1 _08884_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_98_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07835_ _07835_/A _07835_/B vssd1 vssd1 vccd1 vccd1 _07836_/B sky130_fd_sc_hd__xor2_1
XANTENNA__13085__A1 _07508_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07766_ _08724_/A _07766_/B vssd1 vssd1 vccd1 vccd1 _07768_/B sky130_fd_sc_hd__xnor2_1
X_06717_ reg1_val[14] _06981_/A vssd1 vssd1 vccd1 vccd1 _11130_/S sky130_fd_sc_hd__and2_1
X_09505_ _09118_/X _09143_/X _09505_/S vssd1 vssd1 vccd1 vccd1 _09505_/X sky130_fd_sc_hd__mux2_1
XANTENNA__07352__A _10707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09436_ _12844_/A _10167_/A1 _10022_/B1 _12846_/A vssd1 vssd1 vccd1 vccd1 _09437_/B
+ sky130_fd_sc_hd__o22a_1
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07697_ _07719_/A vssd1 vssd1 vccd1 vccd1 _07697_/Y sky130_fd_sc_hd__inv_2
X_06648_ _08980_/B _12110_/A _12176_/A _06648_/D vssd1 vssd1 vccd1 vccd1 _06649_/B
+ sky130_fd_sc_hd__and4b_1
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06579_ instruction[0] instruction[1] instruction[2] pred_val vssd1 vssd1 vccd1 vccd1
+ _06581_/B sky130_fd_sc_hd__or4bb_4
X_09367_ _09367_/A vssd1 vssd1 vccd1 vccd1 _09367_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_117_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_50 reg1_val[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09298_ _09298_/A _09298_/B vssd1 vssd1 vccd1 vccd1 _09299_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_62_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08318_ _07885_/B _08741_/A2 _08617_/B _08721_/B1 vssd1 vssd1 vccd1 vccd1 _08319_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08183__A _08745_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_61 instruction[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10071__A1 _11146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10071__B2 _11294_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08249_ _08249_/A _08249_/B vssd1 vssd1 vccd1 vccd1 _08254_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11260_ _11653_/A _12213_/A fanout56/X _08752_/B vssd1 vssd1 vccd1 vccd1 _11261_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_113_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07224__C1 _07135_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10211_ _10211_/A _10211_/B _10211_/C vssd1 vssd1 vccd1 vccd1 _10212_/B sky130_fd_sc_hd__or3_1
X_11191_ _11191_/A _11191_/B vssd1 vssd1 vccd1 vccd1 _11205_/A sky130_fd_sc_hd__xnor2_1
X_10142_ _10093_/A _10093_/B _10091_/X vssd1 vssd1 vccd1 vccd1 _10231_/A sky130_fd_sc_hd__a21oi_4
XFILLER_0_30_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11571__B2 _11923_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11571__A1 _11847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10073_ _10073_/A _10073_/B vssd1 vssd1 vccd1 vccd1 _10076_/C sky130_fd_sc_hd__xnor2_2
XFILLER_0_27_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10888__A _11886_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12714_ reg1_val[17] _12741_/B vssd1 vssd1 vccd1 vccd1 _12725_/B sky130_fd_sc_hd__xnor2_4
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10975_ _10976_/A _10976_/B _10976_/C vssd1 vssd1 vccd1 vccd1 _11088_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_85_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12645_ _12643_/Y _12645_/B vssd1 vssd1 vccd1 vccd1 _12646_/B sky130_fd_sc_hd__and2b_1
XANTENNA__13203__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12576_ _12581_/C _12576_/B vssd1 vssd1 vccd1 vccd1 new_PC[19] sky130_fd_sc_hd__xnor2_4
XANTENNA__12051__A2 _12404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11527_ _11524_/X _11526_/Y _06693_/X vssd1 vssd1 vccd1 vccd1 _11527_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_80_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11458_ _11430_/Y _11433_/Y _11457_/X _11359_/Y vssd1 vssd1 vccd1 vccd1 dest_val[17]
+ sky130_fd_sc_hd__o31a_4
XFILLER_0_40_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09917__A _10959_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10409_ _10656_/B _10409_/B vssd1 vssd1 vccd1 vccd1 _10409_/X sky130_fd_sc_hd__and2_1
X_11389_ _11389_/A _11389_/B vssd1 vssd1 vccd1 vccd1 _11390_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_0_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13128_ _13128_/A hold274/X vssd1 vssd1 vccd1 vccd1 _13355_/D sky130_fd_sc_hd__and2_1
XANTENNA__11562__B2 _09614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11562__A1 _09613_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13059_ _11385_/A _13087_/B2 hold138/X vssd1 vssd1 vccd1 vccd1 hold139/A sky130_fd_sc_hd__o21a_1
XFILLER_0_84_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13067__A1 _10422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07620_ _10448_/A _07620_/B vssd1 vssd1 vccd1 vccd1 _07983_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__08191__B1 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08730__A2 _08038_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07551_ _12264_/B _07551_/B vssd1 vssd1 vccd1 vccd1 _07564_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__08268__A _08728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10310__B _12316_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07482_ _10445_/A _12832_/A _12834_/A _10706_/B2 vssd1 vssd1 vccd1 vccd1 _07483_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07297__A2 _10167_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09221_ _12842_/A _10167_/A1 _10022_/B1 _12844_/A vssd1 vssd1 vccd1 vccd1 _09222_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07900__A _11758_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09152_ _12423_/A _09152_/B vssd1 vssd1 vccd1 vccd1 _09152_/Y sky130_fd_sc_hd__nor2_4
XFILLER_0_90_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09994__A1 _09156_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08103_ _08038_/A _11472_/A _11558_/A _08730_/A1 vssd1 vssd1 vccd1 vccd1 _08104_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_114_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09083_ _12388_/S _09152_/B vssd1 vssd1 vccd1 vccd1 _09083_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__09994__B2 _09111_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout215_A _06939_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10038__A _12076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08034_ _08034_/A _08034_/B _08034_/C vssd1 vssd1 vccd1 vccd1 _08845_/A sky130_fd_sc_hd__or3_1
XANTENNA__08731__A _08731_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07347__A _09442_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07757__B1 _07819_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09985_ _06775_/Y _12403_/A1 _09165_/X _06777_/B _09984_/X vssd1 vssd1 vccd1 vccd1
+ _09985_/X sky130_fd_sc_hd__o221a_1
XANTENNA__06980__A1 _11020_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08936_ _08936_/A _08936_/B vssd1 vssd1 vccd1 vccd1 _08937_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_99_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08867_ _08869_/A _08869_/B vssd1 vssd1 vccd1 vccd1 _08867_/X sky130_fd_sc_hd__or2_1
X_07818_ _07818_/A _07818_/B _07818_/C vssd1 vssd1 vccd1 vccd1 _07840_/A sky130_fd_sc_hd__or3_1
XANTENNA__08721__A2 _07885_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08182__B1 _08564_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08798_ _08752_/A _07087_/A _07087_/B _08752_/B _08798_/B2 vssd1 vssd1 vccd1 vccd1
+ _08799_/B sky130_fd_sc_hd__o32a_1
X_07749_ _08727_/B1 _11847_/A _11766_/A _08727_/A2 vssd1 vssd1 vccd1 vccd1 _07750_/B
+ sky130_fd_sc_hd__o22a_1
X_10760_ _09664_/X _09668_/X _11231_/S vssd1 vssd1 vccd1 vccd1 _10761_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_67_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07288__A2 _11989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09501__S _09666_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09419_ _09420_/A _09420_/B vssd1 vssd1 vccd1 vccd1 _09558_/B sky130_fd_sc_hd__nand2_1
X_10691_ _11172_/A _10691_/B vssd1 vssd1 vccd1 vccd1 _10693_/B sky130_fd_sc_hd__xnor2_1
X_12430_ _12430_/A _12430_/B vssd1 vssd1 vccd1 vccd1 _12430_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_47_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12361_ _12356_/Y _12357_/X _12360_/X _12354_/X vssd1 vssd1 vccd1 vccd1 _12361_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_117_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12292_ _06857_/Y _12291_/X _12388_/S vssd1 vssd1 vccd1 vccd1 _12293_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_62_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09737__A _10448_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11312_ _11313_/A _11313_/B vssd1 vssd1 vccd1 vccd1 _11417_/B sky130_fd_sc_hd__or2_1
X_11243_ _11243_/A _11243_/B vssd1 vssd1 vccd1 vccd1 _11243_/Y sky130_fd_sc_hd__nor2_2
XANTENNA__07257__A _12317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11174_ _07087_/A _07087_/B _12150_/A _12213_/A fanout66/X vssd1 vssd1 vccd1 vccd1
+ _11175_/B sky130_fd_sc_hd__o32a_1
X_10125_ _11452_/B1 _10256_/B hold242/A vssd1 vssd1 vccd1 vccd1 _10125_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_89_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10056_ _10056_/A _10056_/B _10056_/C vssd1 vssd1 vccd1 vccd1 _10057_/B sky130_fd_sc_hd__or3_1
XANTENNA__13049__A1 _06954_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08173__B1 _12820_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07920__B1 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07279__A2 _10567_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10807__B1 fanout27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10958_ _11146_/A _10797_/B fanout5/X _11065_/A vssd1 vssd1 vccd1 vccd1 _10959_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_73_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11480__B1 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10889_ _12244_/S _10883_/A _10888_/X vssd1 vssd1 vccd1 vccd1 _10889_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_72_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08228__A1 _07896_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12628_ reg1_val[1] _12629_/B vssd1 vssd1 vccd1 vccd1 _12630_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_26_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08228__B2 _08723_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12559_ _12623_/A _12559_/B vssd1 vssd1 vccd1 vccd1 _12566_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_53_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_717 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold106 hold106/A vssd1 vssd1 vccd1 vccd1 hold106/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold117 hold117/A vssd1 vssd1 vccd1 vccd1 hold117/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08551__A _09441_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold128 hold128/A vssd1 vssd1 vccd1 vccd1 hold128/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold139 hold139/A vssd1 vssd1 vccd1 vccd1 hold139/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11535__A1 _12394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12073__A _12073_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08400__A1 _07821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08400__B2 _09423_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06982_ reg1_val[14] _06982_/B vssd1 vssd1 vccd1 vccd1 _06986_/B sky130_fd_sc_hd__xnor2_4
X_09770_ _09771_/A _09771_/B vssd1 vssd1 vccd1 vccd1 _09770_/X sky130_fd_sc_hd__and2b_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08721_ _10537_/A1 _07885_/B _08721_/B1 _08432_/B vssd1 vssd1 vccd1 vccd1 _08722_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08652_ _08652_/A _08652_/B vssd1 vssd1 vccd1 vccd1 _08653_/B sky130_fd_sc_hd__xor2_2
X_07603_ _07603_/A _07603_/B vssd1 vssd1 vccd1 vccd1 _07604_/B sky130_fd_sc_hd__nand2_1
XANTENNA_fanout165_A _08979_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08583_ _08612_/A _08612_/B vssd1 vssd1 vccd1 vccd1 _08613_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_49_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07534_ _07533_/B _07533_/C _09746_/A vssd1 vssd1 vccd1 vccd1 _07540_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_48_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07465_ _07568_/A _07568_/B vssd1 vssd1 vccd1 vccd1 _07569_/A sky130_fd_sc_hd__and2_1
XFILLER_0_48_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09204_ _09205_/A _09205_/B _09205_/C vssd1 vssd1 vccd1 vccd1 _09469_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_8_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07396_ _07396_/A _07396_/B vssd1 vssd1 vccd1 vccd1 _07399_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09135_ reg1_val[3] reg1_val[28] _09142_/S vssd1 vssd1 vccd1 vccd1 _09135_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_8_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07442__A2 _12808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08461__A _09441_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09066_ _09066_/A _09066_/B vssd1 vssd1 vccd1 vccd1 _09067_/B sky130_fd_sc_hd__nand2_1
X_08017_ _08017_/A _08017_/B vssd1 vssd1 vccd1 vccd1 _08019_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_4_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10329__A2 _10574_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07508__C _10959_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09968_ _09968_/A vssd1 vssd1 vccd1 vccd1 _09968_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_99_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08919_ _08919_/A _08919_/B vssd1 vssd1 vccd1 vccd1 _08920_/B sky130_fd_sc_hd__xnor2_2
X_09899_ _09900_/A _09900_/B vssd1 vssd1 vccd1 vccd1 _09899_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__08155__B1 _07955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11930_ _11931_/A _11931_/B _11931_/C vssd1 vssd1 vccd1 vccd1 _11932_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_99_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10231__A _10231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11861_ _11861_/A _11861_/B _11861_/C vssd1 vssd1 vccd1 vccd1 _11862_/A sky130_fd_sc_hd__and3_1
XANTENNA__12254__A2 _09821_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06681__A_N _07210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11792_ _11792_/A _11792_/B vssd1 vssd1 vccd1 vccd1 _11793_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_39_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10812_ _11172_/A _10812_/B vssd1 vssd1 vccd1 vccd1 _10813_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_67_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10743_ _09652_/B _10232_/X _10741_/X _10742_/X _10740_/X vssd1 vssd1 vccd1 vccd1
+ _10744_/B sky130_fd_sc_hd__o311a_2
XFILLER_0_55_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11462__B1 fanout12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10377__S _12388_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10674_ _11261_/A _10674_/B vssd1 vssd1 vccd1 vccd1 _10676_/B sky130_fd_sc_hd__xnor2_1
X_13393_ instruction[9] vssd1 vssd1 vccd1 vccd1 pred_idx[1] sky130_fd_sc_hd__buf_12
XFILLER_0_106_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12413_ _12413_/A _12413_/B vssd1 vssd1 vccd1 vccd1 _12414_/C sky130_fd_sc_hd__nand2_1
XANTENNA__12962__B1 _13213_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12344_ _06647_/B _12341_/X _12342_/Y _11624_/A vssd1 vssd1 vccd1 vccd1 _12345_/B
+ sky130_fd_sc_hd__a31o_1
XANTENNA__08630__A1 _08646_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08630__B2 _07752_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06603__B _07144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12275_ _12275_/A _12275_/B vssd1 vssd1 vccd1 vccd1 _12277_/C sky130_fd_sc_hd__xnor2_1
X_11226_ reg1_val[15] curr_PC[15] vssd1 vssd1 vccd1 vccd1 _11226_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_4_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11157_ _12210_/A _11157_/B vssd1 vssd1 vccd1 vccd1 _11158_/B sky130_fd_sc_hd__xnor2_1
X_10108_ _06813_/Y _10107_/Y _12388_/S vssd1 vssd1 vccd1 vccd1 _10109_/B sky130_fd_sc_hd__mux2_1
XANTENNA__07715__A _07833_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11088_ _11088_/A _11088_/B _11088_/C vssd1 vssd1 vccd1 vccd1 _11089_/B sky130_fd_sc_hd__and3_1
X_10039_ _10040_/A _10040_/B _10040_/C vssd1 vssd1 vccd1 vccd1 _10042_/B sky130_fd_sc_hd__and3_1
XFILLER_0_86_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11453__B1 _09167_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09141__S _09142_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07250_ _12832_/A _10167_/A1 _12834_/A _10022_/B1 vssd1 vssd1 vccd1 vccd1 _07251_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_53_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07181_ _07603_/A _07603_/B vssd1 vssd1 vccd1 vccd1 _07604_/A sky130_fd_sc_hd__or2_1
XFILLER_0_41_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10008__B2 _10445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10008__A1 _06971_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11756__A1 fanout24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11756__B2 _07819_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09822_ _09098_/X _09113_/X _10250_/S vssd1 vssd1 vccd1 vccd1 _09824_/B sky130_fd_sc_hd__mux2_1
X_09753_ _10941_/A _11558_/A _11751_/A fanout94/X vssd1 vssd1 vccd1 vccd1 _09754_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06965_ _06988_/A _06981_/A vssd1 vssd1 vccd1 vccd1 _06967_/D sky130_fd_sc_hd__or2_1
X_08704_ _09002_/A _08699_/A _08699_/B _09006_/A _08702_/Y vssd1 vssd1 vccd1 vccd1
+ _09008_/B sky130_fd_sc_hd__a41o_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09684_ _12341_/A _09684_/B _09684_/C vssd1 vssd1 vccd1 vccd1 _09684_/X sky130_fd_sc_hd__or3_1
X_06896_ instruction[13] _06896_/B vssd1 vssd1 vccd1 vccd1 dest_pred[2] sky130_fd_sc_hd__and2_4
XFILLER_0_96_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08635_ _09442_/A _08635_/B _08635_/C vssd1 vssd1 vccd1 vccd1 _08636_/C sky130_fd_sc_hd__and3_1
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08566_ _08591_/A _08591_/B vssd1 vssd1 vccd1 vccd1 _08575_/A sky130_fd_sc_hd__and2b_1
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07517_ _07517_/A _07517_/B vssd1 vssd1 vccd1 vccd1 _07519_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_76_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout12 _12854_/A vssd1 vssd1 vccd1 vccd1 fanout12/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_37_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08497_ _09441_/A _08497_/B vssd1 vssd1 vccd1 vccd1 _08501_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_64_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout45 _12840_/A vssd1 vssd1 vccd1 vccd1 _10570_/B sky130_fd_sc_hd__buf_4
Xfanout56 _10941_/B vssd1 vssd1 vccd1 vccd1 fanout56/X sky130_fd_sc_hd__buf_6
Xfanout34 _12264_/B vssd1 vssd1 vccd1 vccd1 _12261_/A sky130_fd_sc_hd__buf_8
Xfanout23 fanout24/X vssd1 vssd1 vccd1 vccd1 fanout23/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__11995__A1 _12213_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07448_ _11673_/A _07448_/B vssd1 vssd1 vccd1 vccd1 _07449_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_52_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout67 _07090_/Y vssd1 vssd1 vccd1 vccd1 _08752_/B sky130_fd_sc_hd__buf_6
Xfanout89 _07178_/Y vssd1 vssd1 vccd1 vccd1 _10963_/A sky130_fd_sc_hd__clkbuf_8
Xfanout78 _07256_/Y vssd1 vssd1 vccd1 vccd1 _09548_/A sky130_fd_sc_hd__buf_8
XFILLER_0_9_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11995__B2 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07379_ _07579_/B _07377_/B _07395_/B _07378_/B _07378_/A vssd1 vssd1 vccd1 vccd1
+ _07393_/A sky130_fd_sc_hd__o32a_1
XFILLER_0_122_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09118_ _09116_/X _09117_/X _09330_/S vssd1 vssd1 vccd1 vccd1 _09118_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_45_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10390_ _10391_/A2 _10518_/B hold220/A vssd1 vssd1 vccd1 vccd1 _10390_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__07415__A2 _10941_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09049_ _09049_/A _09049_/B vssd1 vssd1 vccd1 vccd1 _09049_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_20_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12060_ _12455_/S _12056_/X _12057_/X _12059_/Y vssd1 vssd1 vccd1 vccd1 dest_val[24]
+ sky130_fd_sc_hd__a22o_4
XANTENNA__07179__A1 _08741_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11011_ _09496_/Y _11010_/X _11233_/S vssd1 vssd1 vccd1 vccd1 _11012_/B sky130_fd_sc_hd__mux2_2
XANTENNA__07179__B2 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10183__B1 _10570_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12962_ hold290/A _13213_/B2 _13213_/A2 hold248/X vssd1 vssd1 vccd1 vccd1 hold249/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08679__A1 _12626_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08679__B2 _09351_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12893_ hold37/X hold269/X vssd1 vssd1 vccd1 vccd1 _12893_/X sky130_fd_sc_hd__and2b_1
X_11913_ _11992_/B _11913_/B vssd1 vssd1 vccd1 vccd1 _11915_/B sky130_fd_sc_hd__or2_1
XFILLER_0_68_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07351__A1 _10445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07351__B2 _10706_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11844_ _12261_/A _11844_/B vssd1 vssd1 vccd1 vccd1 _11846_/B sky130_fd_sc_hd__xnor2_1
XTAP_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08366__A _10949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11775_ _11775_/A _11775_/B vssd1 vssd1 vccd1 vccd1 _11777_/B sky130_fd_sc_hd__xnor2_1
XTAP_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10726_ _10727_/B _10727_/A vssd1 vssd1 vccd1 vccd1 _10854_/A sky130_fd_sc_hd__and2b_1
X_10657_ _10655_/X _10656_/Y _11142_/S vssd1 vssd1 vccd1 vccd1 dest_val[10] sky130_fd_sc_hd__mux2_8
XFILLER_0_82_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09197__A _09716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13376_ _13376_/CLK _13376_/D vssd1 vssd1 vccd1 vccd1 hold268/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07406__A2 _10941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10588_ _10425_/B _10428_/B _10423_/Y vssd1 vssd1 vccd1 vccd1 _10592_/A sky130_fd_sc_hd__a21o_1
X_12327_ _12327_/A _12327_/B _12327_/C vssd1 vssd1 vccd1 vccd1 _12328_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_11_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12258_ _06882_/Y _12204_/X _12232_/Y _12257_/X vssd1 vssd1 vccd1 vccd1 dest_val[27]
+ sky130_fd_sc_hd__o22a_4
XANTENNA__07709__A3 _07087_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11209_ _11210_/A _11210_/B _11210_/C vssd1 vssd1 vccd1 vccd1 _11209_/X sky130_fd_sc_hd__a21o_1
X_12189_ hold281/A _11636_/B _12245_/B _12247_/C1 vssd1 vssd1 vccd1 vccd1 _12190_/B
+ sky130_fd_sc_hd__a31o_1
X_06750_ _06750_/A _06750_/B vssd1 vssd1 vccd1 vccd1 _10507_/A sky130_fd_sc_hd__or2_1
X_06681_ _07210_/A reg1_val[19] vssd1 vssd1 vccd1 vccd1 _11638_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_116_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09882__A3 _12264_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08420_ _08429_/A _08429_/B vssd1 vssd1 vccd1 vccd1 _08421_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_116_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07180__A _11163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08351_ _08742_/A _08351_/B vssd1 vssd1 vccd1 vccd1 _08413_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07302_ _07302_/A _07302_/B vssd1 vssd1 vccd1 vccd1 _07628_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_41_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08282_ _08282_/A _08282_/B vssd1 vssd1 vccd1 vccd1 _08291_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_18_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07233_ _07233_/A _07233_/B vssd1 vssd1 vccd1 vccd1 _07270_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__13121__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12526__A _12686_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11729__A1 _07223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout128_A _07222_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07164_ _09445_/A _07164_/B vssd1 vssd1 vccd1 vccd1 _09758_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_26_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07095_ _07095_/A _07095_/B vssd1 vssd1 vccd1 vccd1 _12812_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout202 _12830_/B vssd1 vssd1 vccd1 vccd1 _12798_/B sky130_fd_sc_hd__buf_4
XFILLER_0_100_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout213 _07120_/Y vssd1 vssd1 vccd1 vccd1 _09445_/A sky130_fd_sc_hd__buf_12
XANTENNA__08358__B1 _12820_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout246 _09355_/X vssd1 vssd1 vccd1 vccd1 _11636_/B sky130_fd_sc_hd__buf_4
Xfanout235 _09503_/S vssd1 vssd1 vccd1 vccd1 _09974_/A sky130_fd_sc_hd__clkbuf_8
Xfanout224 _09311_/S vssd1 vssd1 vccd1 vccd1 _09351_/B sky130_fd_sc_hd__clkbuf_8
XANTENNA__12261__A _12261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout279 _12790_/A vssd1 vssd1 vccd1 vccd1 _13246_/B2 sky130_fd_sc_hd__clkbuf_4
Xfanout268 _06770_/X vssd1 vssd1 vccd1 vccd1 _12244_/S sky130_fd_sc_hd__clkbuf_8
Xfanout257 _07149_/Y vssd1 vssd1 vccd1 vccd1 _08436_/B sky130_fd_sc_hd__clkbuf_8
X_09805_ _09805_/A _09805_/B vssd1 vssd1 vccd1 vccd1 _09808_/B sky130_fd_sc_hd__xnor2_4
X_07997_ _07997_/A _07997_/B vssd1 vssd1 vccd1 vccd1 _08006_/A sky130_fd_sc_hd__xnor2_1
X_06948_ reg1_val[11] _06948_/B vssd1 vssd1 vccd1 vccd1 _09431_/A sky130_fd_sc_hd__xnor2_4
X_09736_ _10706_/B2 _10571_/B _11923_/A _10445_/A vssd1 vssd1 vccd1 vccd1 _09737_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09858__B1 _10575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09667_ _09327_/X _09329_/X _09669_/S vssd1 vssd1 vccd1 vccd1 _09667_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09570__A _10165_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11665__B1 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06879_ _06926_/A _06862_/Y _06877_/X vssd1 vssd1 vccd1 vccd1 _06880_/B sky130_fd_sc_hd__o21a_1
X_08618_ _08671_/B2 _09238_/B _09440_/B1 _08646_/B2 vssd1 vssd1 vccd1 vccd1 _08619_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_69_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09598_ _09598_/A _12264_/B vssd1 vssd1 vccd1 vccd1 _09604_/A sky130_fd_sc_hd__nand2_1
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08186__A _08742_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08549_ _08549_/A _08549_/B vssd1 vssd1 vccd1 vccd1 _08572_/A sky130_fd_sc_hd__xnor2_1
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11560_ _11682_/B _11560_/B vssd1 vssd1 vccd1 vccd1 _11570_/A sky130_fd_sc_hd__and2_1
XFILLER_0_107_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10640__A1 _12244_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10511_ reg1_val[9] curr_PC[9] vssd1 vssd1 vccd1 vccd1 _10512_/B sky130_fd_sc_hd__nand2_1
XANTENNA_fanout7_A fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13230_ hold268/A _13229_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13230_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_45_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11491_ _11405_/A _11405_/B _11403_/Y vssd1 vssd1 vccd1 vccd1 _11499_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10442_ _10288_/A _10288_/B _10285_/A vssd1 vssd1 vccd1 vccd1 _10455_/A sky130_fd_sc_hd__a21o_1
X_13161_ hold279/A _13160_/Y fanout2/A vssd1 vssd1 vccd1 vccd1 _13161_/X sky130_fd_sc_hd__mux2_1
XANTENNA__08597__B1 _08673_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10373_ _11874_/A _10410_/A _10658_/B vssd1 vssd1 vccd1 vccd1 _10373_/X sky130_fd_sc_hd__and3_1
XFILLER_0_32_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13092_ _13092_/A _13092_/B vssd1 vssd1 vccd1 vccd1 _13092_/X sky130_fd_sc_hd__xor2_1
X_12112_ _12041_/A _12038_/Y _12040_/B vssd1 vssd1 vccd1 vccd1 _12112_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_60_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12043_ hold192/A _12043_/B vssd1 vssd1 vccd1 vccd1 _12123_/B sky130_fd_sc_hd__or2_1
XANTENNA__10156__B1 _10963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07265__A _12138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09849__B1 _06881_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12853__C1 _13128_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12945_ _13197_/B _13198_/A _12872_/X vssd1 vssd1 vccd1 vccd1 _13202_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_87_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12876_ hold275/A hold9/X vssd1 vssd1 vccd1 vccd1 _13188_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__07204__S _10444_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11234__B _11234_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11827_ _12317_/A _11827_/B vssd1 vssd1 vccd1 vccd1 _11831_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_28_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11758_ _11758_/A _11758_/B vssd1 vssd1 vccd1 vccd1 _11762_/B sky130_fd_sc_hd__xnor2_1
X_10709_ _11163_/A _10709_/B vssd1 vssd1 vccd1 vccd1 _10710_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_16_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_55 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11689_ _11689_/A _11689_/B vssd1 vssd1 vccd1 vccd1 _11691_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_11_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13359_ _13365_/CLK _13359_/D vssd1 vssd1 vccd1 vccd1 hold287/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09655__A _11707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07920_ fanout99/X fanout87/X fanout82/X _12818_/A vssd1 vssd1 vccd1 vccd1 _07921_/B
+ sky130_fd_sc_hd__o22a_1
X_07851_ _07824_/X _07849_/Y _07848_/X _07807_/B vssd1 vssd1 vccd1 vccd1 _07854_/A
+ sky130_fd_sc_hd__o211ai_1
X_06802_ _09343_/A _09663_/S vssd1 vssd1 vccd1 vccd1 _06802_/X sky130_fd_sc_hd__and2_1
X_07782_ _07782_/A _07782_/B vssd1 vssd1 vccd1 vccd1 _07783_/B sky130_fd_sc_hd__nor2_1
X_09521_ hold238/A _10391_/A2 _09519_/X _12401_/B1 vssd1 vssd1 vccd1 vccd1 _09521_/X
+ sky130_fd_sc_hd__a31o_1
X_06733_ _06805_/A _06702_/A _12686_/B _06732_/X vssd1 vssd1 vccd1 vccd1 _06963_/A
+ sky130_fd_sc_hd__a31o_4
XANTENNA__13116__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06664_ _06686_/A _12649_/B vssd1 vssd1 vccd1 vccd1 _06664_/Y sky130_fd_sc_hd__nor2_1
X_09452_ _09452_/A _09452_/B vssd1 vssd1 vccd1 vccd1 _09453_/B sky130_fd_sc_hd__nand2_1
X_06595_ instruction[24] _06587_/X _06897_/B instruction[41] _06591_/X vssd1 vssd1
+ vccd1 vccd1 _06596_/B sky130_fd_sc_hd__a221o_1
X_09383_ _09716_/A _09383_/B vssd1 vssd1 vccd1 vccd1 _09385_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_59_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08403_ _08673_/A _10537_/A1 _08432_/B _08798_/B2 vssd1 vssd1 vccd1 vccd1 _08404_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_52_60 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08334_ _08331_/A _08331_/B _08384_/A vssd1 vssd1 vccd1 vccd1 _08347_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_19_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08265_ _08266_/A _08266_/B vssd1 vssd1 vccd1 vccd1 _08265_/X sky130_fd_sc_hd__or2_1
XFILLER_0_27_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07216_ _10165_/A _07217_/B vssd1 vssd1 vccd1 vccd1 _10321_/A sky130_fd_sc_hd__or2_1
XFILLER_0_61_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08196_ _08722_/A _08196_/B vssd1 vssd1 vccd1 vccd1 _08245_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__08579__B1 _08673_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07147_ _09594_/A _07147_/B vssd1 vssd1 vccd1 vccd1 _07174_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_30_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08043__A2 _11472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12127__A1 _12307_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07078_ _11470_/A _07078_/B vssd1 vssd1 vccd1 vccd1 _07093_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__12703__B _12703_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11350__A2 _11234_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12835__C1 _13214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09719_ _09719_/A _09719_/B vssd1 vssd1 vccd1 vccd1 _09722_/A sky130_fd_sc_hd__nand2_4
X_10991_ _10738_/X _11215_/A _10989_/Y vssd1 vssd1 vccd1 vccd1 _11424_/A sky130_fd_sc_hd__o21ba_1
Xclkbuf_4_6_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13311_/CLK sky130_fd_sc_hd__clkbuf_8
XANTENNA__07532__B _10571_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07857__A2 _08741_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12730_ reg1_val[21] _12741_/B vssd1 vssd1 vccd1 vccd1 _12730_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_84_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12661_ _12661_/A _12661_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[7] sky130_fd_sc_hd__xor2_4
XFILLER_0_77_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11612_ _11785_/A _11613_/B vssd1 vssd1 vccd1 vccd1 _11614_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_107_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12592_ _12623_/A _12592_/B vssd1 vssd1 vccd1 vccd1 _12593_/B sky130_fd_sc_hd__or2_1
XFILLER_0_65_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11989__B _12214_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11543_ _10113_/A _11012_/B _11024_/Y _12254_/A1 _11542_/X vssd1 vssd1 vccd1 vccd1
+ _11543_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_65_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11474_ _11475_/A _11475_/B _11475_/C vssd1 vssd1 vccd1 vccd1 _11476_/A sky130_fd_sc_hd__o21ai_1
X_13213_ hold281/X _13213_/A2 _13212_/X _13213_/B2 vssd1 vssd1 vccd1 vccd1 _13214_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10425_ _10423_/Y _10425_/B vssd1 vssd1 vccd1 vccd1 _10428_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_21_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13144_ _12891_/X _13144_/B vssd1 vssd1 vccd1 vccd1 _13145_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_110_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12118__A1 _12394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10356_ _10356_/A _10356_/B vssd1 vssd1 vccd1 vccd1 _10358_/B sky130_fd_sc_hd__xnor2_2
X_13075_ _09716_/A _13077_/A2 hold98/X vssd1 vssd1 vccd1 vccd1 _13340_/D sky130_fd_sc_hd__o21a_1
XANTENNA__06611__B _06612_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10287_ _11269_/A _10287_/B vssd1 vssd1 vccd1 vccd1 _10288_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_20_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12026_ _12025_/A _12026_/B vssd1 vssd1 vccd1 vccd1 _12026_/X sky130_fd_sc_hd__and2b_1
XANTENNA__07723__A _08745_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13094__A2 _06892_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06765__A_N _07036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12928_ _13139_/B _13140_/A _12893_/X vssd1 vssd1 vccd1 vccd1 _13145_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_87_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12859_ hold268/A hold11/X vssd1 vssd1 vccd1 vccd1 _12860_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_118_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_4_3_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08273__A2 _08741_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12076__A _12076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08050_ _08069_/A _08069_/B vssd1 vssd1 vccd1 vccd1 _08050_/Y sky130_fd_sc_hd__nand2b_1
X_07001_ reg1_val[26] _07254_/B _06999_/X _07364_/B1 vssd1 vssd1 vccd1 vccd1 _07002_/B
+ sky130_fd_sc_hd__o31a_2
XFILLER_0_12_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12804__A _12804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06802__A _09343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08952_ _08954_/A _08954_/B vssd1 vssd1 vccd1 vccd1 _08952_/Y sky130_fd_sc_hd__nand2_1
X_08883_ _08885_/A _08885_/B vssd1 vssd1 vccd1 vccd1 _08883_/X sky130_fd_sc_hd__and2b_1
X_07903_ _07903_/A _07913_/A _07903_/C vssd1 vssd1 vccd1 vccd1 _07972_/A sky130_fd_sc_hd__or3_1
X_07834_ _07853_/A _07853_/B _07830_/X vssd1 vssd1 vccd1 vccd1 _07836_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07765_ fanout75/X fanout99/X _12818_/A _08304_/B vssd1 vssd1 vccd1 vccd1 _07766_/B
+ sky130_fd_sc_hd__o22a_1
X_06716_ _06981_/A reg1_val[14] vssd1 vssd1 vccd1 vccd1 _06716_/Y sky130_fd_sc_hd__nand2b_1
X_09504_ _09500_/X _09503_/X _11231_/S vssd1 vssd1 vccd1 vccd1 _09504_/X sky130_fd_sc_hd__mux2_1
X_07696_ _07986_/B _07696_/B vssd1 vssd1 vccd1 vccd1 _07719_/A sky130_fd_sc_hd__or2_1
XFILLER_0_39_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11155__A _12261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06647_ _12389_/A _06647_/B _12293_/A vssd1 vssd1 vccd1 vccd1 _06647_/X sky130_fd_sc_hd__or3_1
XFILLER_0_79_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09435_ _09435_/A _09435_/B vssd1 vssd1 vccd1 vccd1 _09439_/A sky130_fd_sc_hd__xor2_1
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06578_ rst vssd1 vssd1 vccd1 vccd1 _06578_/Y sky130_fd_sc_hd__inv_2
X_09366_ _10250_/S _09365_/X _09176_/B vssd1 vssd1 vccd1 vccd1 _09367_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_93_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_40 pred_val vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09297_ _09298_/A _09298_/B vssd1 vssd1 vccd1 vccd1 _09297_/X sky130_fd_sc_hd__and2_1
X_08317_ _08327_/A _08327_/B vssd1 vssd1 vccd1 vccd1 _08317_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_35_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_62 instruction[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07472__B1 _12836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_51 reg1_val[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10071__A2 _10574_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08248_ _08248_/A _08297_/A vssd1 vssd1 vccd1 vccd1 _08254_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_22_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10210_ _10211_/A _10211_/B _10211_/C vssd1 vssd1 vccd1 vccd1 _10210_/X sky130_fd_sc_hd__o21a_1
X_08179_ _08240_/A _08240_/B _08172_/X vssd1 vssd1 vccd1 vccd1 _08200_/A sky130_fd_sc_hd__a21o_1
X_11190_ _11188_/X _11190_/B vssd1 vssd1 vccd1 vccd1 _11191_/B sky130_fd_sc_hd__nand2b_1
X_10141_ _09854_/B _09958_/B _10275_/B _12426_/A vssd1 vssd1 vccd1 vccd1 _10141_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__11571__A2 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10072_ _11180_/A _10072_/B vssd1 vssd1 vccd1 vccd1 _10073_/B sky130_fd_sc_hd__xor2_2
XANTENNA__10531__B1 _10530_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07543__A _10422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10974_ _10974_/A _10974_/B vssd1 vssd1 vccd1 vccd1 _10976_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__11065__A _11065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12823__A2 _12830_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12713_ _12709_/B _12725_/A vssd1 vssd1 vccd1 vccd1 _12715_/A sky130_fd_sc_hd__nand2b_2
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12644_ reg1_val[4] _12644_/B vssd1 vssd1 vccd1 vccd1 _12645_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_108_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12575_ _12582_/A _12575_/B vssd1 vssd1 vccd1 vccd1 _12576_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_93_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11526_ _12174_/S _11526_/B vssd1 vssd1 vccd1 vccd1 _11526_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__07463__B1 _12814_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11457_ _09156_/Y _11437_/X _11444_/X _11456_/Y vssd1 vssd1 vccd1 vccd1 _11457_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_110_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10408_ curr_PC[9] _10779_/D vssd1 vssd1 vccd1 vccd1 _10409_/B sky130_fd_sc_hd__or2_1
X_11388_ _11389_/A _11389_/B vssd1 vssd1 vccd1 vccd1 _11475_/B sky130_fd_sc_hd__and2_1
XFILLER_0_21_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13127_ hold273/X _12789_/B _13126_/X _12790_/A vssd1 vssd1 vccd1 vccd1 hold274/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11562__A2 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10339_ _10454_/B _10339_/B vssd1 vssd1 vccd1 vccd1 _10341_/B sky130_fd_sc_hd__nor2_1
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13058_ _13331_/Q _12791_/A _13080_/B1 hold137/X _13128_/A vssd1 vssd1 vccd1 vccd1
+ hold138/A sky130_fd_sc_hd__o221a_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12009_ _12009_/A _12009_/B vssd1 vssd1 vccd1 vccd1 _12010_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_17_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08191__A1 _08723_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13067__A2 _13087_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08191__B2 _07885_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08730__A3 _08038_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07550_ _08671_/B2 fanout9/A fanout5/X _12794_/A vssd1 vssd1 vccd1 vccd1 _07551_/B
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_17_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09220_ _09220_/A _09220_/B vssd1 vssd1 vccd1 vccd1 _09223_/B sky130_fd_sc_hd__xor2_1
X_07481_ _07481_/A _07481_/B vssd1 vssd1 vccd1 vccd1 _07502_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_76_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_84 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09151_ _12429_/B _09147_/X _09150_/X _06923_/Y vssd1 vssd1 vccd1 vccd1 _09151_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_8_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09082_ _09542_/A _09079_/B _09079_/Y _11707_/A vssd1 vssd1 vccd1 vccd1 _09082_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_44_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10319__A _10444_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08102_ _08733_/A _08102_/B vssd1 vssd1 vccd1 vccd1 _08106_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_71_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08033_ _08033_/A _08033_/B vssd1 vssd1 vccd1 vccd1 _08034_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__12534__A _12692_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07206__B1 _06691_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07757__A1 _08752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07757__B2 _08798_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09984_ _09837_/A _09982_/X _09983_/Y _06939_/Y _06774_/B vssd1 vssd1 vccd1 vccd1
+ _09984_/X sky130_fd_sc_hd__o32a_1
XANTENNA__06980__A2 _07074_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08935_ _08936_/A _08936_/B vssd1 vssd1 vccd1 vccd1 _08935_/X sky130_fd_sc_hd__and2_1
X_08866_ _08835_/A _08833_/X _08832_/X vssd1 vssd1 vccd1 vccd1 _08869_/B sky130_fd_sc_hd__a21oi_4
XANTENNA__08182__A1 _08721_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07817_ _07816_/B _07816_/C _07816_/A vssd1 vssd1 vccd1 vccd1 _07818_/C sky130_fd_sc_hd__a21oi_1
X_08797_ _11385_/A _08797_/B vssd1 vssd1 vccd1 vccd1 _08801_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__08182__B2 _08739_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07748_ _08731_/A _07748_/B vssd1 vssd1 vccd1 vccd1 _07856_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__12805__A2 _12818_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10816__A1 _10444_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07679_ _08959_/B _08959_/A vssd1 vssd1 vccd1 vccd1 _07679_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_90_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09418_ _09418_/A _09418_/B vssd1 vssd1 vccd1 vccd1 _09420_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10690_ fanout23/X _09745_/B _10574_/B _11171_/A vssd1 vssd1 vccd1 vccd1 _10691_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout23_A fanout24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08194__A _08724_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09349_ hold248/A hold290/A _10391_/A2 _12401_/B1 _09348_/Y vssd1 vssd1 vccd1 vccd1
+ _09361_/B sky130_fd_sc_hd__a311o_1
XFILLER_0_109_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12360_ _09153_/Y _09497_/Y _09512_/Y _09142_/S _12359_/X vssd1 vssd1 vccd1 vccd1
+ _12360_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_62_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10229__A _10231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11311_ _11311_/A _11311_/B vssd1 vssd1 vccd1 vccd1 _11313_/B sky130_fd_sc_hd__and2_1
X_12291_ _06605_/Y _12195_/S _12176_/Y _06606_/A vssd1 vssd1 vccd1 vccd1 _12291_/X
+ sky130_fd_sc_hd__o31a_1
X_11242_ hold271/A _11452_/B1 _11339_/B _12247_/C1 vssd1 vssd1 vccd1 vccd1 _11243_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_120_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11173_ _11172_/B _11172_/C _11172_/A vssd1 vssd1 vccd1 vccd1 _11177_/B sky130_fd_sc_hd__a21o_1
X_10124_ hold258/A hold291/A _10124_/C vssd1 vssd1 vccd1 vccd1 _10256_/B sky130_fd_sc_hd__or3_2
XFILLER_0_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10055_ _10056_/A _10056_/B _10056_/C vssd1 vssd1 vccd1 vccd1 _10218_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_54_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08173__A1 _08741_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08173__B2 _08727_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07920__A1 fanout99/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07920__B2 _12818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10807__A1 _10418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10807__B2 _09745_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10957_ _10957_/A _10957_/B vssd1 vssd1 vccd1 vccd1 _10966_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_45_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11480__A1 _11766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11480__B2 _11847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10888_ _11886_/A _10888_/B _10887_/X vssd1 vssd1 vccd1 vccd1 _10888_/X sky130_fd_sc_hd__or3b_1
XFILLER_0_38_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12627_ _12631_/A _12627_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[0] sky130_fd_sc_hd__and2_4
XFILLER_0_115_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08228__A2 fanout87/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12558_ reg1_val[17] curr_PC[17] _12586_/S vssd1 vssd1 vccd1 vccd1 _12559_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_81_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold107 hold107/A vssd1 vssd1 vccd1 vccd1 hold107/X sky130_fd_sc_hd__dlygate4sd3_1
X_12489_ _12495_/B _12489_/B vssd1 vssd1 vccd1 vccd1 new_PC[6] sky130_fd_sc_hd__and2_4
XFILLER_0_81_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09647__B _09647_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11509_ _11507_/Y _11509_/B vssd1 vssd1 vccd1 vccd1 _11700_/A sky130_fd_sc_hd__nand2b_2
Xhold118 hold118/A vssd1 vssd1 vccd1 vccd1 hold118/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold129 hold129/A vssd1 vssd1 vccd1 vccd1 hold129/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09139__S _09142_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07448__A _11673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08400__A2 fanout87/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06981_ _06981_/A _06981_/B vssd1 vssd1 vccd1 vccd1 _12822_/A sky130_fd_sc_hd__xnor2_4
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08720_ _09028_/A _09028_/B _09036_/A _08718_/Y vssd1 vssd1 vccd1 vccd1 _09033_/A
+ sky130_fd_sc_hd__a31o_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08651_ _08652_/A _08643_/B _08643_/C _08689_/A vssd1 vssd1 vccd1 vccd1 _08653_/A
+ sky130_fd_sc_hd__a31o_1
XANTENNA__10321__B fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07602_ _07602_/A _07602_/B vssd1 vssd1 vccd1 vccd1 _07678_/A sky130_fd_sc_hd__xnor2_4
X_08582_ _08681_/A _08582_/B vssd1 vssd1 vccd1 vccd1 _08612_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_88_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07533_ _09746_/A _07533_/B _07533_/C vssd1 vssd1 vccd1 vccd1 _07540_/A sky130_fd_sc_hd__and3_1
XFILLER_0_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout158_A _08980_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07464_ _10422_/A _07464_/B vssd1 vssd1 vccd1 vccd1 _07568_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_48_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11471__B2 _11269_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09203_ _09203_/A _09203_/B vssd1 vssd1 vccd1 vccd1 _09205_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_76_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09134_ reg1_val[2] reg1_val[29] _09142_/S vssd1 vssd1 vccd1 vccd1 _09134_/X sky130_fd_sc_hd__mux2_1
X_07395_ _07395_/A _07395_/B vssd1 vssd1 vccd1 vccd1 _07399_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_44_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12420__B1 _12290_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08742__A _08742_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12264__A _12264_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09065_ _09065_/A _09065_/B _09065_/C _09065_/D vssd1 vssd1 vccd1 vccd1 _09066_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_0_4_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08016_ _08016_/A _08016_/B vssd1 vssd1 vccd1 vccd1 _08017_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_4_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09967_ _11233_/S _09966_/A _09182_/B vssd1 vssd1 vccd1 vccd1 _09968_/A sky130_fd_sc_hd__a21o_1
X_08918_ _08918_/A _08918_/B vssd1 vssd1 vccd1 vccd1 _08920_/A sky130_fd_sc_hd__or2_1
XANTENNA__09352__B1 _11624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09898_ _09898_/A _09898_/B vssd1 vssd1 vccd1 vccd1 _09900_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__08155__A1 fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08155__B2 _08304_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10231__B _10231_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08849_ _08849_/A _08849_/B vssd1 vssd1 vccd1 vccd1 _08863_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_79_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11860_ _11861_/A _11861_/B _11861_/C vssd1 vssd1 vccd1 vccd1 _11863_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_79_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11791_ _11790_/A _11822_/B _12290_/A vssd1 vssd1 vccd1 vccd1 _11791_/X sky130_fd_sc_hd__a21o_1
XANTENNA__07821__A _07821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10811_ fanout23/X _10574_/B _10575_/B _11171_/A vssd1 vssd1 vccd1 vccd1 _10812_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11343__A _11343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10742_ _10233_/X _10234_/X _10741_/X vssd1 vssd1 vccd1 vccd1 _10742_/X sky130_fd_sc_hd__a21o_1
XANTENNA__11462__A1 _11653_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11462__B2 _08752_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10673_ _07087_/A _07087_/B fanout48/X _10570_/B fanout66/X vssd1 vssd1 vccd1 vccd1
+ _10674_/B sky130_fd_sc_hd__o32a_1
X_13392_ instruction[8] vssd1 vssd1 vccd1 vccd1 pred_idx[0] sky130_fd_sc_hd__buf_12
XFILLER_0_63_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12412_ _12412_/A _12412_/B vssd1 vssd1 vccd1 vccd1 _12417_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_105_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12343_ _12341_/X _12342_/Y _06647_/B vssd1 vssd1 vccd1 vccd1 _12345_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_63_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08091__B1 _08617_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08630__A2 _08661_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12274_ _12275_/A _12275_/B vssd1 vssd1 vccd1 vccd1 _12327_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_120_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11225_ _11224_/A _11224_/B _11224_/Y _09156_/Y vssd1 vssd1 vccd1 vccd1 _11250_/A
+ sky130_fd_sc_hd__o211a_1
XANTENNA__09186__A3 _09168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11156_ fanout29/X _11751_/A _11766_/A fanout27/X vssd1 vssd1 vccd1 vccd1 _11157_/B
+ sky130_fd_sc_hd__o22a_1
X_10107_ _06775_/Y _09962_/X _06777_/B vssd1 vssd1 vccd1 vccd1 _10107_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_65_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11518__A _11649_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10422__A _10422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11087_ _11088_/A _11088_/B _11088_/C vssd1 vssd1 vccd1 vccd1 _11089_/A sky130_fd_sc_hd__a21oi_1
X_10038_ _12076_/A _10038_/B vssd1 vssd1 vccd1 vccd1 _10040_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_105_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11989_ _11989_/A _12214_/B vssd1 vssd1 vccd1 vccd1 _11990_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_46_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07180_ _11163_/A _07180_/B vssd1 vssd1 vccd1 vccd1 _07603_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10008__A2 _12214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11756__A2 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07178__A _11020_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12812__A _12812_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09821_ _11233_/S _09820_/Y _09182_/B vssd1 vssd1 vccd1 vccd1 _09821_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_39_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11428__A _11649_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09752_ _09752_/A _09752_/B vssd1 vssd1 vccd1 vccd1 _09755_/A sky130_fd_sc_hd__nor2_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06964_ _06964_/A _06964_/B _06967_/C vssd1 vssd1 vccd1 vccd1 _07074_/C sky130_fd_sc_hd__or3_2
X_08703_ _08703_/A _08703_/B vssd1 vssd1 vccd1 vccd1 _09006_/A sky130_fd_sc_hd__nor2_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10332__A _11673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09683_ _09523_/A _09523_/B _06798_/B vssd1 vssd1 vccd1 vccd1 _09684_/C sky130_fd_sc_hd__a21boi_1
X_06895_ instruction[12] _06896_/B vssd1 vssd1 vccd1 vccd1 dest_pred[1] sky130_fd_sc_hd__and2_4
X_08634_ _08635_/B _08635_/C _09442_/A vssd1 vssd1 vccd1 vccd1 _08636_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_68_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_82 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08565_ _08584_/A _08565_/B vssd1 vssd1 vccd1 vccd1 _08591_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__07641__A _11908_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11444__A1 _12394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07516_ _07517_/A _07517_/B vssd1 vssd1 vccd1 vccd1 _07516_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_77_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07648__B1 _11766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout13 _12854_/A vssd1 vssd1 vccd1 vccd1 fanout13/X sky130_fd_sc_hd__buf_4
XANTENNA__11163__A _11163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08496_ _07896_/A _09238_/B _08656_/B _08723_/B1 vssd1 vssd1 vccd1 vccd1 _08497_/B
+ sky130_fd_sc_hd__o22a_1
Xfanout46 _07194_/X vssd1 vssd1 vccd1 vccd1 _12840_/A sky130_fd_sc_hd__clkbuf_8
Xfanout35 _07504_/Y vssd1 vssd1 vccd1 vccd1 _12264_/B sky130_fd_sc_hd__buf_8
XFILLER_0_64_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout24 _07048_/X vssd1 vssd1 vccd1 vccd1 fanout24/X sky130_fd_sc_hd__buf_6
XFILLER_0_9_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout57 _07150_/Y vssd1 vssd1 vccd1 vccd1 _10941_/B sky130_fd_sc_hd__buf_6
X_07447_ fanout30/X _12804_/A _09768_/A1 _07688_/B vssd1 vssd1 vccd1 vccd1 _07448_/B
+ sky130_fd_sc_hd__o22a_1
Xfanout79 _12832_/A vssd1 vssd1 vccd1 vccd1 _11558_/A sky130_fd_sc_hd__buf_6
Xfanout68 fanout69/X vssd1 vssd1 vccd1 vccd1 _10941_/A sky130_fd_sc_hd__clkbuf_8
XANTENNA__11995__A2 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07378_ _07378_/A _07378_/B vssd1 vssd1 vccd1 vccd1 _07395_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__09568__A _09568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09117_ reg1_val[9] reg1_val[22] _09142_/S vssd1 vssd1 vccd1 vccd1 _09117_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_17_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06704__B _11343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09048_ _08884_/Y _08897_/X _08899_/B vssd1 vssd1 vccd1 vccd1 _09048_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_5_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07820__B1 _08671_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout90_A _07178_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11010_ _09972_/B _09975_/Y _11010_/S vssd1 vssd1 vccd1 vccd1 _11010_/X sky130_fd_sc_hd__mux2_1
XANTENNA__07179__A2 _10948_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10183__A1 _10941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10183__B2 fanout94/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12961_ _13214_/A _12961_/B vssd1 vssd1 vccd1 vccd1 _13283_/D sky130_fd_sc_hd__and2_1
XANTENNA__08679__A2 _09251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12892_ hold285/X hold45/X vssd1 vssd1 vccd1 vccd1 _13144_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_87_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08647__A _08728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07887__B1 _11385_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11912_ _11912_/A _11912_/B vssd1 vssd1 vccd1 vccd1 _11913_/B sky130_fd_sc_hd__nor2_1
XANTENNA__10388__S _11886_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07551__A _12264_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07351__A2 _12828_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11843_ _11989_/A fanout9/X fanout4/X _11923_/A vssd1 vssd1 vccd1 vccd1 _11844_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11774_ _11775_/A _11775_/B vssd1 vssd1 vccd1 vccd1 _11824_/B sky130_fd_sc_hd__nand2b_1
XTAP_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10725_ _10725_/A _10725_/B vssd1 vssd1 vccd1 vccd1 _10727_/B sky130_fd_sc_hd__xnor2_1
X_10656_ curr_PC[10] _10656_/B vssd1 vssd1 vccd1 vccd1 _10656_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08064__B1 _07885_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13375_ _13376_/CLK _13375_/D vssd1 vssd1 vccd1 vccd1 hold266/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_4_8_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10587_ _10465_/A _10465_/B _10468_/X vssd1 vssd1 vccd1 vccd1 _10594_/A sky130_fd_sc_hd__o21ba_1
X_12326_ _12373_/B _12326_/B vssd1 vssd1 vccd1 vccd1 _12327_/C sky130_fd_sc_hd__or2_1
X_12257_ _12428_/A _12238_/Y _12256_/Y _12236_/X vssd1 vssd1 vccd1 vccd1 _12257_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12188_ _11636_/B _12245_/B hold281/A vssd1 vssd1 vccd1 vccd1 _12190_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__07726__A _08742_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11208_ _11210_/A _11210_/B _11210_/C vssd1 vssd1 vccd1 vccd1 _11211_/A sky130_fd_sc_hd__a21oi_1
X_11139_ curr_PC[13] curr_PC[14] _11139_/C vssd1 vssd1 vccd1 vccd1 _11253_/B sky130_fd_sc_hd__and3_1
XANTENNA__13112__B2 _06572_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06680_ reg1_val[19] _07210_/A vssd1 vssd1 vccd1 vccd1 _06680_/X sky130_fd_sc_hd__and2_1
XFILLER_0_116_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08350_ _09768_/A1 _09567_/B _09568_/B _07885_/B vssd1 vssd1 vccd1 vccd1 _08351_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_74_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07301_ _08000_/A _07303_/B vssd1 vssd1 vccd1 vccd1 _07301_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08281_ _08301_/A _08301_/B _08270_/X vssd1 vssd1 vccd1 vccd1 _08291_/A sky130_fd_sc_hd__a21boi_1
XFILLER_0_128_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09388__A _11673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07232_ _07604_/A _07232_/B vssd1 vssd1 vccd1 vccd1 _07233_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_41_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11729__A2 _11343_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07163_ _09897_/A _07167_/A vssd1 vssd1 vccd1 vccd1 _07163_/X sky130_fd_sc_hd__or2_1
XFILLER_0_54_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07094_ _07089_/A _06964_/A _06964_/B _07074_/B vssd1 vssd1 vccd1 vccd1 _07095_/B
+ sky130_fd_sc_hd__o31a_2
XFILLER_0_14_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout203 _12790_/Y vssd1 vssd1 vccd1 vccd1 _12830_/B sky130_fd_sc_hd__buf_4
XANTENNA__08358__B2 _07149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08358__A1 _12818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout247 _11452_/B1 vssd1 vssd1 vccd1 vccd1 _09835_/B sky130_fd_sc_hd__buf_4
Xfanout236 _11231_/S vssd1 vssd1 vccd1 vccd1 _11010_/S sky130_fd_sc_hd__buf_4
X_09804_ _09804_/A _09804_/B vssd1 vssd1 vccd1 vccd1 _09805_/B sky130_fd_sc_hd__xor2_4
Xfanout225 _12794_/A vssd1 vssd1 vccd1 vccd1 _08752_/A sky130_fd_sc_hd__clkbuf_8
Xfanout269 _06770_/X vssd1 vssd1 vccd1 vccd1 _12429_/B sky130_fd_sc_hd__clkbuf_4
Xfanout258 _09442_/A vssd1 vssd1 vccd1 vccd1 _08731_/A sky130_fd_sc_hd__buf_12
X_07996_ _07996_/A _07996_/B vssd1 vssd1 vccd1 vccd1 _07997_/B sky130_fd_sc_hd__xnor2_1
X_06947_ reg1_val[10] _07200_/B _07200_/A vssd1 vssd1 vccd1 vccd1 _06948_/B sky130_fd_sc_hd__o21a_1
X_09735_ _10710_/A _09735_/B vssd1 vssd1 vccd1 vccd1 _09743_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__09858__A1 _11065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09666_ _09326_/X _09336_/X _09666_/S vssd1 vssd1 vccd1 vccd1 _09666_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12311__C1 _12310_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09858__B2 _11146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11665__B2 _11989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11665__A1 _11923_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06878_ _06926_/A instruction[4] vssd1 vssd1 vccd1 vccd1 _09165_/A sky130_fd_sc_hd__or2_2
X_08617_ _08673_/A _08617_/B vssd1 vssd1 vccd1 vccd1 _08628_/A sky130_fd_sc_hd__nor2_1
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09597_ _09597_/A _09597_/B vssd1 vssd1 vccd1 vccd1 _09606_/A sky130_fd_sc_hd__xor2_2
X_08548_ _08549_/A _08549_/B vssd1 vssd1 vccd1 vccd1 _08571_/A sky130_fd_sc_hd__nor2_1
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07090__B _07090_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08479_ _08508_/A _08508_/B vssd1 vssd1 vccd1 vccd1 _08518_/A sky130_fd_sc_hd__nor2_1
XANTENNA__11621__A _12423_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10510_ reg1_val[9] curr_PC[9] vssd1 vssd1 vccd1 vccd1 _10510_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_80_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09298__A _09298_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11490_ _11398_/A _11397_/B _11397_/A vssd1 vssd1 vccd1 vccd1 _11501_/A sky130_fd_sc_hd__o21ba_1
X_10441_ _10441_/A _10441_/B vssd1 vssd1 vccd1 vccd1 _10459_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_17_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08597__A1 _07752_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13160_ _13160_/A _13160_/B vssd1 vssd1 vccd1 vccd1 _13160_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_115_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08597__B2 _12802_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10372_ _11874_/A _10410_/A _10658_/B vssd1 vssd1 vccd1 vccd1 _10372_/Y sky130_fd_sc_hd__a21oi_1
X_13091_ _13109_/A hold303/X vssd1 vssd1 vccd1 vccd1 _13347_/D sky130_fd_sc_hd__and2_1
XFILLER_0_103_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12111_ _12110_/A _12110_/B _12110_/Y _11624_/A vssd1 vssd1 vccd1 vccd1 _12111_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__09745__B _09745_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12042_ _10246_/X _12041_/Y _12244_/S vssd1 vssd1 vccd1 vccd1 _12042_/X sky130_fd_sc_hd__mux2_1
Xhold290 hold290/A vssd1 vssd1 vccd1 vccd1 hold290/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11353__B1 _11352_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10156__A1 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10156__B2 _07688_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11105__B1 _11707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12944_ _13193_/A _12943_/B _12874_/X vssd1 vssd1 vccd1 vccd1 _13198_/A sky130_fd_sc_hd__a21o_1
XANTENNA__06780__B1 _06778_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12875_ hold9/X hold275/A vssd1 vssd1 vccd1 vccd1 _12875_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_87_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11826_ _12067_/A fanout15/X fanout36/X _12150_/A vssd1 vssd1 vccd1 vccd1 _11827_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11757_ _12073_/A _11757_/B vssd1 vssd1 vccd1 vccd1 _11758_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_126_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10708_ fanout74/X fanout56/X _09568_/A _10948_/B2 vssd1 vssd1 vccd1 vccd1 _10709_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_71_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11688_ _11688_/A _11688_/B vssd1 vssd1 vccd1 vccd1 _11689_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_11_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10639_ _10635_/Y _10636_/X _12244_/S vssd1 vssd1 vccd1 vccd1 _10639_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_3_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10919__B1 _11923_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13358_ _13365_/CLK _13358_/D vssd1 vssd1 vccd1 vccd1 hold285/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12309_ _09111_/S _09672_/X _12299_/B _09152_/Y _12308_/X vssd1 vssd1 vccd1 vccd1
+ _12309_/Y sky130_fd_sc_hd__a221oi_2
XFILLER_0_51_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07260__A1 _12076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13289_ _13311_/CLK _13289_/D vssd1 vssd1 vccd1 vccd1 hold157/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09147__S _09147_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07850_ _07824_/X _07849_/Y _07848_/X _07807_/B vssd1 vssd1 vccd1 vccd1 _07850_/X
+ sky130_fd_sc_hd__o211a_1
X_06801_ _06805_/A _06702_/A _12634_/B _06799_/X vssd1 vssd1 vccd1 vccd1 _09505_/S
+ sky130_fd_sc_hd__a31o_2
X_07781_ _07781_/A _07781_/B _07781_/C vssd1 vssd1 vccd1 vccd1 _07782_/B sky130_fd_sc_hd__and3_1
X_09520_ _10391_/A2 _09519_/X hold238/A vssd1 vssd1 vccd1 vccd1 _09520_/Y sky130_fd_sc_hd__a21oi_1
X_06732_ reg2_val[11] _06799_/B vssd1 vssd1 vccd1 vccd1 _06732_/X sky130_fd_sc_hd__and2_1
XFILLER_0_78_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06663_ instruction[30] _06694_/B vssd1 vssd1 vccd1 vccd1 _12649_/B sky130_fd_sc_hd__and2_4
X_09451_ _09452_/A _09452_/B vssd1 vssd1 vccd1 vccd1 _09453_/A sky130_fd_sc_hd__or2_1
X_06594_ instruction[41] _06897_/B _06591_/X vssd1 vssd1 vccd1 vccd1 _06635_/A sky130_fd_sc_hd__a21oi_4
XFILLER_0_93_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09382_ fanout23/X _12812_/A _12814_/A _07819_/B vssd1 vssd1 vccd1 vccd1 _09383_/B
+ sky130_fd_sc_hd__o22a_1
X_08402_ _08405_/A _08405_/B vssd1 vssd1 vccd1 vccd1 _08402_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_47_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07079__A1 _07036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08333_ _08383_/A _08383_/B vssd1 vssd1 vccd1 vccd1 _08384_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08276__B1 _08564_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout140_A _07089_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08264_ _08731_/A _08264_/B vssd1 vssd1 vccd1 vccd1 _08266_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_116_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07215_ reg1_val[8] _07215_/B vssd1 vssd1 vccd1 vccd1 _07217_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08195_ _08432_/B _07896_/A _07955_/A _10537_/A1 vssd1 vssd1 vccd1 vccd1 _08196_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08579__A1 _12802_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08579__B2 _12804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07146_ _09444_/A _12846_/A _09236_/B2 _12848_/A vssd1 vssd1 vccd1 vccd1 _07147_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_30_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07077_ _10664_/A _10941_/A _10818_/A fanout94/X vssd1 vssd1 vccd1 vccd1 _07078_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07366__A _09548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07979_ _08024_/B _08024_/A vssd1 vssd1 vccd1 vccd1 _07979_/Y sky130_fd_sc_hd__nand2b_1
X_09718_ _09718_/A _09718_/B vssd1 vssd1 vccd1 vccd1 _09719_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_69_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout53_A _12842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10990_ _11102_/B _11100_/A vssd1 vssd1 vccd1 vccd1 _11215_/A sky130_fd_sc_hd__or2_1
XFILLER_0_69_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09649_ _09706_/A _09649_/B _09953_/A _09953_/B vssd1 vssd1 vccd1 vccd1 wire3/A sky130_fd_sc_hd__nor4_1
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12660_ _12658_/Y _12660_/B vssd1 vssd1 vccd1 vccd1 _12661_/B sky130_fd_sc_hd__nand2b_2
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08267__B1 _08727_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11611_ _10744_/B _11215_/X _11609_/Y _11610_/Y vssd1 vssd1 vccd1 vccd1 _11613_/B
+ sky130_fd_sc_hd__o31a_2
X_12591_ _12623_/A _12592_/B vssd1 vssd1 vccd1 vccd1 _12591_/X sky130_fd_sc_hd__and2_1
XFILLER_0_108_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11542_ _07131_/B _11343_/B _11541_/X _06693_/B vssd1 vssd1 vccd1 vccd1 _11542_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_53_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11473_ _11557_/A _11473_/B vssd1 vssd1 vccd1 vccd1 _11475_/C sky130_fd_sc_hd__xnor2_1
X_13212_ hold261/X _13211_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13212_/X sky130_fd_sc_hd__mux2_1
XANTENNA__11023__C1 _11022_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10424_ _10424_/A _10424_/B _10424_/C vssd1 vssd1 vccd1 vccd1 _10425_/B sky130_fd_sc_hd__nand3_1
X_13143_ _13235_/A hold286/X vssd1 vssd1 vccd1 vccd1 _13358_/D sky130_fd_sc_hd__and2_1
XANTENNA__07276__A _10422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10355_ _10356_/A _10356_/B vssd1 vssd1 vccd1 vccd1 _10412_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_20_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13074_ hold97/X _12791_/A _13080_/B1 hold67/X _13113_/A vssd1 vssd1 vccd1 vccd1
+ hold98/A sky130_fd_sc_hd__o221a_1
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10286_ _10571_/A fanout48/X _10930_/B _10570_/A vssd1 vssd1 vccd1 vccd1 _10287_/B
+ sky130_fd_sc_hd__o22a_1
X_12025_ _12025_/A vssd1 vssd1 vccd1 vccd1 _12025_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13217__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11526__A _12174_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12927_ _13134_/B _13135_/A _12895_/X vssd1 vssd1 vccd1 vccd1 _13140_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_88_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12858_ hold11/X hold268/A vssd1 vssd1 vccd1 vccd1 _12860_/A sky130_fd_sc_hd__and2b_1
X_11809_ _11636_/B _11888_/B hold252/A vssd1 vssd1 vccd1 vccd1 _11809_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__12054__A1 _09172_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08258__B1 _08304_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12789_ rst _12789_/B _12789_/C vssd1 vssd1 vccd1 vccd1 _13249_/D sky130_fd_sc_hd__nor3_1
XFILLER_0_113_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11261__A _11261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07000_ _07254_/B _06999_/X _07364_/B1 vssd1 vssd1 vccd1 vccd1 _07010_/B sky130_fd_sc_hd__o21a_1
XANTENNA__12804__B _12818_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11565__B1 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08430__B1 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07186__A _09441_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08981__A1 _09445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08951_ _08951_/A _08951_/B vssd1 vssd1 vccd1 vccd1 _08954_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10324__B _10324_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12820__A _12820_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08882_ _08882_/A _08882_/B vssd1 vssd1 vccd1 vccd1 _08885_/B sky130_fd_sc_hd__xnor2_2
X_07902_ _07902_/A _07902_/B vssd1 vssd1 vccd1 vccd1 _07903_/C sky130_fd_sc_hd__nor2_1
X_07833_ _07833_/A _07833_/B vssd1 vssd1 vccd1 vccd1 _07853_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07764_ _08740_/A _07764_/B vssd1 vssd1 vccd1 vccd1 _07768_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_2_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09503_ _09501_/X _09502_/X _09503_/S vssd1 vssd1 vccd1 vccd1 _09503_/X sky130_fd_sc_hd__mux2_1
X_06715_ _06805_/A _06686_/A _12703_/B _06714_/X vssd1 vssd1 vccd1 vccd1 _06981_/A
+ sky130_fd_sc_hd__a31o_4
XFILLER_0_78_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07695_ _07694_/B _07695_/B vssd1 vssd1 vccd1 vccd1 _07696_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_2_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06646_ _12049_/S _06646_/B vssd1 vssd1 vccd1 vccd1 _06648_/D sky130_fd_sc_hd__nand2_2
X_09434_ _09435_/A _09435_/B vssd1 vssd1 vccd1 vccd1 _09434_/Y sky130_fd_sc_hd__nor2_1
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08745__A _08745_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09365_ _09133_/X _09181_/B _09666_/S vssd1 vssd1 vccd1 vccd1 _09365_/X sky130_fd_sc_hd__mux2_1
X_06577_ _12341_/A vssd1 vssd1 vccd1 vccd1 _06577_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_47_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11171__A _11171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_41 pred_val vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_30 reg2_val[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09296_ _09296_/A _09296_/B vssd1 vssd1 vccd1 vccd1 _09298_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_47_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08316_ _08314_/Y _08371_/B _08311_/Y vssd1 vssd1 vccd1 vccd1 _08327_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_34_215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_63 instruction[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07472__A1 _12838_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07472__B2 _10589_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_52 reg1_val[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08247_ _08296_/A _08296_/B vssd1 vssd1 vccd1 vccd1 _08297_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_15_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07224__A1 _07220_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08178_ _08178_/A _08178_/B vssd1 vssd1 vccd1 vccd1 _08240_/B sky130_fd_sc_hd__xor2_1
XANTENNA__11110__S _12174_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06712__B _06988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07129_ _07130_/A _11343_/A vssd1 vssd1 vccd1 vccd1 _07129_/X sky130_fd_sc_hd__and2_1
X_10140_ _10403_/C _10139_/Y _10780_/A _10137_/X vssd1 vssd1 vccd1 vccd1 dest_val[6]
+ sky130_fd_sc_hd__a2bb2o_4
X_10071_ _11146_/A _10574_/A _10575_/A _11294_/A vssd1 vssd1 vccd1 vccd1 _10072_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_100_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10531__A1 _11876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10973_ _10974_/A _10974_/B vssd1 vssd1 vccd1 vccd1 _11088_/A sky130_fd_sc_hd__or2_1
XANTENNA__11065__B _12412_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12712_ _12712_/A _12712_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[16] sky130_fd_sc_hd__xor2_4
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10295__B1 _10941_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08655__A _08655_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12643_ reg1_val[4] _12644_/B vssd1 vssd1 vccd1 vccd1 _12643_/Y sky130_fd_sc_hd__nor2_1
X_12574_ _12582_/C _12574_/B vssd1 vssd1 vccd1 vccd1 _12581_/C sky130_fd_sc_hd__nand2_2
XFILLER_0_93_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07058__A4 _06994_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11525_ _06700_/B _11435_/A _06698_/X vssd1 vssd1 vccd1 vccd1 _11526_/B sky130_fd_sc_hd__a21o_1
XANTENNA__07463__B2 _11653_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07463__A1 _10664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11547__B1 _11539_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11456_ _10113_/A _11121_/B _11448_/Y _11455_/X vssd1 vssd1 vccd1 vccd1 _11456_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_0_68_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10407_ curr_PC[9] _10779_/D vssd1 vssd1 vccd1 vccd1 _10656_/B sky130_fd_sc_hd__nand2_1
X_11387_ _11564_/A _11387_/B vssd1 vssd1 vccd1 vccd1 _11389_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13126_ hold294/A _13125_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13126_/X sky130_fd_sc_hd__mux2_1
X_10338_ _10338_/A _10338_/B vssd1 vssd1 vccd1 vccd1 _10339_/B sky130_fd_sc_hd__nor2_1
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13057_ _07076_/B _13087_/B2 hold77/X vssd1 vssd1 vccd1 vccd1 hold78/A sky130_fd_sc_hd__o21a_1
Xload_slew214 _09594_/A vssd1 vssd1 vccd1 vccd1 _08598_/A sky130_fd_sc_hd__buf_6
XANTENNA__06974__B1 _10706_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10269_ _09111_/S _10246_/X _10252_/X _09830_/A _10268_/X vssd1 vssd1 vccd1 vccd1
+ _10270_/D sky130_fd_sc_hd__a221o_1
XFILLER_0_84_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07734__A _08724_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12008_ _12010_/A vssd1 vssd1 vccd1 vccd1 _12089_/A sky130_fd_sc_hd__inv_2
XANTENNA__08191__A2 fanout87/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07480_ _10449_/A _07480_/B vssd1 vssd1 vccd1 vccd1 _07481_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_76_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10286__B1 _10930_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08565__A _08584_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11235__C1 _09172_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09150_ _09345_/A _09149_/X _11886_/A vssd1 vssd1 vccd1 vccd1 _09150_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_33_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09081_ _09165_/A _09170_/A vssd1 vssd1 vccd1 vccd1 _09081_/X sky130_fd_sc_hd__or2_1
XFILLER_0_44_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08101_ _08741_/B2 _08732_/A2 _08656_/B _08732_/A1 vssd1 vssd1 vccd1 vccd1 _08102_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09396__A _11294_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08032_ _08031_/A _08031_/C _08031_/B vssd1 vssd1 vccd1 vccd1 _08034_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_31_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08403__B1 _08432_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout103_A _11758_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09983_ hold258/A _09983_/B vssd1 vssd1 vccd1 vccd1 _09983_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__07757__A2 fanout24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08934_ _08934_/A _08934_/B vssd1 vssd1 vccd1 vccd1 _08936_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__07644__A _09716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09903__B1 _08507_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08865_ _08865_/A _08865_/B vssd1 vssd1 vccd1 vccd1 _08869_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_98_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07816_ _07816_/A _07816_/B _07816_/C vssd1 vssd1 vccd1 vccd1 _07818_/B sky130_fd_sc_hd__and3_1
X_08796_ _07955_/A fanout69/X _08216_/B _07896_/A vssd1 vssd1 vccd1 vccd1 _08797_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11166__A _11470_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08182__A2 _08744_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07747_ _06574_/Y _11989_/A _11923_/A _08436_/B vssd1 vssd1 vccd1 vccd1 _07748_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_79_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07678_ _07678_/A _07678_/B vssd1 vssd1 vccd1 vccd1 _08959_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_109_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06629_ _06635_/A _12673_/B vssd1 vssd1 vccd1 vccd1 _06629_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_90_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09417_ _09415_/A _09415_/B _09418_/B vssd1 vssd1 vccd1 vccd1 _09558_/A sky130_fd_sc_hd__o21bai_1
X_09348_ hold290/A _10391_/A2 hold248/A vssd1 vssd1 vccd1 vccd1 _09348_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_124_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10229__B _10231_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09279_ _09280_/A _09280_/B vssd1 vssd1 vccd1 vccd1 _09279_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_7_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11310_ _11310_/A _11310_/B vssd1 vssd1 vccd1 vccd1 _11313_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_105_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12290_ _12290_/A _12290_/B _12290_/C vssd1 vssd1 vccd1 vccd1 _12290_/X sky130_fd_sc_hd__or3_1
XANTENNA__07819__A _08752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11241_ _11341_/B _11339_/B hold271/A vssd1 vssd1 vccd1 vccd1 _11243_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_120_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11172_ _11172_/A _11172_/B _11172_/C vssd1 vssd1 vccd1 vccd1 _11177_/A sky130_fd_sc_hd__nand3_1
XANTENNA__10201__B1 _10930_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10123_ _10123_/A _10123_/B vssd1 vssd1 vccd1 vccd1 _10123_/Y sky130_fd_sc_hd__nor2_1
X_10054_ _10054_/A _10054_/B vssd1 vssd1 vccd1 vccd1 _10056_/C sky130_fd_sc_hd__xor2_1
XFILLER_0_89_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09370__B2 _09142_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09370__A1 _09163_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08173__A2 _08727_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07920__A2 fanout87/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10807__A2 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10956_ _10956_/A _10956_/B vssd1 vssd1 vccd1 vccd1 _10957_/B sky130_fd_sc_hd__or2_1
XFILLER_0_128_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10887_ _10884_/X _10885_/Y _10755_/X _10759_/A vssd1 vssd1 vccd1 vccd1 _10887_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__11480__A2 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06617__B _06838_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12626_ _12626_/A _12626_/B vssd1 vssd1 vccd1 vccd1 _12627_/B sky130_fd_sc_hd__or2_1
XFILLER_0_109_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13230__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12557_ _12566_/A _12557_/B vssd1 vssd1 vccd1 vccd1 new_PC[16] sky130_fd_sc_hd__and2_4
XANTENNA__08633__B1 _06574_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold108 hold108/A vssd1 vssd1 vccd1 vccd1 hold108/X sky130_fd_sc_hd__dlygate4sd3_1
X_12488_ _12488_/A _12488_/B _12488_/C vssd1 vssd1 vccd1 vccd1 _12489_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_79_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11508_ _11508_/A _11508_/B _11508_/C vssd1 vssd1 vccd1 vccd1 _11509_/B sky130_fd_sc_hd__nand3_2
Xhold119 hold119/A vssd1 vssd1 vccd1 vccd1 hold119/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11439_ reg1_val[17] curr_PC[17] vssd1 vssd1 vccd1 vccd1 _11439_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__09189__A1 _11142_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13109_ _13109_/A _13109_/B vssd1 vssd1 vccd1 vccd1 _13351_/D sky130_fd_sc_hd__and2_1
XANTENNA__06947__B1 _07200_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06980_ _11020_/A _07074_/A _07074_/C _07074_/B vssd1 vssd1 vccd1 vccd1 _06981_/B
+ sky130_fd_sc_hd__o31a_2
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07464__A _10422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08650_ _08650_/A _08650_/B _08650_/C vssd1 vssd1 vccd1 vccd1 _08689_/A sky130_fd_sc_hd__and3_1
XFILLER_0_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07601_ _07681_/A _07681_/B vssd1 vssd1 vccd1 vccd1 _07601_/X sky130_fd_sc_hd__and2_1
XFILLER_0_89_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08581_ _08730_/A1 _12808_/A _08038_/A _09768_/A1 vssd1 vssd1 vccd1 vccd1 _08582_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07124__B1 _07200_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06808__A _07149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07532_ _11065_/A _10571_/A vssd1 vssd1 vccd1 vccd1 _07533_/C sky130_fd_sc_hd__or2_1
XFILLER_0_76_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07463_ _10664_/A fanout66/X _12814_/A _11653_/A vssd1 vssd1 vccd1 vccd1 _07464_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_48_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09202_ _11673_/A _09202_/B vssd1 vssd1 vccd1 vccd1 _09203_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_63_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09133_ _09131_/X _09132_/X _09336_/S vssd1 vssd1 vccd1 vccd1 _09133_/X sky130_fd_sc_hd__mux2_1
X_07394_ _07394_/A _07394_/B vssd1 vssd1 vccd1 vccd1 _07401_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_8_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11759__B1 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout220_A _13213_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12264__B _12264_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09064_ _09065_/A _09065_/B _09055_/Y _09073_/C _09073_/A vssd1 vssd1 vccd1 vccd1
+ _09066_/A sky130_fd_sc_hd__o32a_1
XANTENNA__07639__A _12076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10431__B1 _07282_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08015_ _08015_/A _08015_/B vssd1 vssd1 vccd1 vccd1 _08016_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__10065__A _11172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_752 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09966_ _09966_/A vssd1 vssd1 vccd1 vccd1 _09966_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_85_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08917_ _07626_/B _08917_/B vssd1 vssd1 vccd1 vccd1 _08918_/B sky130_fd_sc_hd__and2b_1
X_09897_ _09897_/A _09898_/B vssd1 vssd1 vccd1 vccd1 _09897_/X sky130_fd_sc_hd__or2_1
XFILLER_0_99_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08155__A2 _07752_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08848_ _08848_/A _08848_/B vssd1 vssd1 vccd1 vccd1 _08849_/B sky130_fd_sc_hd__xnor2_4
X_08779_ _08779_/A _08779_/B vssd1 vssd1 vccd1 vccd1 _08780_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__11624__A _11624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11790_ _11790_/A _11822_/B vssd1 vssd1 vccd1 vccd1 _11790_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__07821__B _09614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10810_ _10810_/A _10810_/B vssd1 vssd1 vccd1 vccd1 _10813_/A sky130_fd_sc_hd__xor2_1
XANTENNA__11343__B _11343_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10741_ _10741_/A _10741_/B _10992_/A vssd1 vssd1 vccd1 vccd1 _10741_/X sky130_fd_sc_hd__or3_1
XANTENNA__11462__A2 _12316_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07418__A1 _06612_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12411_ _12287_/A _12287_/B _12382_/Y _12383_/X _12170_/A vssd1 vssd1 vccd1 vccd1
+ _12411_/X sky130_fd_sc_hd__o41a_1
X_10672_ _11470_/A _10672_/B vssd1 vssd1 vccd1 vccd1 _10676_/A sky130_fd_sc_hd__xnor2_1
X_13391_ instruction[6] vssd1 vssd1 vccd1 vccd1 loadstore_size[1] sky130_fd_sc_hd__buf_12
XFILLER_0_23_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12342_ _12423_/A _12342_/B vssd1 vssd1 vccd1 vccd1 _12342_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__08091__B2 _12820_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08091__A1 _12818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12273_ fanout59/X _12215_/S _12216_/Y _12217_/A vssd1 vssd1 vccd1 vccd1 _12275_/B
+ sky130_fd_sc_hd__o22ai_2
XFILLER_0_105_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11224_ _11224_/A _11224_/B vssd1 vssd1 vccd1 vccd1 _11224_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__06929__B1 _06771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11155_ _12261_/A _11155_/B vssd1 vssd1 vccd1 vccd1 _11158_/A sky130_fd_sc_hd__xnor2_1
X_10106_ _10106_/A _10106_/B vssd1 vssd1 vccd1 vccd1 _10106_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_65_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07284__A _09441_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11086_ _11086_/A _11086_/B vssd1 vssd1 vccd1 vccd1 _11088_/C sky130_fd_sc_hd__xnor2_1
X_10037_ fanout29/X _10664_/A _10818_/A fanout27/X vssd1 vssd1 vccd1 vccd1 _10038_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_86_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11988_ _07048_/A fanout6/X _11987_/X _11172_/A vssd1 vssd1 vccd1 vccd1 _12065_/A
+ sky130_fd_sc_hd__a2bb2o_2
X_10939_ _10938_/A _10938_/B _10938_/C vssd1 vssd1 vccd1 vccd1 _10940_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_128_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12609_ reg1_val[25] curr_PC[25] _12622_/S vssd1 vssd1 vccd1 vccd1 _12611_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_54_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13196__A _13214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09820_ _11010_/S _09670_/X _09179_/B vssd1 vssd1 vccd1 vccd1 _09820_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__07042__C1 _12341_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10613__A _10615_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07194__A _07194_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06963_ _06963_/A _07100_/A _07095_/A _07089_/A vssd1 vssd1 vccd1 vccd1 _06967_/C
+ sky130_fd_sc_hd__or4_1
X_09751_ _09751_/A _09751_/B _09751_/C vssd1 vssd1 vccd1 vccd1 _09752_/B sky130_fd_sc_hd__and3_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08702_ _09004_/A _08701_/Y _08703_/A vssd1 vssd1 vccd1 vccd1 _08702_/Y sky130_fd_sc_hd__a21oi_1
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09682_ _10119_/S _09681_/X _09181_/X vssd1 vssd1 vccd1 vccd1 _12299_/B sky130_fd_sc_hd__o21a_1
X_06894_ instruction[11] _06896_/B vssd1 vssd1 vccd1 vccd1 dest_pred[0] sky130_fd_sc_hd__and2_4
XANTENNA_fanout170_A _07192_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08633_ _07026_/A _07026_/B _06574_/Y vssd1 vssd1 vccd1 vccd1 _08635_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_55_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout268_A _06770_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08564_ _08673_/A _08564_/B vssd1 vssd1 vccd1 vccd1 _08565_/B sky130_fd_sc_hd__nor2_1
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07515_ _07515_/A _07515_/B vssd1 vssd1 vccd1 vccd1 _07517_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07648__A1 _08656_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout14 _07345_/Y vssd1 vssd1 vccd1 vccd1 _12854_/A sky130_fd_sc_hd__buf_4
X_08495_ _08495_/A _08495_/B vssd1 vssd1 vccd1 vccd1 _08506_/A sky130_fd_sc_hd__xor2_1
Xfanout25 _09613_/A vssd1 vssd1 vccd1 vccd1 _10574_/A sky130_fd_sc_hd__clkbuf_8
Xfanout47 _12838_/A vssd1 vssd1 vccd1 vccd1 _11847_/A sky130_fd_sc_hd__buf_6
XANTENNA__07648__B2 _08732_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout36 _07282_/B vssd1 vssd1 vccd1 vccd1 fanout36/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_76_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07446_ _07446_/A _07446_/B vssd1 vssd1 vccd1 vccd1 _07449_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_71_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout58 fanout59/X vssd1 vssd1 vccd1 vccd1 _12213_/A sky130_fd_sc_hd__clkbuf_8
Xfanout69 _07072_/X vssd1 vssd1 vccd1 vccd1 fanout69/X sky130_fd_sc_hd__buf_8
XANTENNA__08753__A _11758_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07377_ _07579_/B _07377_/B vssd1 vssd1 vccd1 vccd1 _07395_/A sky130_fd_sc_hd__or2_1
XANTENNA__09568__B _09568_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09116_ reg1_val[8] reg1_val[23] _09142_/S vssd1 vssd1 vccd1 vccd1 _09116_/X sky130_fd_sc_hd__mux2_1
XANTENNA__07369__A _09548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09047_ _09049_/B _09047_/B vssd1 vssd1 vccd1 vccd1 _12031_/C sky130_fd_sc_hd__xor2_2
XANTENNA__07820__A1 _07033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_335 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11619__A _12174_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout83_A _07208_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09949_ _09949_/A _09949_/B vssd1 vssd1 vccd1 vccd1 _10496_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__10183__A2 fanout48/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12960_ hold290/X _13213_/A2 fanout2/X _13213_/B2 vssd1 vssd1 vccd1 vccd1 _12961_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11132__A1 _06981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12891_ hold45/X hold285/X vssd1 vssd1 vccd1 vccd1 _12891_/X sky130_fd_sc_hd__and2b_1
XANTENNA__07887__A1 _07886_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11911_ _11912_/A _11912_/B vssd1 vssd1 vccd1 vccd1 _11992_/B sky130_fd_sc_hd__and2_1
XTAP_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11842_ _11758_/A _11758_/B _11763_/A vssd1 vssd1 vccd1 vccd1 _11846_/A sky130_fd_sc_hd__o21bai_2
XTAP_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11773_ _11824_/A _11773_/B vssd1 vssd1 vccd1 vccd1 _11775_/B sky130_fd_sc_hd__and2_1
XTAP_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10724_ _10724_/A _10724_/B vssd1 vssd1 vccd1 vccd1 _10725_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_70_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10655_ _11707_/A _10623_/Y _10624_/X _10654_/X vssd1 vssd1 vccd1 vccd1 _10655_/X
+ sky130_fd_sc_hd__a31o_1
X_13374_ _13376_/CLK _13374_/D vssd1 vssd1 vccd1 vccd1 hold256/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08064__A1 fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12325_ _12325_/A _12325_/B _12325_/C vssd1 vssd1 vccd1 vccd1 _12326_/B sky130_fd_sc_hd__and3_1
X_10586_ _10586_/A _10586_/B vssd1 vssd1 vccd1 vccd1 _10596_/A sky130_fd_sc_hd__xor2_2
XANTENNA__08064__B2 _08304_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12256_ _06924_/X _12244_/X _12255_/X vssd1 vssd1 vccd1 vccd1 _12256_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_31_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12187_ hold261/A _12187_/B vssd1 vssd1 vccd1 vccd1 _12245_/B sky130_fd_sc_hd__or2_1
XANTENNA__07024__C1 _06960_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11207_ _11207_/A _11207_/B vssd1 vssd1 vccd1 vccd1 _11210_/C sky130_fd_sc_hd__xor2_1
XANTENNA__07218__S _08584_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11138_ _11876_/A _11107_/X _11108_/Y _11137_/X _11106_/Y vssd1 vssd1 vccd1 vccd1
+ _11138_/X sky130_fd_sc_hd__a311o_1
XANTENNA__13112__A2 _06892_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11069_ _11069_/A _11069_/B vssd1 vssd1 vccd1 vccd1 _11070_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_92_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10947__A_N _10448_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07300_ _07300_/A _07300_/B vssd1 vssd1 vccd1 vccd1 _07303_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_46_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08280_ _08280_/A _08280_/B vssd1 vssd1 vccd1 vccd1 _08301_/B sky130_fd_sc_hd__xnor2_2
X_07231_ _07604_/A _07232_/B vssd1 vssd1 vccd1 vccd1 _07231_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_6_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07162_ _09445_/A _07164_/B vssd1 vssd1 vccd1 vccd1 _07167_/A sky130_fd_sc_hd__or2_1
XANTENNA__06805__B _12629_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07093_ _07093_/A _07093_/B vssd1 vssd1 vccd1 vccd1 _07636_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_41_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout204 _09170_/X vssd1 vssd1 vccd1 vccd1 _11968_/B1 sky130_fd_sc_hd__buf_4
XANTENNA__07015__C1 _07064_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12034__S _12388_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08358__A2 _08436_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout237 _06787_/X vssd1 vssd1 vccd1 vccd1 _11231_/S sky130_fd_sc_hd__clkbuf_8
XANTENNA__07128__S _09594_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout215 _06939_/Y vssd1 vssd1 vccd1 vccd1 _11343_/B sky130_fd_sc_hd__buf_6
Xfanout226 _12794_/A vssd1 vssd1 vccd1 vccd1 _08673_/A sky130_fd_sc_hd__buf_4
X_09803_ _09804_/A _09804_/B vssd1 vssd1 vccd1 vccd1 _09803_/X sky130_fd_sc_hd__and2_1
Xfanout248 _11452_/B1 vssd1 vssd1 vccd1 vccd1 _11341_/B sky130_fd_sc_hd__buf_4
Xfanout259 _09442_/A vssd1 vssd1 vccd1 vccd1 _08681_/A sky130_fd_sc_hd__buf_4
X_07995_ _07995_/A _07995_/B vssd1 vssd1 vccd1 vccd1 _07996_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06946_ reg1_val[13] _06946_/B vssd1 vssd1 vccd1 vccd1 _06946_/X sky130_fd_sc_hd__xor2_2
X_09734_ fanout51/X _10589_/A _08507_/B _12214_/A vssd1 vssd1 vccd1 vccd1 _09735_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09858__A2 _10574_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09665_ _09661_/X _09664_/X _11231_/S vssd1 vssd1 vccd1 vccd1 _09665_/X sky130_fd_sc_hd__mux2_1
X_06877_ _09163_/A _06875_/X _09168_/A _06874_/X vssd1 vssd1 vccd1 vccd1 _06877_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11665__A2 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08616_ _08615_/A _08615_/C _08615_/B vssd1 vssd1 vccd1 vccd1 _08621_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_82_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09596_ _09596_/A _09596_/B vssd1 vssd1 vccd1 vccd1 _09597_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_49_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08547_ _08547_/A _08547_/B vssd1 vssd1 vccd1 vccd1 _08549_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_65_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08478_ _09445_/A _08478_/B vssd1 vssd1 vccd1 vccd1 _08508_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_64_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07429_ _10710_/A _07429_/B vssd1 vssd1 vccd1 vccd1 _07433_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_80_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07099__A _07099_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10440_ _10440_/A _10440_/B vssd1 vssd1 vccd1 vccd1 _10441_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_18_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09243__B1 _09593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08597__A2 _08727_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10371_ _10741_/B _10371_/B vssd1 vssd1 vccd1 vccd1 _10658_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__11050__B1 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13090_ _06572_/A hold302/X _13089_/X _06892_/B hold260/X vssd1 vssd1 vccd1 vccd1
+ hold303/A sky130_fd_sc_hd__a32o_1
X_12110_ _12110_/A _12110_/B vssd1 vssd1 vccd1 vccd1 _12110_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__07827__A _11385_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold280 hold280/A vssd1 vssd1 vccd1 vccd1 hold280/X sky130_fd_sc_hd__dlygate4sd3_1
X_12041_ _12041_/A _12041_/B vssd1 vssd1 vccd1 vccd1 _12041_/Y sky130_fd_sc_hd__xnor2_1
Xhold291 hold291/A vssd1 vssd1 vccd1 vccd1 hold291/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11353__A1 _11876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10156__A2 _10818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09761__B _09761_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12943_ _12874_/X _12943_/B vssd1 vssd1 vccd1 vccd1 _13193_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_99_132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12874_ hold3/X hold252/X vssd1 vssd1 vccd1 vccd1 _12874_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_62_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11825_ _11747_/Y _11750_/B _11746_/A vssd1 vssd1 vccd1 vccd1 _11833_/A sky130_fd_sc_hd__o21a_1
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08393__A _08645_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11756_ fanout24/X fanout56/X _12316_/A _07819_/B vssd1 vssd1 vccd1 vccd1 _11757_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_28_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10707_ _10707_/A _10707_/B vssd1 vssd1 vccd1 vccd1 _10712_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_126_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11687_ _11687_/A _11687_/B _11687_/C vssd1 vssd1 vccd1 vccd1 _11688_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_125_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10638_ _09966_/Y _10637_/X _11233_/S vssd1 vssd1 vccd1 vccd1 _10638_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_3_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10919__B2 _10575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10919__A1 _10574_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13357_ _13357_/CLK _13357_/D vssd1 vssd1 vccd1 vccd1 hold269/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10569_ _10569_/A _10569_/B vssd1 vssd1 vccd1 vccd1 _10585_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_3_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11041__B1 fanout12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13288_ _13311_/CLK _13288_/D vssd1 vssd1 vccd1 vccd1 hold185/A sky130_fd_sc_hd__dfxtp_1
X_12308_ _06625_/X _11973_/B _12307_/Y _06627_/B _12404_/A vssd1 vssd1 vccd1 vccd1
+ _12308_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_87_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07737__A _08722_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07260__A2 _07263_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07796__B1 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12239_ _12185_/A _12182_/Y _12184_/B vssd1 vssd1 vccd1 vccd1 _12243_/A sky130_fd_sc_hd__o21a_1
XANTENNA__11259__A _11908_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11895__A2 _09527_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06800_ _06805_/A _06702_/A _12634_/B _06799_/X vssd1 vssd1 vccd1 vccd1 _06800_/Y
+ sky130_fd_sc_hd__a31oi_2
X_07780_ _07781_/B _07781_/C _07781_/A vssd1 vssd1 vccd1 vccd1 _07782_/A sky130_fd_sc_hd__a21oi_1
X_06731_ _10897_/S _06731_/B vssd1 vssd1 vccd1 vccd1 _10879_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_36_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09450_ _11384_/A _09450_/B vssd1 vssd1 vccd1 vccd1 _09452_/B sky130_fd_sc_hd__xnor2_1
X_06662_ _11894_/A _06662_/B vssd1 vssd1 vccd1 vccd1 _11880_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_59_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08401_ _10444_/A _08401_/B vssd1 vssd1 vccd1 vccd1 _08405_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07720__B1 _11766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12818__A _12818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06593_ instruction[41] _06897_/B _06591_/X vssd1 vssd1 vccd1 vccd1 _06771_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_93_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09381_ _09548_/A _09381_/B vssd1 vssd1 vccd1 vccd1 _09385_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11804__C1 _06924_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07079__A2 _06960_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08276__A1 _08723_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08276__B2 _07885_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08332_ _08332_/A _08332_/B vssd1 vssd1 vccd1 vccd1 _08383_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08263_ _08730_/A1 _08732_/A1 _08038_/A _08741_/B2 vssd1 vssd1 vccd1 vccd1 _08264_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout133_A _09238_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07214_ _07214_/A _07214_/B vssd1 vssd1 vccd1 vccd1 _07230_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_27_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08194_ _08724_/A _08194_/B vssd1 vssd1 vccd1 vccd1 _08197_/B sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout300_A _13242_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08579__A2 _08661_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07145_ _07141_/X _07144_/X _07151_/B _07144_/A vssd1 vssd1 vccd1 vccd1 _07145_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_42_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07787__B1 _08564_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07076_ _11164_/A _07076_/B vssd1 vssd1 vccd1 vccd1 _07076_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_0_112_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07366__B _07508_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07978_ _07978_/A _07978_/B vssd1 vssd1 vccd1 vccd1 _08024_/B sky130_fd_sc_hd__xnor2_1
X_06929_ instruction[17] _06924_/X _09152_/B _06771_/A vssd1 vssd1 vccd1 vccd1 _06929_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__08478__A _09445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09717_ _09718_/A _09718_/B vssd1 vssd1 vccd1 vccd1 _09719_/A sky130_fd_sc_hd__or2_2
X_09648_ _09953_/A _09953_/B vssd1 vssd1 vccd1 vccd1 _09648_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_69_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12048__C1 _12247_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09579_ _10445_/A _11847_/A _10570_/B _10706_/B2 vssd1 vssd1 vccd1 vccd1 _09580_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12590_ reg1_val[22] curr_PC[22] _12622_/S vssd1 vssd1 vccd1 vccd1 _12592_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_77_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08267__A1 _12818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08267__B2 _12820_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11610_ _11214_/X _11609_/A _11607_/Y vssd1 vssd1 vccd1 vccd1 _11610_/Y sky130_fd_sc_hd__a21oi_1
X_11541_ _11540_/A _09527_/B _11540_/Y _12307_/B1 vssd1 vssd1 vccd1 vccd1 _11541_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_80_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11472_ _11472_/A _12214_/B vssd1 vssd1 vccd1 vccd1 _11473_/B sky130_fd_sc_hd__nor2_1
X_13211_ _13211_/A _13211_/B vssd1 vssd1 vccd1 vccd1 _13211_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__12463__A _12639_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09767__A1 _09594_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10423_ _10424_/A _10424_/B _10424_/C vssd1 vssd1 vccd1 vccd1 _10423_/Y sky130_fd_sc_hd__a21oi_1
X_13142_ hold285/X _12789_/B _13141_/X _12790_/A vssd1 vssd1 vccd1 vccd1 hold286/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10354_ _10221_/A _10221_/B _10219_/X vssd1 vssd1 vccd1 vccd1 _10356_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_20_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13073_ _11987_/B _13077_/A2 hold108/X vssd1 vssd1 vccd1 vccd1 _13339_/D sky130_fd_sc_hd__o21a_1
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10285_ _10285_/A _10285_/B vssd1 vssd1 vccd1 vccd1 _10288_/A sky130_fd_sc_hd__nor2_1
X_12024_ _12165_/A _12024_/B _12165_/B vssd1 vssd1 vccd1 vccd1 _12025_/A sky130_fd_sc_hd__or3_1
XANTENNA__13079__A1 _07522_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07950__B1 _08721_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12926_ _13129_/B _13130_/A _12897_/X vssd1 vssd1 vccd1 vccd1 _13135_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_87_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12857_ _12412_/A _13087_/B2 hold87/X _13235_/A vssd1 vssd1 vccd1 vccd1 _13282_/D
+ sky130_fd_sc_hd__o211a_1
X_11808_ hold275/A _11808_/B vssd1 vssd1 vccd1 vccd1 _11888_/B sky130_fd_sc_hd__or2_1
XFILLER_0_68_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08258__A1 _08752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12788_ _12788_/A hold168/X vssd1 vssd1 vccd1 vccd1 _12789_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_113_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08258__B2 _08798_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11739_ _11689_/A _11689_/B _11688_/A vssd1 vssd1 vccd1 vccd1 _11779_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_22_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09947__A _09949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11565__A1 _11653_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11565__B2 _08752_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10773__C1 _10772_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08430__B2 _08646_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08430__A1 _08798_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08950_ _08950_/A _08950_/B vssd1 vssd1 vccd1 vccd1 _08951_/B sky130_fd_sc_hd__xor2_4
XANTENNA__10525__C1 _06881_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08881_ _08882_/A _08882_/B vssd1 vssd1 vccd1 vccd1 _08898_/B sky130_fd_sc_hd__nand2_1
X_07901_ _07911_/A _07911_/B _07911_/C vssd1 vssd1 vccd1 vccd1 _07913_/A sky130_fd_sc_hd__a21o_1
XANTENNA__12820__B _12830_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07832_ _07896_/A _09609_/B _09396_/B _08723_/B1 vssd1 vssd1 vccd1 vccd1 _07833_/B
+ sky130_fd_sc_hd__o22a_1
X_09502_ _09105_/X _09109_/X _09663_/S vssd1 vssd1 vccd1 vccd1 _09502_/X sky130_fd_sc_hd__mux2_1
X_07763_ _08732_/A1 fanout87/X fanout82/X _10927_/A1 vssd1 vssd1 vccd1 vccd1 _07764_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09694__B1 _09354_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06714_ reg2_val[14] _06799_/B vssd1 vssd1 vccd1 vccd1 _06714_/X sky130_fd_sc_hd__and2_1
X_07694_ _07695_/B _07694_/B vssd1 vssd1 vccd1 vccd1 _07986_/B sky130_fd_sc_hd__and2b_1
XANTENNA_fanout250_A _12247_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06645_ reg1_val[24] _07166_/A vssd1 vssd1 vccd1 vccd1 _06646_/B sky130_fd_sc_hd__or2_1
X_09433_ _09433_/A _09433_/B vssd1 vssd1 vccd1 vccd1 _09435_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__12548__A _12703_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09364_ _09364_/A _09364_/B vssd1 vssd1 vccd1 vccd1 _09364_/Y sky130_fd_sc_hd__xnor2_1
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06576_ reg1_val[29] vssd1 vssd1 vccd1 vccd1 _06838_/A sky130_fd_sc_hd__inv_2
XFILLER_0_74_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08315_ _08315_/A _08315_/B vssd1 vssd1 vccd1 vccd1 _08371_/B sky130_fd_sc_hd__xor2_2
XANTENNA__11171__B _11923_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_31 reg2_val[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_20 reg2_val[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09295_ _09296_/B _09296_/A vssd1 vssd1 vccd1 vccd1 _09295_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_47_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_42 pred_val vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_64 reg1_val[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07472__A2 _08507_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_53 reg1_val[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08246_ _08246_/A _08246_/B vssd1 vssd1 vccd1 vccd1 _08296_/B sky130_fd_sc_hd__and2_1
XFILLER_0_104_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08177_ _08215_/A _08215_/B vssd1 vssd1 vccd1 vccd1 _08240_/A sky130_fd_sc_hd__nor2_1
X_07128_ _07139_/A _07139_/B _09594_/A vssd1 vssd1 vccd1 vccd1 _07128_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_30_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07224__A2 _07220_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07059_ reg1_val[16] _07254_/B _07364_/B1 reg1_val[17] vssd1 vssd1 vccd1 vccd1 _07071_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_100_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09592__A _09593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10070_ _10070_/A _10070_/B vssd1 vssd1 vccd1 vccd1 _10073_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_10_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08185__B1 _08617_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10972_ _10821_/A _10821_/B _10819_/Y vssd1 vssd1 vccd1 vccd1 _10974_/B sky130_fd_sc_hd__a21boi_1
X_12711_ _12712_/A _12712_/B vssd1 vssd1 vccd1 vccd1 _12725_/A sky130_fd_sc_hd__or2_1
XANTENNA__10295__B2 _10706_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10295__A1 _10445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12642_ _12641_/A _12638_/Y _12640_/B vssd1 vssd1 vccd1 vccd1 _12646_/A sky130_fd_sc_hd__o21a_2
XANTENNA__11244__A0 _09527_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12573_ _12623_/A _12573_/B vssd1 vssd1 vccd1 vccd1 _12574_/B sky130_fd_sc_hd__or2_1
XFILLER_0_65_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11524_ _12174_/S _11524_/B vssd1 vssd1 vccd1 vccd1 _11524_/X sky130_fd_sc_hd__or2_1
XFILLER_0_80_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07463__A2 fanout66/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11455_ _11968_/B1 _11450_/X _11451_/Y _11454_/X vssd1 vssd1 vccd1 vccd1 _11455_/X
+ sky130_fd_sc_hd__o31a_1
XANTENNA__06903__B _06921_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10406_ _11142_/S _10402_/X _10405_/X vssd1 vssd1 vccd1 vccd1 dest_val[8] sky130_fd_sc_hd__o21ai_4
XFILLER_0_61_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11386_ _09609_/B fanout12/X fanout8/X _09396_/B vssd1 vssd1 vccd1 vccd1 _11387_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_0_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13125_ _13125_/A _13125_/B vssd1 vssd1 vccd1 vccd1 _13125_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_103_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06974__A1 _10445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10337_ _10338_/A _10338_/B vssd1 vssd1 vccd1 vccd1 _10454_/B sky130_fd_sc_hd__and2_1
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10268_ _12244_/S _09172_/B _10267_/Y _10262_/Y vssd1 vssd1 vccd1 vccd1 _10268_/X
+ sky130_fd_sc_hd__a31o_1
X_13056_ hold76/X _12791_/A _13080_/B1 _13331_/Q _13128_/A vssd1 vssd1 vccd1 vccd1
+ hold77/A sky130_fd_sc_hd__o221a_1
XANTENNA__06974__B2 _10418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12007_ _12009_/A _12009_/B vssd1 vssd1 vccd1 vccd1 _12010_/A sky130_fd_sc_hd__and2_1
XFILLER_0_84_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10199_ _11294_/A _10574_/A _10575_/A _10418_/A vssd1 vssd1 vccd1 vccd1 _10200_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_17_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11256__B _11650_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_76 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12909_ hold284/X hold49/X vssd1 vssd1 vccd1 vccd1 _12910_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__07750__A _08728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10286__A1 _10571_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10286__B2 _10570_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09691__A3 hold260/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09080_ _09165_/A _09170_/A vssd1 vssd1 vccd1 vccd1 _11707_/A sky130_fd_sc_hd__nor2_4
X_08100_ _08728_/A _08100_/B vssd1 vssd1 vccd1 vccd1 _08108_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_71_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08031_ _08031_/A _08031_/B _08031_/C vssd1 vssd1 vccd1 vccd1 _08034_/A sky130_fd_sc_hd__and3_1
XANTENNA__09396__B _09396_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09600__B1 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08403__B2 _08798_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08403__A1 _08673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09982_ hold258/A _09983_/B vssd1 vssd1 vccd1 vccd1 _09982_/X sky130_fd_sc_hd__and2_1
X_08933_ _08934_/B _08934_/A vssd1 vssd1 vccd1 vccd1 _08933_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__07925__A _08745_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout298_A _13242_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09903__A1 _12214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12042__S _12244_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09903__B2 fanout59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08864_ _08864_/A _08864_/B vssd1 vssd1 vccd1 vccd1 _08865_/B sky130_fd_sc_hd__or2_2
X_07815_ _07814_/A _07814_/B _07813_/X vssd1 vssd1 vccd1 vccd1 _07816_/C sky130_fd_sc_hd__o21bai_1
X_08795_ _08795_/A _08795_/B vssd1 vssd1 vccd1 vccd1 _08817_/A sky130_fd_sc_hd__xnor2_1
X_07746_ _07746_/A _07746_/B vssd1 vssd1 vccd1 vccd1 _07784_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_67_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07660__A _10165_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09416_ _09274_/B _09277_/B _09272_/X vssd1 vssd1 vccd1 vccd1 _09418_/B sky130_fd_sc_hd__a21oi_2
X_07677_ _08942_/A _08942_/B _07676_/A vssd1 vssd1 vccd1 vccd1 _08959_/A sky130_fd_sc_hd__a21o_1
X_06628_ instruction[35] _06634_/B vssd1 vssd1 vccd1 vccd1 _12673_/B sky130_fd_sc_hd__and2_4
XFILLER_0_94_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09347_ _12254_/A1 _09346_/X _09341_/Y vssd1 vssd1 vccd1 vccd1 _09347_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_75_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09278_ _09351_/B _12264_/B _07515_/B _07513_/X vssd1 vssd1 vccd1 vccd1 _09280_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_35_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11910__A _12073_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08229_ _08740_/A _08229_/B vssd1 vssd1 vccd1 vccd1 _08235_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_7_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06723__B _11020_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07819__B _07819_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11240_ hold279/A _11240_/B vssd1 vssd1 vccd1 vccd1 _11339_/B sky130_fd_sc_hd__or2_1
XFILLER_0_120_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11171_ _11171_/A _11923_/A vssd1 vssd1 vccd1 vccd1 _11172_/C sky130_fd_sc_hd__or2_1
XANTENNA__10201__B2 _10571_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10201__A1 _10570_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10122_ hold157/A _10391_/A2 _10253_/B _12401_/B1 vssd1 vssd1 vccd1 vccd1 _10123_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_100_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10053_ _10054_/A _10054_/B vssd1 vssd1 vccd1 vccd1 _10174_/A sky130_fd_sc_hd__and2_1
XFILLER_0_98_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10268__A1 _12244_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10955_ _10956_/A _10956_/B vssd1 vssd1 vccd1 vccd1 _10957_/A sky130_fd_sc_hd__nand2_1
X_10886_ _10755_/X _10759_/A _10884_/X _10885_/Y vssd1 vssd1 vccd1 vccd1 _10888_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_57_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12625_ _12626_/A _12626_/B vssd1 vssd1 vccd1 vccd1 _12631_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_26_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12916__A hold260/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12556_ _12556_/A _12556_/B _12556_/C vssd1 vssd1 vccd1 vccd1 _12557_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_5_419 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11507_ _11508_/A _11508_/B _11508_/C vssd1 vssd1 vccd1 vccd1 _11507_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_124_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12487_ _12488_/A _12488_/B _12488_/C vssd1 vssd1 vccd1 vccd1 _12495_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_80_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold109 hold109/A vssd1 vssd1 vccd1 vccd1 hold109/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11438_ _11337_/A _11334_/Y _11336_/B vssd1 vssd1 vccd1 vccd1 _11442_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_1_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11369_ _11369_/A _11369_/B vssd1 vssd1 vccd1 vccd1 _11370_/B sky130_fd_sc_hd__and2_1
X_13108_ hold291/X _06892_/B _13107_/X _06572_/A vssd1 vssd1 vccd1 vccd1 _13109_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13039_ _10165_/A _12798_/B hold156/X vssd1 vssd1 vccd1 vccd1 _13322_/D sky130_fd_sc_hd__a21boi_1
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08580_ _08728_/A _08580_/B vssd1 vssd1 vccd1 vccd1 _08612_/A sky130_fd_sc_hd__xnor2_1
X_07600_ _07600_/A _07600_/B vssd1 vssd1 vccd1 vccd1 _07681_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__07480__A _10449_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07531_ _07099_/A _07099_/B _10963_/A vssd1 vssd1 vccd1 vccd1 _07533_/B sky130_fd_sc_hd__a21o_1
XANTENNA__07124__A1 _12626_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06808__B _09351_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07462_ _09746_/A _07462_/B vssd1 vssd1 vccd1 vccd1 _07568_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_119_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09201_ fanout30/X _09768_/A1 _12808_/A _07688_/B vssd1 vssd1 vccd1 vccd1 _09202_/B
+ sky130_fd_sc_hd__o22a_1
X_07393_ _07393_/A _07393_/B vssd1 vssd1 vccd1 vccd1 _07394_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_8_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12826__A _12826_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09132_ _09343_/A reg1_val[30] _09142_/S vssd1 vssd1 vccd1 vccd1 _09132_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_72_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11759__A1 _09613_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11759__B2 _09614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10431__A1 _10818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09063_ _09065_/A _09065_/B vssd1 vssd1 vccd1 vccd1 _09063_/X sky130_fd_sc_hd__or2_1
XANTENNA__10431__B2 _10963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08014_ _08013_/A _08013_/B _08015_/A vssd1 vssd1 vccd1 vccd1 _08014_/X sky130_fd_sc_hd__o21a_1
XANTENNA__08388__B1 _09440_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09965_ _11010_/S _09509_/X _09179_/B vssd1 vssd1 vccd1 vccd1 _09966_/A sky130_fd_sc_hd__o21ai_1
X_08916_ _08916_/A _08916_/B vssd1 vssd1 vccd1 vccd1 _08922_/A sky130_fd_sc_hd__xnor2_1
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09896_ _10449_/A _09896_/B vssd1 vssd1 vccd1 vccd1 _09898_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_85_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08847_ _08847_/A _08847_/B vssd1 vssd1 vccd1 vccd1 _08849_/A sky130_fd_sc_hd__nor2_2
X_08778_ _08778_/A _08778_/B vssd1 vssd1 vccd1 vccd1 _08779_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__06718__B _06981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07729_ _07729_/A _07729_/B vssd1 vssd1 vccd1 vccd1 _07730_/B sky130_fd_sc_hd__and2_1
XANTENNA__08312__B1 _08727_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10740_ _10494_/X _10992_/A _10738_/X vssd1 vssd1 vccd1 vccd1 _10740_/X sky130_fd_sc_hd__o21a_1
XANTENNA__06722__A_N _11020_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10671_ _10941_/A _12150_/A _12213_/A fanout94/X vssd1 vssd1 vccd1 vccd1 _10672_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_125_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12410_ _06612_/B _06939_/Y _12386_/X _12409_/X _12455_/S vssd1 vssd1 vccd1 vccd1
+ dest_val[30] sky130_fd_sc_hd__o221a_4
XFILLER_0_48_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13390_ instruction[5] vssd1 vssd1 vccd1 vccd1 loadstore_size[0] sky130_fd_sc_hd__buf_12
XFILLER_0_35_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12341_ _12341_/A _12341_/B vssd1 vssd1 vccd1 vccd1 _12341_/X sky130_fd_sc_hd__or2_1
XFILLER_0_62_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08091__A2 _08741_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12272_ _12327_/A _12272_/B vssd1 vssd1 vccd1 vccd1 _12275_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_16_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11223_ _06822_/X _11222_/X _12174_/S vssd1 vssd1 vccd1 vccd1 _11224_/B sky130_fd_sc_hd__mux2_1
XANTENNA__12471__A _12644_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11154_ _10418_/A fanout9/X fanout4/X _11294_/A vssd1 vssd1 vccd1 vccd1 _11155_/B
+ sky130_fd_sc_hd__o22a_1
X_10105_ _10748_/A _10105_/B vssd1 vssd1 vccd1 vccd1 _10106_/B sky130_fd_sc_hd__nor2_1
XANTENNA__09879__B1 _10574_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11085_ _11085_/A _11085_/B vssd1 vssd1 vccd1 vccd1 _11086_/B sky130_fd_sc_hd__xnor2_1
X_10036_ _10959_/A _10036_/B _10036_/C vssd1 vssd1 vccd1 vccd1 _10040_/B sky130_fd_sc_hd__or3_1
XANTENNA__09780__A _11261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08396__A _08598_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11987_ _11987_/A _11987_/B fanout6/X vssd1 vssd1 vccd1 vccd1 _11987_/X sky130_fd_sc_hd__or3_1
XFILLER_0_105_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10110__B1 _09156_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10938_ _10938_/A _10938_/B _10938_/C vssd1 vssd1 vccd1 vccd1 _11076_/B sky130_fd_sc_hd__and3_1
XFILLER_0_105_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10869_ _10870_/B _10870_/C _10870_/D _11100_/A vssd1 vssd1 vccd1 vccd1 _10871_/A
+ sky130_fd_sc_hd__a31o_1
X_12608_ _12608_/A _12608_/B vssd1 vssd1 vccd1 vccd1 new_PC[24] sky130_fd_sc_hd__xor2_4
XANTENNA__13060__C1 _13128_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12539_ reg1_val[14] curr_PC[14] _12622_/S vssd1 vssd1 vccd1 vccd1 _12541_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_54_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07042__B1 _07064_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07475__A _10165_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06962_ _06964_/A _06964_/B vssd1 vssd1 vccd1 vccd1 _07133_/A sky130_fd_sc_hd__or2_1
X_09750_ _09751_/A _09751_/B _09751_/C vssd1 vssd1 vccd1 vccd1 _09752_/A sky130_fd_sc_hd__a21oi_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09681_ _11010_/S _09680_/X _09179_/B vssd1 vssd1 vccd1 vccd1 _09681_/X sky130_fd_sc_hd__o21a_1
X_08701_ _08571_/A _08571_/B _08571_/C vssd1 vssd1 vccd1 vccd1 _08701_/Y sky130_fd_sc_hd__o21ai_1
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06893_ instruction[2] instruction[1] pred_val instruction[0] vssd1 vssd1 vccd1 vccd1
+ _06896_/B sky130_fd_sc_hd__and4b_4
X_08632_ _08632_/A _08632_/B _08632_/C vssd1 vssd1 vccd1 vccd1 _08635_/B sky130_fd_sc_hd__nand3_1
XANTENNA_fanout163_A _08979_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08563_ _08742_/A _08563_/B vssd1 vssd1 vccd1 vccd1 _08591_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_77_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11429__B1 _12290_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07514_ _07514_/A _07514_/B vssd1 vssd1 vccd1 vccd1 _07515_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_76_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08494_ _08494_/A _08494_/B vssd1 vssd1 vccd1 vccd1 _08517_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__07648__A2 _11847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07445_ _07445_/A _07445_/B vssd1 vssd1 vccd1 vccd1 _07446_/B sky130_fd_sc_hd__nand2_1
Xfanout37 _07263_/Y vssd1 vssd1 vccd1 vccd1 _07282_/B sky130_fd_sc_hd__buf_8
Xfanout26 _07033_/X vssd1 vssd1 vccd1 vccd1 _09613_/A sky130_fd_sc_hd__clkbuf_8
Xfanout15 fanout16/X vssd1 vssd1 vccd1 vccd1 fanout15/X sky130_fd_sc_hd__buf_6
XANTENNA__13151__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout59 _12848_/A vssd1 vssd1 vccd1 vccd1 fanout59/X sky130_fd_sc_hd__clkbuf_8
Xfanout48 _12838_/A vssd1 vssd1 vccd1 vccd1 fanout48/X sky130_fd_sc_hd__clkbuf_8
X_07376_ _07376_/A _07376_/B _07376_/C vssd1 vssd1 vccd1 vccd1 _07377_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09115_ _09099_/X _09114_/X _11231_/S vssd1 vssd1 vccd1 vccd1 _09115_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_60_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09046_ _11793_/A _11875_/A _11953_/A _11792_/B vssd1 vssd1 vccd1 vccd1 _12031_/B
+ sky130_fd_sc_hd__and4bb_2
XFILLER_0_32_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07820__A2 _07033_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09948_ _09949_/A _09949_/B vssd1 vssd1 vccd1 vccd1 _09948_/X sky130_fd_sc_hd__and2_1
XANTENNA_fanout76_A _09548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11132__A2 _12404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08533__B1 _08617_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09879_ _09609_/B _09745_/B _10574_/B _09396_/B vssd1 vssd1 vccd1 vccd1 _09880_/B
+ sky130_fd_sc_hd__o22a_1
X_12890_ hold287/A hold43/X vssd1 vssd1 vccd1 vccd1 _13149_/B sky130_fd_sc_hd__nand2b_1
X_11910_ _12073_/A _11910_/B vssd1 vssd1 vccd1 vccd1 _11912_/B sky130_fd_sc_hd__xnor2_1
XTAP_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11841_ _11755_/B _11764_/B _11753_/A vssd1 vssd1 vccd1 vccd1 _11854_/A sky130_fd_sc_hd__o21a_1
XTAP_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11772_ _11772_/A _11772_/B _11772_/C vssd1 vssd1 vccd1 vccd1 _11773_/B sky130_fd_sc_hd__or3_1
XTAP_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10723_ _10722_/A _10722_/B _10724_/A vssd1 vssd1 vccd1 vccd1 _10723_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_27_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10654_ _11876_/A _10625_/X _10626_/Y _10653_/X vssd1 vssd1 vccd1 vccd1 _10654_/X
+ sky130_fd_sc_hd__a31o_1
X_13373_ _13376_/CLK _13373_/D vssd1 vssd1 vccd1 vccd1 hold281/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10585_ _10585_/A _10585_/B vssd1 vssd1 vccd1 vccd1 _10586_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__08064__A2 _08723_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12324_ _12325_/A _12325_/B _12325_/C vssd1 vssd1 vccd1 vccd1 _12373_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_35_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06911__B _06921_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12255_ _12249_/Y _12250_/X _12254_/X _12247_/X vssd1 vssd1 vccd1 vccd1 _12255_/X
+ sky130_fd_sc_hd__o211a_1
X_12186_ _09968_/A _12185_/Y _12429_/B vssd1 vssd1 vccd1 vccd1 _12186_/X sky130_fd_sc_hd__mux2_1
X_11206_ _11207_/B _11207_/A vssd1 vssd1 vccd1 vccd1 _11315_/B sky130_fd_sc_hd__nand2b_1
X_11137_ _11137_/A _11137_/B _11136_/X vssd1 vssd1 vccd1 vccd1 _11137_/X sky130_fd_sc_hd__or3b_1
XFILLER_0_92_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08524__B1 _08038_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11659__B1 fanout4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11068_ _11069_/A _11069_/B vssd1 vssd1 vccd1 vccd1 _11068_/X sky130_fd_sc_hd__and2b_1
X_10019_ _10019_/A _10019_/B vssd1 vssd1 vccd1 vccd1 _10021_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__10331__B1 _10963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07230_ _07230_/A _07230_/B vssd1 vssd1 vccd1 vccd1 _07232_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_41_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07161_ reg1_val[4] _07161_/B vssd1 vssd1 vccd1 vccd1 _07164_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_54_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07092_ _11261_/A _07092_/B vssd1 vssd1 vccd1 vccd1 _07093_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_41_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout205 _09170_/X vssd1 vssd1 vccd1 vccd1 _12401_/B1 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07015__B1 _12341_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout227 _09336_/S vssd1 vssd1 vccd1 vccd1 _09330_/S sky130_fd_sc_hd__clkbuf_8
Xfanout216 _06923_/Y vssd1 vssd1 vccd1 vccd1 _09172_/B sky130_fd_sc_hd__clkbuf_8
X_09802_ _09802_/A _09802_/B vssd1 vssd1 vccd1 vccd1 _09804_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_10_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout249 _09355_/X vssd1 vssd1 vccd1 vccd1 _11452_/B1 sky130_fd_sc_hd__clkbuf_4
X_07994_ _07994_/A vssd1 vssd1 vccd1 vccd1 _07996_/A sky130_fd_sc_hd__inv_2
XANTENNA_fanout280_A hold65/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06945_ _07200_/A _06994_/D vssd1 vssd1 vccd1 vccd1 _06946_/B sky130_fd_sc_hd__nand2_1
X_09733_ _09869_/B _09733_/B vssd1 vssd1 vccd1 vccd1 _09775_/A sky130_fd_sc_hd__or2_1
XANTENNA__13146__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09664_ _09662_/X _09663_/X _09974_/A vssd1 vssd1 vccd1 vccd1 _09664_/X sky130_fd_sc_hd__mux2_1
X_06876_ instruction[3] instruction[4] vssd1 vssd1 vccd1 vccd1 _09168_/A sky130_fd_sc_hd__nand2_2
X_08615_ _08615_/A _08615_/B _08615_/C vssd1 vssd1 vccd1 vccd1 _08621_/A sky130_fd_sc_hd__and3_1
X_09595_ _09596_/A _09596_/B vssd1 vssd1 vccd1 vccd1 _09595_/Y sky130_fd_sc_hd__nor2_1
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08546_ _08546_/A _08546_/B vssd1 vssd1 vccd1 vccd1 _08547_/B sky130_fd_sc_hd__and2_1
XANTENNA__12075__B1 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08477_ _07885_/B _08661_/A2 _08673_/B _08721_/B1 vssd1 vssd1 vccd1 vccd1 _08478_/B
+ sky130_fd_sc_hd__o22a_1
X_07428_ _10589_/A _12834_/A _12836_/A _08507_/B vssd1 vssd1 vccd1 vccd1 _07429_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_18_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07359_ _11163_/A _07359_/B vssd1 vssd1 vccd1 vccd1 _07360_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__07099__B _07099_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_442 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11050__A1 _10570_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10370_ _09810_/B _10368_/X _10369_/X _10864_/A vssd1 vssd1 vccd1 vccd1 _10371_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_5_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11050__B2 _10571_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09029_ _11521_/B _11521_/C vssd1 vssd1 vccd1 vccd1 _11616_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_20_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold270 hold270/A vssd1 vssd1 vccd1 vccd1 hold270/X sky130_fd_sc_hd__dlygate4sd3_1
X_12040_ _12038_/Y _12040_/B vssd1 vssd1 vccd1 vccd1 _12041_/B sky130_fd_sc_hd__and2b_1
Xhold292 hold292/A vssd1 vssd1 vccd1 vccd1 hold292/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold281 hold281/A vssd1 vssd1 vccd1 vccd1 hold281/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_4_12_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11105__A2 _11650_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12942_ hold252/X hold3/X vssd1 vssd1 vccd1 vccd1 _12943_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_87_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12873_ hold246/X hold1/X vssd1 vssd1 vccd1 vccd1 _13197_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_68_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08674__A _09445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11824_ _11824_/A _11824_/B vssd1 vssd1 vccd1 vccd1 _11859_/A sky130_fd_sc_hd__nand2_1
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11813__B1 _12254_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10709__A _11163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11755_ _11755_/A _11755_/B vssd1 vssd1 vccd1 vccd1 _11764_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_28_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07493__B1 _12854_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10706_ _10445_/A fanout13/X fanout6/X _10706_/B2 vssd1 vssd1 vccd1 vccd1 _10707_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_126_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12369__A1 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11686_ _11687_/A _11687_/B _11687_/C vssd1 vssd1 vccd1 vccd1 _11688_/A sky130_fd_sc_hd__a21o_1
XANTENNA__13030__A2 _06572_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10637_ _09503_/X _09507_/X _11010_/S vssd1 vssd1 vccd1 vccd1 _10637_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_36_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10919__A2 fanout48/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13356_ _13357_/CLK _13356_/D vssd1 vssd1 vccd1 vccd1 hold288/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07796__A1 _12820_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10568_ _10567_/A _10959_/A _10569_/A vssd1 vssd1 vccd1 vccd1 _10568_/X sky130_fd_sc_hd__and3b_1
XANTENNA__11041__B2 fanout94/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11041__A1 _10941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12643__B _12644_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13287_ _13311_/CLK _13287_/D vssd1 vssd1 vccd1 vccd1 hold187/A sky130_fd_sc_hd__dfxtp_1
X_12307_ _06625_/X _12402_/A0 _12307_/B1 vssd1 vssd1 vccd1 vccd1 _12307_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__10658__C_N _10500_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10499_ _10499_/A _10499_/B _10499_/C vssd1 vssd1 vccd1 vccd1 _10500_/B sky130_fd_sc_hd__and3_1
XANTENNA__07796__B2 _08741_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10444__A _10444_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06641__B _12669_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12238_ _12238_/A _12238_/B vssd1 vssd1 vccd1 vccd1 _12238_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__11344__A2 _11973_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12169_ _12169_/A _12169_/B _12169_/C _12169_/D vssd1 vssd1 vccd1 vccd1 _12287_/A
+ sky130_fd_sc_hd__or4_4
XANTENNA__10552__B1 _07282_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07753__A _11908_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06730_ reg1_val[12] _07074_/A vssd1 vssd1 vccd1 vccd1 _06731_/B sky130_fd_sc_hd__nor2_1
X_06661_ reg1_val[22] _07191_/A vssd1 vssd1 vccd1 vccd1 _06662_/B sky130_fd_sc_hd__nor2_1
X_08400_ _07821_/A fanout87/X fanout82/X _09423_/B2 vssd1 vssd1 vccd1 vccd1 _08401_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07720__B2 _08656_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07720__A1 _08732_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06592_ instruction[1] instruction[2] instruction[25] pred_val vssd1 vssd1 vccd1
+ vccd1 _06592_/Y sky130_fd_sc_hd__o211ai_1
XANTENNA__08584__A _08584_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09380_ _12804_/A fanout16/X _07282_/B _09768_/A1 vssd1 vssd1 vccd1 vccd1 _09381_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_59_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12818__B _12818_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07079__A3 _09147_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08331_ _08331_/A _08331_/B vssd1 vssd1 vccd1 vccd1 _08383_/A sky130_fd_sc_hd__xor2_1
XANTENNA__08276__A2 _08744_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07484__B1 _07076_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08262_ _08733_/A _08262_/B vssd1 vssd1 vccd1 vccd1 _08266_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_117_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07213_ _07214_/A _07214_/B vssd1 vssd1 vccd1 vccd1 _07376_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_62_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12834__A _12834_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08193_ fanout75/X _07821_/A _07752_/B _08304_/B vssd1 vssd1 vccd1 vccd1 _08194_/B
+ sky130_fd_sc_hd__o22a_1
X_07144_ _07144_/A _07223_/B vssd1 vssd1 vccd1 vccd1 _07144_/X sky130_fd_sc_hd__or2_1
XFILLER_0_15_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07787__A1 _08732_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07075_ _08391_/B _08391_/C vssd1 vssd1 vccd1 vccd1 _07075_/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07787__B2 _10927_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07977_ _07975_/A _07975_/B _07976_/Y vssd1 vssd1 vccd1 vccd1 _08024_/A sky130_fd_sc_hd__o21ai_2
X_06928_ _09157_/B _09170_/B vssd1 vssd1 vccd1 vccd1 _09152_/B sky130_fd_sc_hd__or2_2
XANTENNA__12296__B1 _09163_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09716_ _09716_/A _09716_/B vssd1 vssd1 vccd1 vccd1 _09718_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_96_103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06859_ _06621_/Y _12342_/B _06838_/Y vssd1 vssd1 vccd1 vccd1 _06859_/Y sky130_fd_sc_hd__a21oi_1
X_09647_ _09647_/A _09647_/B vssd1 vssd1 vccd1 vccd1 _10232_/A sky130_fd_sc_hd__xnor2_4
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09578_ _09578_/A _09578_/B vssd1 vssd1 vccd1 vccd1 _09597_/A sky130_fd_sc_hd__xnor2_2
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08529_ _08530_/A _08530_/B vssd1 vssd1 vccd1 vccd1 _08529_/Y sky130_fd_sc_hd__nand2_1
XANTENNA_fanout39_A _12836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08267__A2 _08727_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11540_ _11540_/A _11973_/B vssd1 vssd1 vccd1 vccd1 _11540_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__06726__B _06799_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11471_ _07099_/A fanout6/X _11470_/X _11269_/A vssd1 vssd1 vccd1 vccd1 _11557_/A
+ sky130_fd_sc_hd__a2bb2o_4
X_13210_ _13210_/A hold262/X vssd1 vssd1 vccd1 vccd1 _13372_/D sky130_fd_sc_hd__and2_1
XANTENNA__07227__B1 _10022_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10422_ _10422_/A _10422_/B vssd1 vssd1 vccd1 vccd1 _10424_/C sky130_fd_sc_hd__xor2_1
X_13141_ hold269/X _13140_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13141_/X sky130_fd_sc_hd__mux2_1
X_10353_ _10353_/A _10353_/B vssd1 vssd1 vccd1 vccd1 _10356_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_0_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13072_ hold107/X _12791_/A _13080_/B1 hold97/X _13113_/A vssd1 vssd1 vccd1 vccd1
+ hold108/A sky130_fd_sc_hd__o221a_1
X_12023_ _11865_/Y _12380_/A _12021_/A vssd1 vssd1 vccd1 vccd1 _12023_/X sky130_fd_sc_hd__a21o_1
X_10284_ _10284_/A _10284_/B vssd1 vssd1 vccd1 vccd1 _10285_/B sky130_fd_sc_hd__nor2_1
XANTENNA__08727__B1 _08727_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13079__A2 _13087_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07950__A1 fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07950__B2 _08304_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12925_ _13124_/B _13125_/A _12899_/X vssd1 vssd1 vccd1 vccd1 _13130_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_87_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12856_ hold86/X _12856_/B vssd1 vssd1 vccd1 vccd1 hold87/A sky130_fd_sc_hd__or2_1
XFILLER_0_87_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11807_ hold236/A _11450_/B _11891_/B _11968_/B1 vssd1 vssd1 vccd1 vccd1 _11807_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08258__A2 fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12638__B _12639_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12787_ hold53/X hold167/X vssd1 vssd1 vccd1 vccd1 hold168/A sky130_fd_sc_hd__nand2_1
XFILLER_0_113_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11738_ _12169_/A _11822_/A _11874_/A vssd1 vssd1 vccd1 vccd1 _11790_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_22_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09947__B _09949_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11669_ _11670_/A _11670_/B vssd1 vssd1 vccd1 vccd1 _11768_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_114_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07748__A _08731_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13339_ _13340_/CLK _13339_/D vssd1 vssd1 vccd1 vccd1 hold97/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11565__A2 fanout12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08430__A2 fanout87/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10525__B1 _11973_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08880_ _08880_/A _08880_/B vssd1 vssd1 vccd1 vccd1 _08882_/B sky130_fd_sc_hd__xor2_2
X_07900_ _11758_/A _07900_/B vssd1 vssd1 vccd1 vccd1 _07911_/C sky130_fd_sc_hd__xor2_1
XFILLER_0_20_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07483__A _10707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07831_ _07831_/A _07831_/B vssd1 vssd1 vccd1 vccd1 _07853_/A sky130_fd_sc_hd__xor2_1
XANTENNA__12817__A2 _12818_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09501_ _09102_/X _09128_/X _09666_/S vssd1 vssd1 vccd1 vccd1 _09501_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_79_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07762_ _08722_/A _07762_/B vssd1 vssd1 vccd1 vccd1 _07770_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__09694__A1 _11118_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06713_ _11244_/S _06713_/B vssd1 vssd1 vccd1 vccd1 _11224_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_79_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07693_ _09716_/A _07693_/B vssd1 vssd1 vccd1 vccd1 _07694_/B sky130_fd_sc_hd__xnor2_1
X_06644_ reg1_val[24] _07166_/A vssd1 vssd1 vccd1 vccd1 _12049_/S sky130_fd_sc_hd__nand2_1
XFILLER_0_78_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09432_ _12848_/A _09567_/B _09568_/B _10941_/B vssd1 vssd1 vccd1 vccd1 _09433_/B
+ sky130_fd_sc_hd__o22a_1
X_06575_ instruction[41] vssd1 vssd1 vccd1 vccd1 _06575_/Y sky130_fd_sc_hd__inv_2
X_09363_ _09442_/A _12426_/A _09362_/Y vssd1 vssd1 vccd1 vccd1 _09364_/B sky130_fd_sc_hd__a21oi_1
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout243_A _12394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08314_ _08371_/A vssd1 vssd1 vccd1 vccd1 _08314_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_32 reg2_val[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_10 reg1_val[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_21 reg2_val[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09294_ _09294_/A _09294_/B vssd1 vssd1 vccd1 vccd1 _09296_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_117_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_43 reg1_val[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_65 reg1_val[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11879__S _12341_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_54 reg1_val[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08245_ _08245_/A _08245_/B vssd1 vssd1 vccd1 vccd1 _08246_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_43_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08176_ _08731_/A _08176_/B vssd1 vssd1 vccd1 vccd1 _08215_/B sky130_fd_sc_hd__xnor2_1
X_07127_ _09442_/A _07127_/B vssd1 vssd1 vccd1 vccd1 _07139_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_42_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07058_ reg1_val[13] reg1_val[14] reg1_val[15] _06994_/D _07200_/A vssd1 vssd1 vccd1
+ vccd1 _07069_/B sky130_fd_sc_hd__o41a_4
XFILLER_0_100_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10812__A _11172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11908__A _11908_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09382__B1 _12814_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08185__B2 fanout99/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08185__A1 _08436_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09685__A1 _12388_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10971_ _10971_/A _10971_/B vssd1 vssd1 vccd1 vccd1 _10974_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_97_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12710_ reg1_val[15] _12703_/B _12706_/A vssd1 vssd1 vccd1 vccd1 _12712_/B sky130_fd_sc_hd__a21oi_4
XANTENNA__10295__A2 fanout59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12641_ _12641_/A _12641_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[3] sky130_fd_sc_hd__xnor2_4
XANTENNA__11244__A1 _09354_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12572_ _12623_/A _12573_/B vssd1 vssd1 vccd1 vccd1 _12582_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_93_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11523_ _11523_/A _11523_/B vssd1 vssd1 vccd1 vccd1 _11523_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_18_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11454_ hold277/A _11452_/X _11453_/Y vssd1 vssd1 vccd1 vccd1 _11454_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_80_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10405_ _10780_/A _10779_/D _10405_/C vssd1 vssd1 vccd1 vccd1 _10405_/X sky130_fd_sc_hd__or3_1
XFILLER_0_33_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11385_ _11385_/A _11385_/B vssd1 vssd1 vccd1 vccd1 _11389_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13124_ _12899_/X _13124_/B vssd1 vssd1 vccd1 vccd1 _13125_/B sky130_fd_sc_hd__nand2b_1
X_10336_ _11172_/A _10336_/B vssd1 vssd1 vccd1 vccd1 _10338_/B sky130_fd_sc_hd__xnor2_1
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13055_ _11164_/A _13087_/B2 hold122/X vssd1 vssd1 vccd1 vccd1 _13330_/D sky130_fd_sc_hd__o21a_1
X_10267_ _10267_/A _10267_/B vssd1 vssd1 vccd1 vccd1 _10267_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__06974__A2 _12826_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12006_ _12081_/B _12006_/B vssd1 vssd1 vccd1 vccd1 _12009_/B sky130_fd_sc_hd__nor2_1
X_10198_ _10017_/X _10018_/Y _10021_/B _10029_/A _10029_/B vssd1 vssd1 vccd1 vccd1
+ _10213_/A sky130_fd_sc_hd__a32o_2
XANTENNA__11256__C _11650_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12908_ hold49/X hold284/X vssd1 vssd1 vccd1 vccd1 _12908_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_88_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10286__A2 fanout48/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12839_ hold3/X _12848_/B _12838_/Y _13214_/A vssd1 vssd1 vccd1 vccd1 hold4/A sky130_fd_sc_hd__o211a_1
XFILLER_0_84_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12432__B1 _09167_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11235__A1 _11886_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08030_ _08030_/A _08030_/B _08030_/C vssd1 vssd1 vccd1 vccd1 _08031_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_114_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_5_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13307_/CLK sky130_fd_sc_hd__clkbuf_8
XANTENNA__10108__S _12388_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09600__B2 _12802_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09600__A1 _07026_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10746__B1 _12290_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08403__A2 _10537_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09981_ hold291/A _10124_/C _09835_/B vssd1 vssd1 vccd1 vccd1 _09983_/B sky130_fd_sc_hd__o21a_1
XANTENNA__07611__B1 _10571_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08932_ _08932_/A _08932_/B vssd1 vssd1 vccd1 vccd1 _08934_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__09903__A2 _10589_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout193_A _09433_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08863_ _08863_/A _08863_/B vssd1 vssd1 vccd1 vccd1 _08865_/A sky130_fd_sc_hd__xor2_4
XANTENNA__08102__A _08733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07814_ _07814_/A _07814_/B _07813_/X vssd1 vssd1 vccd1 vccd1 _07816_/B sky130_fd_sc_hd__or3b_1
X_08794_ _08795_/A _08795_/B vssd1 vssd1 vccd1 vccd1 _08794_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_74_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07745_ _07746_/A _07746_/B vssd1 vssd1 vccd1 vccd1 _07745_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__11463__A _11758_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09415_ _09415_/A _09415_/B vssd1 vssd1 vccd1 vccd1 _09418_/A sky130_fd_sc_hd__or2_1
XFILLER_0_67_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07676_ _07676_/A _07676_/B vssd1 vssd1 vccd1 vccd1 _08942_/B sky130_fd_sc_hd__nor2_2
X_06627_ _06625_/X _06627_/B vssd1 vssd1 vccd1 vccd1 _12293_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_66_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09346_ _12244_/S _09345_/Y _06924_/X vssd1 vssd1 vccd1 vccd1 _09346_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_81_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09277_ _09277_/A _09277_/B vssd1 vssd1 vccd1 vccd1 _09280_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_62_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08228_ _07896_/A fanout87/X fanout82/X _08723_/B1 vssd1 vssd1 vccd1 vccd1 _08229_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_90_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08159_ _08159_/A _08159_/B vssd1 vssd1 vccd1 vccd1 _08161_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_15_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10201__A2 _10575_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11170_ _07048_/A _07048_/B fanout48/X vssd1 vssd1 vccd1 vccd1 _11172_/B sky130_fd_sc_hd__a21o_1
X_10121_ _10391_/A2 _10253_/B hold157/A vssd1 vssd1 vccd1 vccd1 _10123_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_100_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10052_ _11564_/A _10052_/B vssd1 vssd1 vccd1 vccd1 _10054_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_97_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10268__A2 _09172_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12111__C1 _11624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11373__A _12210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10954_ _10954_/A _10954_/B vssd1 vssd1 vccd1 vccd1 _10956_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_128_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10885_ reg1_val[12] curr_PC[12] vssd1 vssd1 vccd1 vccd1 _10885_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_97_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12624_ _12624_/A _12624_/B vssd1 vssd1 vccd1 vccd1 new_PC[27] sky130_fd_sc_hd__xnor2_4
XFILLER_0_65_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09778__A _11180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12555_ _12556_/A _12556_/B _12556_/C vssd1 vssd1 vccd1 vccd1 _12566_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_93_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07298__A _10449_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11506_ _11506_/A _11506_/B vssd1 vssd1 vccd1 vccd1 _11508_/C sky130_fd_sc_hd__xor2_1
X_12486_ _12495_/A _12486_/B vssd1 vssd1 vccd1 vccd1 _12488_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_81_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11437_ _11437_/A _11437_/B vssd1 vssd1 vccd1 vccd1 _11437_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_21_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11368_ _11369_/A _11369_/B vssd1 vssd1 vccd1 vccd1 _11370_/A sky130_fd_sc_hd__nor2_1
X_13107_ hold284/X _13106_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13107_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_95_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10319_ _10444_/A _10319_/B vssd1 vssd1 vccd1 vccd1 _10324_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__13142__B2 _12790_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09346__B1 _06924_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11299_ _11158_/A _11158_/B _11159_/X vssd1 vssd1 vccd1 vccd1 _11301_/A sky130_fd_sc_hd__a21o_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13038_ hold148/X _12788_/A _13236_/B hold155/X _13109_/A vssd1 vssd1 vccd1 vccd1
+ hold156/A sky130_fd_sc_hd__o221a_1
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07530_ _07527_/B _07577_/B _07527_/A vssd1 vssd1 vccd1 vccd1 _07556_/A sky130_fd_sc_hd__o21bai_2
XANTENNA__07124__A2 _09343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07461_ _10818_/A _10570_/A _10571_/A _10963_/A vssd1 vssd1 vccd1 vccd1 _07462_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_9_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09200_ _09200_/A _09200_/B vssd1 vssd1 vccd1 vccd1 _09203_/A sky130_fd_sc_hd__nand2_1
X_07392_ _07393_/A _07393_/B vssd1 vssd1 vccd1 vccd1 _07392_/X sky130_fd_sc_hd__or2_1
XFILLER_0_57_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12826__B _12830_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09131_ reg1_val[0] reg1_val[31] _09142_/S vssd1 vssd1 vccd1 vccd1 _09131_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_60_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11759__A2 fanout12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09062_ _08912_/A _08912_/B _08939_/A _08939_/B vssd1 vssd1 vccd1 vccd1 _09073_/C
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_60_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07832__B1 _09396_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10431__A2 fanout16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12842__A _12842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08013_ _08013_/A _08013_/B vssd1 vssd1 vccd1 vccd1 _08015_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_4_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08388__A1 _07885_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08388__B2 _08721_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_83 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09585__B1 _11766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09964_ _09964_/A _09964_/B vssd1 vssd1 vccd1 vccd1 _09964_/X sky130_fd_sc_hd__xor2_1
XANTENNA__10362__A _10364_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08915_ _08017_/A _08017_/B _08018_/Y vssd1 vssd1 vccd1 vccd1 _08937_/A sky130_fd_sc_hd__a21bo_2
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09895_ _10941_/B _10167_/A1 _10022_/B1 _09568_/A vssd1 vssd1 vccd1 vccd1 _09896_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07899__B1 _08752_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08846_ _08845_/A _08845_/B _08845_/C vssd1 vssd1 vccd1 vccd1 _08847_/B sky130_fd_sc_hd__a21oi_1
X_08777_ _08778_/B _08778_/A vssd1 vssd1 vccd1 vccd1 _08777_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_94_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07728_ _07835_/A _07835_/B _07724_/X vssd1 vssd1 vccd1 vccd1 _07744_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__08312__A1 fanout99/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07659_ _09567_/B _10574_/B _11751_/A _09568_/B vssd1 vssd1 vccd1 vccd1 _07660_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08312__B2 _12818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09598__A _09598_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10670_ _10669_/B _10669_/C _10669_/A vssd1 vssd1 vccd1 vccd1 _10681_/B sky130_fd_sc_hd__a21oi_1
X_09329_ _09120_/X _09123_/X _09330_/S vssd1 vssd1 vccd1 vccd1 _09329_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_75_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10958__B1 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12340_ _06627_/B _12291_/X _06625_/X vssd1 vssd1 vccd1 vccd1 _12341_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_62_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07823__B1 _11908_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12271_ _12271_/A _12321_/B vssd1 vssd1 vccd1 vccd1 _12272_/B sky130_fd_sc_hd__nand2_1
X_11222_ _11111_/A _11109_/X _11130_/S vssd1 vssd1 vccd1 vccd1 _11222_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_105_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09576__B1 _10022_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06929__A2 _06924_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11153_ _12317_/A _11153_/B vssd1 vssd1 vccd1 vccd1 _11160_/A sky130_fd_sc_hd__xnor2_1
X_10104_ _10000_/X _10275_/B _10103_/Y vssd1 vssd1 vccd1 vccd1 _10104_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__09879__A1 _09609_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11084_ _10953_/Y _10957_/A _11085_/B vssd1 vssd1 vccd1 vccd1 _11084_/X sky130_fd_sc_hd__a21o_1
XANTENNA__09879__B2 _09396_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10035_ _10036_/B _10036_/C _10959_/A vssd1 vssd1 vccd1 vccd1 _10040_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__06909__B _06921_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11986_ _12169_/A _12169_/B _12169_/C vssd1 vssd1 vccd1 vccd1 _12030_/B sky130_fd_sc_hd__or3_1
XFILLER_0_98_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10937_ _12076_/A _10937_/B vssd1 vssd1 vccd1 vccd1 _10938_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_14_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12607_ _12607_/A _12607_/B _12607_/C _12607_/D vssd1 vssd1 vccd1 vccd1 _12608_/B
+ sky130_fd_sc_hd__and4_2
XANTENNA__06665__A2_N _06771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10868_ _10868_/A vssd1 vssd1 vccd1 vccd1 _10870_/D sky130_fd_sc_hd__inv_2
XFILLER_0_6_718 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06644__B _07166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10799_ _10959_/A _10799_/B _10799_/C vssd1 vssd1 vccd1 vccd1 _10800_/C sky130_fd_sc_hd__nor3_1
XFILLER_0_121_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12538_ _12544_/B _12538_/B vssd1 vssd1 vccd1 vccd1 new_PC[13] sky130_fd_sc_hd__and2_4
XFILLER_0_54_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12469_ reg1_val[4] curr_PC[4] _12622_/S vssd1 vssd1 vccd1 vccd1 _12471_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11374__B1 _12213_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10182__A _10448_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06961_ _06964_/A _06964_/B vssd1 vssd1 vccd1 vccd1 _06961_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__07066__C_N _06963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_86 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09680_ _10250_/S _09137_/X _09176_/B vssd1 vssd1 vccd1 vccd1 _09680_/X sky130_fd_sc_hd__o21a_1
X_08700_ _08571_/A _08571_/B _08571_/C vssd1 vssd1 vccd1 vccd1 _08703_/B sky130_fd_sc_hd__o21a_1
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06892_ hold160/A _06892_/B vssd1 vssd1 vccd1 vccd1 busy sky130_fd_sc_hd__nor2_8
X_08631_ _09445_/A _08631_/B vssd1 vssd1 vccd1 vccd1 _08636_/A sky130_fd_sc_hd__xnor2_1
X_08562_ _08798_/B2 _09567_/B _09568_/B _08646_/B2 vssd1 vssd1 vccd1 vccd1 _08563_/B
+ sky130_fd_sc_hd__o22a_1
X_07513_ _07514_/A _07514_/B vssd1 vssd1 vccd1 vccd1 _07513_/X sky130_fd_sc_hd__and2b_1
X_08493_ _08493_/A _08493_/B vssd1 vssd1 vccd1 vccd1 _08494_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_49_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07444_ _07445_/A _07445_/B vssd1 vssd1 vccd1 vccd1 _07446_/A sky130_fd_sc_hd__or2_1
Xfanout38 _12836_/A vssd1 vssd1 vccd1 vccd1 _11766_/A sky130_fd_sc_hd__buf_6
Xfanout16 _07262_/X vssd1 vssd1 vccd1 vccd1 fanout16/X sky130_fd_sc_hd__buf_8
Xfanout27 _07688_/B vssd1 vssd1 vccd1 vccd1 fanout27/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__11741__A _12261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout49 _07191_/Y vssd1 vssd1 vccd1 vccd1 _12838_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_9_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07375_ _07376_/A _07376_/B _07376_/C vssd1 vssd1 vccd1 vccd1 _07579_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_45_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09114_ _09106_/X _09113_/X _09974_/A vssd1 vssd1 vccd1 vccd1 _09114_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_45_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09045_ _09049_/A _09045_/B vssd1 vssd1 vccd1 vccd1 _11953_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11365__B1 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08230__B1 _07821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09947_ _09949_/A _09949_/B vssd1 vssd1 vccd1 vccd1 _09947_/X sky130_fd_sc_hd__or2_1
XANTENNA__09092__S _09108_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08497__A _09441_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08533__A1 _08646_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08533__B2 _09423_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09878_ _09878_/A _09878_/B vssd1 vssd1 vccd1 vccd1 _09881_/A sky130_fd_sc_hd__xor2_4
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06729__B _07074_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08829_ _08829_/A _08829_/B vssd1 vssd1 vccd1 vccd1 _08831_/B sky130_fd_sc_hd__xnor2_2
XTAP_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11840_ _11840_/A _11840_/B vssd1 vssd1 vccd1 vccd1 _11856_/A sky130_fd_sc_hd__xor2_1
XTAP_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11771_ _11772_/A _11772_/B _11772_/C vssd1 vssd1 vccd1 vccd1 _11824_/A sky130_fd_sc_hd__o21ai_1
XTAP_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10722_ _10722_/A _10722_/B vssd1 vssd1 vccd1 vccd1 _10724_/B sky130_fd_sc_hd__nor2_1
XTAP_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10653_ _09152_/Y _10638_/X _10640_/X _10652_/Y _10630_/X vssd1 vssd1 vccd1 vccd1
+ _10653_/X sky130_fd_sc_hd__a2111o_1
XFILLER_0_35_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_391 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13372_ _13378_/CLK _13372_/D vssd1 vssd1 vccd1 vccd1 hold261/A sky130_fd_sc_hd__dfxtp_1
X_10584_ _10585_/A _10585_/B vssd1 vssd1 vccd1 vccd1 _10584_/Y sky130_fd_sc_hd__nand2_1
X_12323_ _12373_/A _12323_/B vssd1 vssd1 vccd1 vccd1 _12325_/C sky130_fd_sc_hd__or2_1
XFILLER_0_106_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09549__B1 _10567_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12254_ _12254_/A1 _09821_/X _09828_/Y _10113_/A _12253_/Y vssd1 vssd1 vccd1 vccd1
+ _12254_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_50_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12185_ _12185_/A _12185_/B vssd1 vssd1 vccd1 vccd1 _12185_/Y sky130_fd_sc_hd__xnor2_1
X_11205_ _11205_/A _11205_/B vssd1 vssd1 vccd1 vccd1 _11207_/B sky130_fd_sc_hd__xnor2_1
X_11136_ _12254_/A1 _11121_/B _11135_/Y _10113_/A _11133_/X vssd1 vssd1 vccd1 vccd1
+ _11136_/X sky130_fd_sc_hd__o221a_1
XANTENNA__11659__A1 _11847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08524__B2 _08721_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08524__A1 _08730_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11067_ _12138_/A _11067_/B vssd1 vssd1 vccd1 vccd1 _11069_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__11659__B2 _11766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10018_ _10019_/A _10019_/B vssd1 vssd1 vccd1 vccd1 _10018_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__10331__B2 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10331__A1 _11065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11969_ _11969_/A _11969_/B vssd1 vssd1 vccd1 vccd1 _11969_/X sky130_fd_sc_hd__or2_1
XFILLER_0_86_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07160_ _07200_/A _07160_/B vssd1 vssd1 vccd1 vccd1 _07161_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_27_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07091_ _12808_/A _11653_/A _12810_/A _08752_/B vssd1 vssd1 vccd1 vccd1 _07092_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_14_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08460__B1 _08656_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10624__B _10624_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07015__A1 _09666_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout217 _06891_/Y vssd1 vssd1 vccd1 vccd1 _13080_/B1 sky130_fd_sc_hd__buf_4
Xfanout228 _12794_/A vssd1 vssd1 vccd1 vccd1 _09336_/S sky130_fd_sc_hd__buf_4
Xfanout206 _09165_/X vssd1 vssd1 vccd1 vccd1 _09354_/B sky130_fd_sc_hd__buf_4
X_09801_ _09802_/B _09802_/A vssd1 vssd1 vccd1 vccd1 _09801_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_5_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout239 _07050_/A vssd1 vssd1 vccd1 vccd1 _11233_/S sky130_fd_sc_hd__buf_4
X_09732_ _09732_/A _09732_/B _09732_/C vssd1 vssd1 vccd1 vccd1 _09733_/B sky130_fd_sc_hd__nor3_1
X_07993_ _07993_/A _07993_/B vssd1 vssd1 vccd1 vccd1 _07994_/A sky130_fd_sc_hd__and2_1
X_06944_ reg1_val[10] reg1_val[11] reg1_val[12] _07200_/B vssd1 vssd1 vccd1 vccd1
+ _06994_/D sky130_fd_sc_hd__or4_4
X_09663_ _09319_/X _09321_/X _09663_/S vssd1 vssd1 vccd1 vccd1 _09663_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout273_A _12788_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06875_ _06874_/X _08980_/B instruction[6] vssd1 vssd1 vccd1 vccd1 _06875_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_96_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09594_ _09594_/A _09594_/B vssd1 vssd1 vccd1 vccd1 _09596_/B sky130_fd_sc_hd__xnor2_2
X_08614_ _08606_/A _08605_/C _08605_/B vssd1 vssd1 vccd1 vccd1 _08615_/C sky130_fd_sc_hd__a21o_1
XANTENNA__10873__A2 _10871_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08545_ _08574_/A _08545_/B vssd1 vssd1 vccd1 vccd1 _08549_/A sky130_fd_sc_hd__xnor2_1
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12075__A1 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12075__B2 fanout27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08476_ _08681_/A _08476_/B vssd1 vssd1 vccd1 vccd1 _08508_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_65_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07427_ _07427_/A _07427_/B vssd1 vssd1 vccd1 vccd1 _07438_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_64_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07358_ _12826_/A _10948_/B2 _12824_/A fanout74/X vssd1 vssd1 vccd1 vccd1 _07359_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09876__A _11261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09779__B1 _08752_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07289_ _09445_/A _07289_/B vssd1 vssd1 vccd1 vccd1 _07647_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__11050__A2 _12213_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09028_ _09028_/A _09028_/B vssd1 vssd1 vccd1 vccd1 _11521_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold271 hold271/A vssd1 vssd1 vccd1 vccd1 hold271/X sky130_fd_sc_hd__buf_1
Xhold260 hold260/A vssd1 vssd1 vccd1 vccd1 hold260/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold293 hold293/A vssd1 vssd1 vccd1 vccd1 hold293/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 hold282/A vssd1 vssd1 vccd1 vccd1 hold282/X sky130_fd_sc_hd__dlygate4sd3_1
X_12941_ _13188_/B _13189_/A _12875_/X vssd1 vssd1 vccd1 vccd1 _13193_/A sky130_fd_sc_hd__a21o_1
XANTENNA__06780__A3 _12649_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12872_ hold1/X hold246/X vssd1 vssd1 vccd1 vccd1 _12872_/X sky130_fd_sc_hd__and2b_1
X_11823_ _12169_/A _12169_/B vssd1 vssd1 vccd1 vccd1 _11872_/B sky130_fd_sc_hd__or2_1
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12477__A _12649_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11813__A1 _07135_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11754_ _11754_/A _11754_/B vssd1 vssd1 vccd1 vccd1 _11755_/B sky130_fd_sc_hd__and2_1
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07493__B2 _09236_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07493__A1 _09444_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08393__C _08393_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11685_ _11685_/A _11685_/B vssd1 vssd1 vccd1 vccd1 _11687_/C sky130_fd_sc_hd__xnor2_1
X_10705_ _10566_/A _10566_/B _10568_/X vssd1 vssd1 vccd1 vccd1 _10716_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_125_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10636_ _10636_/A _10636_/B _10636_/C vssd1 vssd1 vccd1 vccd1 _10636_/X sky130_fd_sc_hd__and3_1
XFILLER_0_70_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12369__A2 _12316_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13355_ _13355_/CLK _13355_/D vssd1 vssd1 vccd1 vccd1 hold273/A sky130_fd_sc_hd__dfxtp_1
X_10567_ _10567_/A _12316_/B vssd1 vssd1 vccd1 vccd1 _10569_/B sky130_fd_sc_hd__or2_1
XANTENNA__11041__A2 _12316_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12306_ hold169/A _12434_/B1 _12355_/B _12401_/B1 vssd1 vssd1 vccd1 vccd1 _12306_/X
+ sky130_fd_sc_hd__a31o_1
X_13286_ _13311_/CLK hold199/X vssd1 vssd1 vccd1 vccd1 hold234/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10498_ _09307_/A _09307_/B _09953_/X _10496_/X vssd1 vssd1 vccd1 vccd1 _10499_/C
+ sky130_fd_sc_hd__a211o_1
XANTENNA__07796__A2 fanout87/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12237_ _09059_/A _09059_/B _12170_/A vssd1 vssd1 vccd1 vccd1 _12238_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_121_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12168_ _12030_/C _12168_/B vssd1 vssd1 vccd1 vccd1 _12169_/D sky130_fd_sc_hd__nand2b_1
XANTENNA__10552__A1 _10963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10552__B2 _11065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11556__A _11557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11119_ _11010_/S _10115_/X _11118_/X _11233_/S vssd1 vssd1 vccd1 vccd1 _11119_/X
+ sky130_fd_sc_hd__o211a_1
X_12099_ _12099_/A _12099_/B vssd1 vssd1 vccd1 vccd1 _12099_/X sky130_fd_sc_hd__and2_1
X_06660_ reg1_val[22] _07191_/A vssd1 vssd1 vccd1 vccd1 _11894_/A sky130_fd_sc_hd__and2_1
XFILLER_0_78_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07720__A2 _11751_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06591_ instruction[1] instruction[2] instruction[25] pred_val vssd1 vssd1 vccd1
+ vccd1 _06591_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_59_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11804__A1 _11886_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08330_ _08330_/A _08330_/B vssd1 vssd1 vccd1 vccd1 _08331_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_86_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07484__A1 _12824_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07484__B2 _12826_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08261_ _08436_/A _08732_/A2 _08656_/B fanout99/X vssd1 vssd1 vccd1 vccd1 _08262_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_6_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07212_ _10710_/A _07212_/B vssd1 vssd1 vccd1 vccd1 _07214_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08192_ _08740_/A _08192_/B vssd1 vssd1 vccd1 vccd1 _08197_/A sky130_fd_sc_hd__xnor2_2
X_07143_ _07144_/A _07142_/B _07142_/C _07142_/D _07223_/B vssd1 vssd1 vccd1 vccd1
+ _07151_/B sky130_fd_sc_hd__a41o_2
XFILLER_0_42_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07074_ _07074_/A _07074_/B _07074_/C vssd1 vssd1 vccd1 vccd1 _08391_/C sky130_fd_sc_hd__nand3_2
XANTENNA__10240__B1 _09163_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout119_A _11367_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07787__A2 _08744_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11740__B1 fanout4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07976_ _08027_/B _08027_/A vssd1 vssd1 vccd1 vccd1 _07976_/Y sky130_fd_sc_hd__nand2b_1
X_06927_ _09157_/B _09170_/B vssd1 vssd1 vccd1 vccd1 _09153_/B sky130_fd_sc_hd__nor2_1
X_09715_ fanout23/X _10664_/A _10818_/A _07819_/B vssd1 vssd1 vccd1 vccd1 _09716_/B
+ sky130_fd_sc_hd__o22a_1
X_09646_ _09647_/A _09647_/B vssd1 vssd1 vccd1 vccd1 _09646_/X sky130_fd_sc_hd__and2_1
XFILLER_0_96_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06858_ _12293_/A _06857_/Y _06839_/Y vssd1 vssd1 vccd1 vccd1 _12342_/B sky130_fd_sc_hd__o21ai_1
X_06789_ reg1_val[3] _11010_/S vssd1 vssd1 vccd1 vccd1 _06789_/Y sky130_fd_sc_hd__nor2_1
X_09577_ _10449_/A _09577_/B vssd1 vssd1 vccd1 vccd1 _09578_/B sky130_fd_sc_hd__xnor2_2
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08528_ _08598_/A _08528_/B vssd1 vssd1 vccd1 vccd1 _08560_/A sky130_fd_sc_hd__xnor2_1
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08459_ _08459_/A _08459_/B vssd1 vssd1 vccd1 vccd1 _08514_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_38_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11470_ _11470_/A _11470_/B fanout6/X vssd1 vssd1 vccd1 vccd1 _11470_/X sky130_fd_sc_hd__or3_1
XANTENNA__06742__B _07100_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07227__A1 _10167_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07227__B2 _12836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10421_ _07087_/A _07087_/B _10575_/B _10930_/B fanout66/X vssd1 vssd1 vccd1 vccd1
+ _10422_/B sky130_fd_sc_hd__o32a_1
XANTENNA__10545__A _11163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13140_ _13140_/A _13140_/B vssd1 vssd1 vccd1 vccd1 _13140_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_61_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10352_ _10352_/A _10352_/B vssd1 vssd1 vccd1 vccd1 _10353_/B sky130_fd_sc_hd__xor2_2
XANTENNA__06771__C_N _12654_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13071_ _11987_/A _13077_/A2 hold117/X vssd1 vssd1 vccd1 vccd1 _13338_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_20_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12022_ _12165_/A _12165_/B vssd1 vssd1 vccd1 vccd1 _12380_/A sky130_fd_sc_hd__nor2_1
X_10283_ _10284_/A _10284_/B vssd1 vssd1 vccd1 vccd1 _10285_/A sky130_fd_sc_hd__and2_1
XANTENNA__08727__A1 _11367_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08727__B2 _11472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10280__A _11470_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07950__A2 _07885_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12924_ _13119_/B _13120_/A _12901_/X vssd1 vssd1 vccd1 vccd1 _13125_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_88_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12855_ hold11/X _12856_/B _12854_/Y _13235_/A vssd1 vssd1 vccd1 vccd1 hold12/A sky130_fd_sc_hd__o211a_1
XANTENNA__06917__B _06921_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11806_ _11450_/B _11891_/B hold236/A vssd1 vssd1 vccd1 vccd1 _11806_/Y sky130_fd_sc_hd__a21oi_1
X_12786_ hold167/A vssd1 vssd1 vccd1 vccd1 _12786_/Y sky130_fd_sc_hd__inv_2
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12000__A _12210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11737_ _11142_/S _11733_/X _11736_/X vssd1 vssd1 vccd1 vccd1 dest_val[20] sky130_fd_sc_hd__o21ai_4
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08663__B1 _08436_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06933__A _12455_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12654__B _12654_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11668_ _12073_/A _11668_/B vssd1 vssd1 vccd1 vccd1 _11670_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10619_ _10861_/C _10491_/Y _10492_/X vssd1 vssd1 vccd1 vccd1 _10619_/Y sky130_fd_sc_hd__a21oi_1
X_11599_ _11599_/A _11599_/B vssd1 vssd1 vccd1 vccd1 _11601_/B sky130_fd_sc_hd__nor2_1
X_13338_ _13340_/CLK _13338_/D vssd1 vssd1 vccd1 vccd1 hold107/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_605 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13269_ _13365_/CLK hold48/X vssd1 vssd1 vccd1 vccd1 hold47/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10525__A1 _07095_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07764__A _08740_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07830_ _07831_/A _07831_/B vssd1 vssd1 vccd1 vccd1 _07830_/X sky130_fd_sc_hd__and2_1
X_07761_ _08432_/B _08741_/B2 _12820_/A _10537_/A1 vssd1 vssd1 vccd1 vccd1 _07762_/B
+ sky130_fd_sc_hd__o22a_1
X_06712_ reg1_val[15] _06988_/A vssd1 vssd1 vccd1 vccd1 _06713_/B sky130_fd_sc_hd__nor2_1
X_09500_ _09498_/X _09499_/X _10250_/S vssd1 vssd1 vccd1 vccd1 _09500_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09679__C1 _09172_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09694__A2 _06939_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07692_ _08671_/B2 fanout24/X _07819_/B _07821_/A vssd1 vssd1 vccd1 vccd1 _07693_/B
+ sky130_fd_sc_hd__o22a_1
X_06643_ _06641_/Y _06703_/B1 _06720_/B reg2_val[24] vssd1 vssd1 vccd1 vccd1 _07166_/A
+ sky130_fd_sc_hd__a2bb2o_2
X_09431_ _09431_/A _09431_/B vssd1 vssd1 vccd1 vccd1 _09435_/A sky130_fd_sc_hd__xnor2_1
X_09362_ _09442_/A _12426_/A _08680_/A vssd1 vssd1 vccd1 vccd1 _09362_/Y sky130_fd_sc_hd__o21ai_1
X_06574_ _12626_/A vssd1 vssd1 vccd1 vccd1 _06574_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_47_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07004__A _12341_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08313_ _08728_/A _08313_/B vssd1 vssd1 vccd1 vccd1 _08371_/A sky130_fd_sc_hd__xnor2_2
XANTENNA_11 reg1_val[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_22 reg2_val[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09293_ _07590_/A _07590_/B _07588_/Y vssd1 vssd1 vccd1 vccd1 _09294_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_19_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_44 reg1_val[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_33 reg2_val[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_66 _12804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_55 reg1_val[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10461__B1 fanout59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08244_ _08244_/A _08244_/B vssd1 vssd1 vccd1 vccd1 _08296_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__07209__A1 _07131_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08175_ _08730_/A1 _10927_/A1 _08732_/A1 _08038_/A vssd1 vssd1 vccd1 vccd1 _08176_/B
+ sky130_fd_sc_hd__o22a_1
X_07126_ _09442_/A _07127_/B vssd1 vssd1 vccd1 vccd1 _07139_/A sky130_fd_sc_hd__or2_1
XFILLER_0_43_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09365__S _09666_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07057_ _07057_/A _07057_/B vssd1 vssd1 vccd1 vccd1 _07671_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__09382__B2 _07819_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09382__A1 fanout23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08185__A2 _08741_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12269__A1 _12210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07959_ _11758_/A _07959_/B vssd1 vssd1 vccd1 vccd1 _08030_/C sky130_fd_sc_hd__xor2_1
XANTENNA_fanout51_A _12844_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10970_ _10825_/B _10839_/B _10823_/A vssd1 vssd1 vccd1 vccd1 _10981_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_97_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09629_ _09629_/A _09629_/B vssd1 vssd1 vccd1 vccd1 _09630_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_38_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12640_ _12638_/Y _12640_/B vssd1 vssd1 vccd1 vccd1 _12641_/B sky130_fd_sc_hd__and2b_2
XFILLER_0_77_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12571_ reg1_val[19] curr_PC[19] _12586_/S vssd1 vssd1 vccd1 vccd1 _12573_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_26_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11522_ _11792_/A _11521_/B _11521_/C vssd1 vssd1 vccd1 vccd1 _11523_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_18_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11453_ hold277/A _11452_/X _09167_/Y vssd1 vssd1 vccd1 vccd1 _11453_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_92_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10404_ curr_PC[7] _10403_/C curr_PC[8] vssd1 vssd1 vccd1 vccd1 _10405_/C sky130_fd_sc_hd__a21oi_1
XFILLER_0_21_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13123_ _13128_/A _13123_/B vssd1 vssd1 vccd1 vccd1 _13354_/D sky130_fd_sc_hd__and2_1
XFILLER_0_61_593 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11384_ _11384_/A _11385_/B vssd1 vssd1 vccd1 vccd1 _11475_/A sky130_fd_sc_hd__and2_1
X_10335_ _11146_/A fanout23/X _11171_/A _11294_/A vssd1 vssd1 vccd1 vccd1 _10336_/B
+ sky130_fd_sc_hd__o22a_1
X_13054_ hold121/X _12791_/A _13080_/B1 hold76/X _13113_/A vssd1 vssd1 vccd1 vccd1
+ hold122/A sky130_fd_sc_hd__o221a_1
X_10266_ _10264_/Y _10266_/B vssd1 vssd1 vccd1 vccd1 _10267_/B sky130_fd_sc_hd__and2b_1
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12005_ _12005_/A _12005_/B vssd1 vssd1 vccd1 vccd1 _12006_/B sky130_fd_sc_hd__and2_1
XFILLER_0_108_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10197_ _10197_/A _10197_/B vssd1 vssd1 vccd1 vccd1 _10214_/A sky130_fd_sc_hd__nor2_2
X_12907_ _12905_/X _12907_/B vssd1 vssd1 vccd1 vccd1 _13110_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_88_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12649__B _12649_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12838_ _12838_/A _12848_/B vssd1 vssd1 vccd1 vccd1 _12838_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_33_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12769_ _12773_/B _12769_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[28] sky130_fd_sc_hd__nor2_8
XFILLER_0_127_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10443__B1 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09600__A2 fanout9/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09980_ hold185/A _09980_/B vssd1 vssd1 vccd1 vccd1 _09980_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__07611__B2 _10413_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07611__A1 _12810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07494__A _09594_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08931_ _08016_/A _08016_/B _08014_/X vssd1 vssd1 vccd1 vccd1 _08932_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08862_ _08863_/A _08863_/B vssd1 vssd1 vccd1 vccd1 _08862_/X sky130_fd_sc_hd__and2_1
X_07813_ _07813_/A _07813_/B vssd1 vssd1 vccd1 vccd1 _07813_/X sky130_fd_sc_hd__xor2_1
XANTENNA_fanout186_A _08740_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08793_ _08793_/A _08793_/B vssd1 vssd1 vccd1 vccd1 _08795_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_74_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07744_ _07744_/A _07744_/B vssd1 vssd1 vccd1 vccd1 _07746_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07675_ _07675_/A _07675_/B vssd1 vssd1 vccd1 vccd1 _07676_/B sky130_fd_sc_hd__and2_1
X_06626_ reg1_val[28] _07343_/B vssd1 vssd1 vccd1 vccd1 _06627_/B sky130_fd_sc_hd__nand2b_1
X_09414_ _09235_/A _09235_/B _09232_/A vssd1 vssd1 vccd1 vccd1 _09420_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_90_50 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09345_ _09345_/A _09345_/B vssd1 vssd1 vccd1 vccd1 _09345_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11631__C1 _09172_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09276_ _10422_/A _09276_/B vssd1 vssd1 vccd1 vccd1 _09277_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_47_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10434__B1 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08227_ _08238_/A _08238_/B vssd1 vssd1 vccd1 vccd1 _08227_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_16_730 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10095__A _10096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08158_ _08158_/A _08158_/B vssd1 vssd1 vccd1 vccd1 _08159_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_113_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07109_ _07522_/A _07109_/B vssd1 vssd1 vccd1 vccd1 _07113_/A sky130_fd_sc_hd__xnor2_1
X_08089_ _08745_/A _08089_/B vssd1 vssd1 vccd1 vccd1 _08146_/B sky130_fd_sc_hd__xnor2_1
X_10120_ hold185/A hold187/A _10120_/C vssd1 vssd1 vccd1 vccd1 _10253_/B sky130_fd_sc_hd__or3_1
XANTENNA__11638__B _11973_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09095__S _09108_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout99_A _12816_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10051_ _10570_/A _10574_/B _11751_/A _10571_/A vssd1 vssd1 vccd1 vccd1 _10052_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_100_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07118__B1 _07200_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11654__A _11758_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10953_ _10954_/A _10954_/B vssd1 vssd1 vccd1 vccd1 _10953_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_58_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10673__B1 _10570_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10884_ reg1_val[12] curr_PC[12] vssd1 vssd1 vccd1 vccd1 _10884_/X sky130_fd_sc_hd__or2_1
XFILLER_0_85_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12623_ _12623_/A _12623_/B vssd1 vssd1 vccd1 vccd1 _12624_/B sky130_fd_sc_hd__xor2_2
XANTENNA__12485__A _12654_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08618__B1 _09440_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12554_ _12623_/A _12554_/B vssd1 vssd1 vccd1 vccd1 _12556_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_66_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11505_ _11506_/A _11506_/B vssd1 vssd1 vccd1 vccd1 _11603_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_124_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12485_ _12654_/B _12485_/B vssd1 vssd1 vccd1 vccd1 _12486_/B sky130_fd_sc_hd__or2_1
XFILLER_0_41_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11436_ _06824_/Y _11435_/Y _12174_/S vssd1 vssd1 vccd1 vccd1 _11437_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_61_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11367_ _11367_/A _12214_/B vssd1 vssd1 vccd1 vccd1 _11369_/B sky130_fd_sc_hd__or2_1
XANTENNA__11829__A _12210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_max_cap151_A _11164_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13106_ _13106_/A _13106_/B vssd1 vssd1 vccd1 vccd1 _13106_/Y sky130_fd_sc_hd__xnor2_1
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10318_ _09568_/A _10589_/A _08507_/B fanout13/X vssd1 vssd1 vccd1 vccd1 _10319_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__13142__A2 _12789_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13037_ _07188_/B _12798_/B hold149/X vssd1 vssd1 vccd1 vccd1 _13321_/D sky130_fd_sc_hd__a21boi_1
XANTENNA__09346__A1 _12244_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11298_ _11191_/A _11190_/B _11188_/X vssd1 vssd1 vccd1 vccd1 _11308_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_119_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10249_ _10247_/X _10248_/X _11231_/S vssd1 vssd1 vccd1 vccd1 _10249_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12350__B1 _12429_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11564__A _11564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11456__A2 _11121_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07460_ _07460_/A _07460_/B vssd1 vssd1 vccd1 vccd1 _07470_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_9_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12405__A1 _09127_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07391_ _07389_/A _07389_/B _07390_/X vssd1 vssd1 vccd1 vccd1 _07393_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_57_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09130_ _09122_/X _09129_/X _09974_/A vssd1 vssd1 vccd1 vccd1 _10385_/B sky130_fd_sc_hd__mux2_1
XANTENNA__07489__A _08724_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09061_ _09061_/A _09061_/B vssd1 vssd1 vccd1 vccd1 _09077_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_60_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08012_ _07697_/Y _07719_/B _07717_/X vssd1 vssd1 vccd1 vccd1 _08015_/A sky130_fd_sc_hd__a21o_2
XANTENNA__07832__A1 _07896_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07832__B2 _08723_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08388__A2 _08732_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09585__A1 fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09585__B2 _08304_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout101_A _07485_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09963_ _06812_/X _09962_/X _12388_/S vssd1 vssd1 vccd1 vccd1 _09964_/B sky130_fd_sc_hd__mux2_1
XANTENNA__06840__B _07144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08914_ _08022_/A _08022_/B _08020_/X vssd1 vssd1 vccd1 vccd1 _08939_/A sky130_fd_sc_hd__a21o_2
XANTENNA__10362__B _10364_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08113__A _08722_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09894_ _10165_/A _09894_/B vssd1 vssd1 vccd1 vccd1 _09900_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_0_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07899__B2 _07752_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07899__A1 _07821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08845_ _08845_/A _08845_/B _08845_/C vssd1 vssd1 vccd1 vccd1 _08847_/A sky130_fd_sc_hd__and3_1
XFILLER_0_109_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08776_ _08208_/A _08206_/Y _08205_/Y vssd1 vssd1 vccd1 vccd1 _08778_/B sky130_fd_sc_hd__o21a_1
X_07727_ _07727_/A _07727_/B vssd1 vssd1 vccd1 vccd1 _07835_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__11447__A2 _11973_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08312__A2 _08727_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07658_ _07664_/B _07664_/A vssd1 vssd1 vccd1 vccd1 _07658_/Y sky130_fd_sc_hd__nand2b_1
X_06609_ _06608_/Y _06703_/B1 _06720_/B reg2_val[30] vssd1 vssd1 vccd1 vccd1 _06612_/B
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_94_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07589_ _07589_/A _07589_/B vssd1 vssd1 vccd1 vccd1 _07590_/B sky130_fd_sc_hd__xor2_4
XANTENNA__09598__B _12264_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09328_ _09326_/X _09327_/X _09669_/S vssd1 vssd1 vccd1 vccd1 _09328_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_75_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10818__A _10818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10958__A1 _11146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10958__B2 _11065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09259_ _09379_/B _09258_/B _09258_/C vssd1 vssd1 vccd1 vccd1 _09260_/C sky130_fd_sc_hd__a21oi_2
XFILLER_0_63_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12270_ _12271_/A _12321_/B vssd1 vssd1 vccd1 vccd1 _12327_/A sky130_fd_sc_hd__or2_1
XANTENNA__12244__S _12244_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09576__B2 _12848_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09576__A1 _12846_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11221_ _11221_/A _11221_/B vssd1 vssd1 vccd1 vccd1 _11221_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__11649__A _11649_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10553__A _10928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11152_ _11472_/A fanout15/X fanout36/X _11558_/A vssd1 vssd1 vccd1 vccd1 _11153_/B
+ sky130_fd_sc_hd__o22a_1
X_10103_ _10000_/X _10275_/B _11707_/A vssd1 vssd1 vccd1 vccd1 _10103_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__07339__B1 _10941_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09879__A2 _09745_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11083_ _10964_/A _10964_/B _10962_/A vssd1 vssd1 vccd1 vccd1 _11085_/B sky130_fd_sc_hd__o21a_1
X_10034_ _12810_/A _10797_/B vssd1 vssd1 vccd1 vccd1 _10036_/C sky130_fd_sc_hd__nor2_1
XANTENNA__11384__A _11384_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11985_ _11985_/A _11985_/B vssd1 vssd1 vccd1 vccd1 _12169_/C sky130_fd_sc_hd__nand2_1
XANTENNA__07511__B1 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_438 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10936_ fanout30/X _09745_/B _10574_/B fanout27/X vssd1 vssd1 vccd1 vccd1 _10937_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_128_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10867_ _10619_/Y _10861_/B _10866_/A vssd1 vssd1 vccd1 vccd1 _10868_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_14_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12606_ _12592_/B _12600_/B _12623_/A vssd1 vssd1 vccd1 vccd1 _12607_/D sky130_fd_sc_hd__o21ai_1
XFILLER_0_85_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10798_ _10799_/B _10799_/C _10959_/A vssd1 vssd1 vccd1 vccd1 _10800_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_121_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12537_ _12537_/A _12537_/B _12537_/C vssd1 vssd1 vccd1 vccd1 _12538_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_81_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_45 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06941__A _12626_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12468_ _12474_/B _12468_/B vssd1 vssd1 vccd1 vccd1 new_PC[3] sky130_fd_sc_hd__and2_4
XFILLER_0_53_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11419_ _11209_/X _11316_/A _11316_/B vssd1 vssd1 vccd1 vccd1 _11420_/A sky130_fd_sc_hd__a21boi_1
X_12399_ _13312_/Q _12399_/B vssd1 vssd1 vccd1 vccd1 _12399_/X sky130_fd_sc_hd__or2_1
XFILLER_0_111_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11374__B2 _09614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11374__A1 _09613_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07042__A2 _09666_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06960_ _07080_/A _07036_/A _06960_/C _09147_/S vssd1 vssd1 vccd1 vccd1 _06964_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_0_39_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06891_ _12788_/A _12790_/B vssd1 vssd1 vccd1 vccd1 _06891_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_55_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07772__A _11385_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08630_ _08646_/B2 _08661_/A2 _08673_/B _07752_/B vssd1 vssd1 vccd1 vccd1 _08631_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_55_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11294__A _11294_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08561_ _08567_/A _08567_/B vssd1 vssd1 vccd1 vccd1 _08561_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_77_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07512_ _12264_/B _07512_/B vssd1 vssd1 vccd1 vccd1 _07514_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08492_ _08492_/A _08492_/B vssd1 vssd1 vccd1 vccd1 _08494_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_92_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07443_ _09716_/A _07443_/B vssd1 vssd1 vccd1 vccd1 _07445_/B sky130_fd_sc_hd__xor2_1
Xfanout17 _12852_/A vssd1 vssd1 vccd1 vccd1 _12316_/A sky130_fd_sc_hd__clkbuf_8
Xfanout28 _07017_/X vssd1 vssd1 vccd1 vccd1 _07688_/B sky130_fd_sc_hd__buf_6
XFILLER_0_9_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout39 _12836_/A vssd1 vssd1 vccd1 vccd1 _10930_/B sky130_fd_sc_hd__buf_4
XFILLER_0_9_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout149_A _08724_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09113_ _09109_/X _09112_/X _09663_/S vssd1 vssd1 vccd1 vccd1 _09113_/X sky130_fd_sc_hd__mux2_1
XANTENNA__13051__A1 _10707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07374_ _07374_/A _07374_/B vssd1 vssd1 vccd1 vccd1 _07376_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_17_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09044_ _09032_/B _09036_/Y _09042_/Y _09043_/X _09041_/X vssd1 vssd1 vccd1 vccd1
+ _09045_/B sky130_fd_sc_hd__o311a_1
XFILLER_0_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07947__A _11384_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11365__A1 _11751_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11365__B2 _11766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08230__A1 fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08230__B2 _08304_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09946_ _09946_/A _09946_/B vssd1 vssd1 vccd1 vccd1 _09949_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__12314__B1 fanout4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08533__A2 _09567_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09877_ _09878_/A _09878_/B vssd1 vssd1 vccd1 vccd1 _09877_/X sky130_fd_sc_hd__and2_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08828_ _08829_/A _08829_/B vssd1 vssd1 vccd1 vccd1 _08864_/A sky130_fd_sc_hd__and2b_1
X_08759_ _08759_/A _08759_/B vssd1 vssd1 vccd1 vccd1 _08761_/B sky130_fd_sc_hd__xnor2_1
XTAP_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11770_ _11770_/A _11770_/B vssd1 vssd1 vccd1 vccd1 _11772_/C sky130_fd_sc_hd__xnor2_1
XTAP_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10721_ _10586_/A _10586_/B _10584_/Y vssd1 vssd1 vccd1 vccd1 _10724_/A sky130_fd_sc_hd__o21ai_2
XTAP_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10652_ _10113_/A _10651_/Y _10650_/X vssd1 vssd1 vccd1 vccd1 _10652_/Y sky130_fd_sc_hd__o21ai_1
X_13371_ _13371_/CLK _13371_/D vssd1 vssd1 vccd1 vccd1 hold254/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10583_ _10583_/A _10583_/B vssd1 vssd1 vccd1 vccd1 _10585_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_106_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12322_ _12321_/B _12322_/B vssd1 vssd1 vccd1 vccd1 _12323_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_23_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12253_ _06606_/A _12251_/X _12252_/X vssd1 vssd1 vccd1 vccd1 _12253_/Y sky130_fd_sc_hd__a21boi_1
XANTENNA__09549__B2 fanout23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11204_ _11205_/A _11205_/B vssd1 vssd1 vccd1 vccd1 _11315_/A sky130_fd_sc_hd__nand2_1
X_12184_ _12182_/Y _12184_/B vssd1 vssd1 vccd1 vccd1 _12185_/B sky130_fd_sc_hd__nand2b_1
X_11135_ _11443_/B vssd1 vssd1 vccd1 vccd1 _11135_/Y sky130_fd_sc_hd__inv_2
X_11066_ _10418_/A fanout15/X fanout36/X _09745_/B vssd1 vssd1 vccd1 vccd1 _11067_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08524__A2 _08739_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10017_ _10019_/A _10019_/B vssd1 vssd1 vccd1 vccd1 _10017_/X sky130_fd_sc_hd__or2_1
XANTENNA__11659__A2 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10331__A2 _07688_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11968_ hold192/A _12434_/B1 _12043_/B _11968_/B1 vssd1 vssd1 vccd1 vccd1 _11969_/B
+ sky130_fd_sc_hd__a31o_1
X_11899_ _11624_/A _11880_/Y _11887_/X _11898_/X vssd1 vssd1 vccd1 vccd1 _11899_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_74_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10919_ _10574_/A fanout48/X _11923_/A _10575_/A vssd1 vssd1 vccd1 vccd1 _10920_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_27_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08460__A1 _08723_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07090_ _09746_/A _07090_/B vssd1 vssd1 vccd1 vccd1 _07090_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08460__B2 _07885_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07015__A2 _09351_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout218 _06891_/Y vssd1 vssd1 vccd1 vccd1 _13236_/B sky130_fd_sc_hd__clkbuf_4
Xfanout207 _09155_/X vssd1 vssd1 vccd1 vccd1 _12307_/B1 sky130_fd_sc_hd__buf_4
Xfanout229 _06806_/Y vssd1 vssd1 vccd1 vccd1 _12794_/A sky130_fd_sc_hd__clkbuf_8
X_09800_ _09800_/A _09800_/B vssd1 vssd1 vccd1 vccd1 _09802_/B sky130_fd_sc_hd__xnor2_2
X_07992_ _07992_/A _07992_/B vssd1 vssd1 vccd1 vccd1 _07993_/B sky130_fd_sc_hd__or2_1
XFILLER_0_10_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06943_ reg1_val[7] reg1_val[8] reg1_val[9] _07182_/B vssd1 vssd1 vccd1 vccd1 _07200_/B
+ sky130_fd_sc_hd__or4_2
XANTENNA__08598__A _08598_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09731_ _09732_/A _09732_/B _09732_/C vssd1 vssd1 vccd1 vccd1 _09869_/B sky130_fd_sc_hd__o21a_1
X_09662_ _09318_/X _09330_/X _09666_/S vssd1 vssd1 vccd1 vccd1 _09662_/X sky130_fd_sc_hd__mux2_1
X_06874_ _06874_/A _06874_/B _06874_/C vssd1 vssd1 vccd1 vccd1 _06874_/X sky130_fd_sc_hd__or3_1
XFILLER_0_96_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08613_ _08613_/A _08613_/B vssd1 vssd1 vccd1 vccd1 _08615_/B sky130_fd_sc_hd__nor2_1
X_09593_ _09593_/A _09593_/B vssd1 vssd1 vccd1 vccd1 _09594_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_77_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12848__A _12848_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout266_A _06882_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08544_ _08542_/Y _08544_/B vssd1 vssd1 vccd1 vccd1 _09008_/A sky130_fd_sc_hd__and2b_1
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09222__A _10449_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11283__B1 _11766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12075__A2 fanout12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08475_ _07149_/A _08436_/A _08038_/A _08739_/A1 vssd1 vssd1 vccd1 vccd1 _08476_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_65_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07426_ _07426_/A _07426_/B vssd1 vssd1 vccd1 vccd1 _07427_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_80_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09228__B1 _08216_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07357_ _07357_/A _07357_/B vssd1 vssd1 vccd1 vccd1 _07360_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09779__B2 _11294_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09779__A1 _11146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11035__B1 _10575_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09027_ _11328_/B _11328_/C _09027_/C vssd1 vssd1 vccd1 vccd1 _11521_/B sky130_fd_sc_hd__and3_1
X_07288_ _09444_/A _11989_/A _12067_/A _09236_/B2 vssd1 vssd1 vccd1 vccd1 _07289_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_103_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold250 hold298/A vssd1 vssd1 vccd1 vccd1 hold250/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold261 hold261/A vssd1 vssd1 vccd1 vccd1 hold261/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold272 hold272/A vssd1 vssd1 vccd1 vccd1 hold272/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold283 hold283/A vssd1 vssd1 vccd1 vccd1 hold283/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold294 hold294/A vssd1 vssd1 vccd1 vccd1 hold294/X sky130_fd_sc_hd__dlygate4sd3_1
X_09929_ _09929_/A _09929_/B vssd1 vssd1 vccd1 vccd1 _09931_/B sky130_fd_sc_hd__xnor2_4
X_12940_ _13184_/A _12939_/B _12877_/X vssd1 vssd1 vccd1 vccd1 _13189_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_99_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07714__B1 _09396_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12871_ hold19/X hold265/A vssd1 vssd1 vccd1 vccd1 _12871_/X sky130_fd_sc_hd__and2b_1
XANTENNA__07190__A1 _07220_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11822_ _11822_/A _11822_/B vssd1 vssd1 vccd1 vccd1 _12169_/B sky130_fd_sc_hd__or2_1
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11813__A2 _11343_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11753_ _11753_/A vssd1 vssd1 vccd1 vccd1 _11755_/A sky130_fd_sc_hd__inv_2
XFILLER_0_126_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06602__A2_N _06771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07493__A2 _12852_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10704_ _10704_/A _10704_/B vssd1 vssd1 vccd1 vccd1 _10717_/A sky130_fd_sc_hd__nand2_1
X_11684_ _11685_/A _11685_/B vssd1 vssd1 vccd1 vccd1 _11772_/B sky130_fd_sc_hd__and2_1
XFILLER_0_125_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10635_ _10636_/A _10636_/B _10636_/C vssd1 vssd1 vccd1 vccd1 _10635_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_83_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13354_ _13355_/CLK _13354_/D vssd1 vssd1 vccd1 vccd1 hold294/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12305_ _12434_/B1 _12355_/B hold169/A vssd1 vssd1 vccd1 vccd1 _12305_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_106_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10566_ _10566_/A _10566_/B vssd1 vssd1 vccd1 vccd1 _10569_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_23_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13285_ _13285_/CLK _13285_/D vssd1 vssd1 vccd1 vccd1 hold238/A sky130_fd_sc_hd__dfxtp_1
X_10497_ _09952_/A _09952_/B _10496_/X vssd1 vssd1 vccd1 vccd1 _10499_/B sky130_fd_sc_hd__o21bai_2
XFILLER_0_51_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12236_ _06846_/A _12234_/Y _12235_/Y vssd1 vssd1 vccd1 vccd1 _12236_/X sky130_fd_sc_hd__o21a_1
X_12167_ _12280_/A _12167_/B vssd1 vssd1 vccd1 vccd1 _12170_/B sky130_fd_sc_hd__xnor2_2
X_11118_ _11118_/A _11118_/B vssd1 vssd1 vccd1 vccd1 _11118_/X sky130_fd_sc_hd__or2_1
XANTENNA__10552__A2 fanout16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12098_ _12098_/A _12098_/B _12228_/A vssd1 vssd1 vccd1 vccd1 _12099_/B sky130_fd_sc_hd__and3_1
XFILLER_0_127_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11049_ _11196_/A _11049_/B vssd1 vssd1 vccd1 vccd1 _11061_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_36_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11572__A _12317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06590_ instruction[25] _06694_/B vssd1 vssd1 vccd1 vccd1 _12626_/B sky130_fd_sc_hd__and2_4
XFILLER_0_46_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07484__A2 _10941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08260_ _08330_/A _08330_/B vssd1 vssd1 vccd1 vccd1 _08280_/A sky130_fd_sc_hd__nor2_1
X_07211_ _10589_/A _12830_/A _08507_/B _12832_/A vssd1 vssd1 vccd1 vccd1 _07212_/B
+ sky130_fd_sc_hd__o22a_1
X_08191_ _08723_/B1 fanout87/X fanout82/X _07885_/B vssd1 vssd1 vccd1 vccd1 _08192_/B
+ sky130_fd_sc_hd__o22a_1
X_07142_ _07144_/A _07142_/B _07142_/C _07142_/D vssd1 vssd1 vccd1 vccd1 _07142_/Y
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_6_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08433__A1 _08722_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07073_ _07074_/B _07074_/C _07074_/A vssd1 vssd1 vccd1 vccd1 _08391_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_70_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07944__B1 _08436_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11740__B2 _11847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11740__A1 _11923_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07975_ _07975_/A _07975_/B vssd1 vssd1 vccd1 vccd1 _08027_/B sky130_fd_sc_hd__xnor2_2
X_06926_ _06926_/A instruction[4] vssd1 vssd1 vccd1 vccd1 _09170_/B sky130_fd_sc_hd__nand2_4
X_09714_ _10928_/A _09714_/B vssd1 vssd1 vccd1 vccd1 _09718_/A sky130_fd_sc_hd__xnor2_1
X_06857_ _06846_/A _12233_/B _06840_/Y vssd1 vssd1 vccd1 vccd1 _06857_/Y sky130_fd_sc_hd__a21boi_1
X_09645_ _09647_/A _09647_/B vssd1 vssd1 vccd1 vccd1 _09645_/X sky130_fd_sc_hd__or2_2
X_06788_ reg1_val[3] _11118_/A vssd1 vssd1 vccd1 vccd1 _06788_/X sky130_fd_sc_hd__and2_1
X_09576_ _12846_/A _10167_/A1 _10022_/B1 _12848_/A vssd1 vssd1 vccd1 vccd1 _09577_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09449__B1 _08216_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08527_ _08723_/B1 _08661_/A2 _08727_/B1 _12808_/A vssd1 vssd1 vccd1 vccd1 _08528_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_77_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08458_ _08459_/A _08459_/B vssd1 vssd1 vccd1 vccd1 _08489_/A sky130_fd_sc_hd__nor2_1
X_07409_ _07409_/A _07409_/B vssd1 vssd1 vccd1 vccd1 _07413_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_107_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08389_ _09897_/A _08389_/B vssd1 vssd1 vccd1 vccd1 _08394_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__11559__A1 _11558_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10420_ _10419_/B _10419_/C _11172_/A vssd1 vssd1 vccd1 vccd1 _10424_/B sky130_fd_sc_hd__a21o_1
XANTENNA__07227__A2 _12834_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07200__A _07200_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10351_ _10352_/A _10352_/B vssd1 vssd1 vccd1 vccd1 _10351_/Y sky130_fd_sc_hd__nor2_1
X_13070_ hold116/X _12791_/A _13080_/B1 hold107/X _13113_/A vssd1 vssd1 vccd1 vccd1
+ hold117/A sky130_fd_sc_hd__o221a_1
X_10282_ _11261_/A _10282_/B vssd1 vssd1 vccd1 vccd1 _10284_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_103_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12021_ _12021_/A vssd1 vssd1 vccd1 vccd1 _12021_/Y sky130_fd_sc_hd__inv_2
XANTENNA__08727__A2 _08727_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12923_ _13114_/B _13115_/A _12903_/X vssd1 vssd1 vccd1 vccd1 _13120_/A sky130_fd_sc_hd__a21o_1
X_12854_ _12854_/A _12856_/B vssd1 vssd1 vccd1 vccd1 _12854_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_87_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11805_ hold210/A _11805_/B vssd1 vssd1 vccd1 vccd1 _11891_/B sky130_fd_sc_hd__or2_1
X_12785_ hold101/X hold166/X hold297/A hold63/X vssd1 vssd1 vccd1 vccd1 hold167/A
+ sky130_fd_sc_hd__and4_1
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08663__A1 _08730_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11736_ _12448_/S _11819_/B _11736_/C vssd1 vssd1 vccd1 vccd1 _11736_/X sky130_fd_sc_hd__or3_1
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08112__B1 _07885_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08663__B2 _07821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09860__B1 _10567_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11667_ fanout24/X _12213_/A fanout56/X _07819_/B vssd1 vssd1 vccd1 vccd1 _11668_/B
+ sky130_fd_sc_hd__o22a_1
X_10618_ _10100_/A _10100_/B _10617_/X vssd1 vssd1 vccd1 vccd1 _10618_/Y sky130_fd_sc_hd__o21bai_2
X_11598_ _11598_/A _11598_/B vssd1 vssd1 vccd1 vccd1 _11601_/A sky130_fd_sc_hd__xor2_1
X_13337_ _13340_/CLK _13337_/D vssd1 vssd1 vccd1 vccd1 hold126/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10549_ _10549_/A _10549_/B vssd1 vssd1 vccd1 vccd1 _10551_/B sky130_fd_sc_hd__xor2_2
X_13268_ _13365_/CLK hold26/X vssd1 vssd1 vccd1 vccd1 hold25/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13199_ hold246/X _13198_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13199_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10525__A2 _12404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12219_ _12219_/A _12219_/B vssd1 vssd1 vccd1 vccd1 _12219_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_47_76 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07760_ _07759_/B _07759_/C _07759_/A vssd1 vssd1 vccd1 vccd1 _07783_/A sky130_fd_sc_hd__a21bo_1
X_06711_ reg1_val[15] _06988_/A vssd1 vssd1 vccd1 vccd1 _11244_/S sky130_fd_sc_hd__and2_1
XFILLER_0_2_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09430_ _12840_/A _10589_/A _08507_/B _12842_/A vssd1 vssd1 vccd1 vccd1 _09431_/B
+ sky130_fd_sc_hd__o22a_1
X_07691_ _07691_/A _07691_/B vssd1 vssd1 vccd1 vccd1 _07695_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_2_56 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13227__B2 _12790_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06642_ reg2_val[24] _06720_/B _06703_/B1 _06641_/Y vssd1 vssd1 vccd1 vccd1 _07140_/C
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_78_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09361_ _09347_/Y _09361_/B _09361_/C _09361_/D vssd1 vssd1 vccd1 vccd1 _09371_/B
+ sky130_fd_sc_hd__and4b_1
X_06573_ instruction[3] vssd1 vssd1 vccd1 vccd1 _06926_/A sky130_fd_sc_hd__inv_2
X_09292_ _09292_/A _09292_/B vssd1 vssd1 vccd1 vccd1 _09294_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__07004__B _07064_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08312_ fanout99/X _08727_/A2 _08727_/B1 _12818_/A vssd1 vssd1 vccd1 vccd1 _08313_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08103__B1 _11558_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_12 reg1_val[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_23 reg2_val[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10461__A1 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08243_ _08244_/A _08244_/B vssd1 vssd1 vccd1 vccd1 _08248_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_28_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_34 reg2_val[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout131_A _09567_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_45 reg1_val[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_56 reg1_val[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10461__B2 _10948_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08174_ _08728_/A _08174_/B vssd1 vssd1 vccd1 vccd1 _08215_/A sky130_fd_sc_hd__xnor2_1
X_07125_ reg1_val[2] _07125_/B vssd1 vssd1 vccd1 vccd1 _07127_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_15_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07056_ _07057_/A _07057_/B vssd1 vssd1 vccd1 vccd1 _07107_/A sky130_fd_sc_hd__and2_1
XANTENNA__07955__A _07955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09382__A2 _12812_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12269__A2 _12317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07958_ _08798_/B2 _07087_/A _07087_/B _08752_/B _07821_/A vssd1 vssd1 vccd1 vccd1
+ _07959_/B sky130_fd_sc_hd__o32a_1
X_06909_ instruction[21] _06921_/B vssd1 vssd1 vccd1 vccd1 _06909_/X sky130_fd_sc_hd__or2_1
XFILLER_0_97_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07145__B2 _07144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07889_ _07889_/A _07889_/B _07889_/C vssd1 vssd1 vccd1 vccd1 _07890_/B sky130_fd_sc_hd__and3_1
XANTENNA__13218__B2 _12790_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09628_ _09628_/A _09628_/B vssd1 vssd1 vccd1 vccd1 _09629_/B sky130_fd_sc_hd__nor2_1
XANTENNA_fanout44_A _12840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09559_ _09559_/A _09559_/B vssd1 vssd1 vccd1 vccd1 _09560_/B sky130_fd_sc_hd__nor2_2
X_12570_ _12575_/B _12570_/B vssd1 vssd1 vccd1 vccd1 new_PC[18] sky130_fd_sc_hd__and2_4
XFILLER_0_65_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09410__A _09411_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11521_ _11792_/A _11521_/B _11521_/C vssd1 vssd1 vccd1 vccd1 _11523_/A sky130_fd_sc_hd__or3_1
XFILLER_0_46_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10556__A _11172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11452_ hold292/A _11536_/C _11452_/B1 vssd1 vssd1 vccd1 vccd1 _11452_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_123_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10403_ curr_PC[7] curr_PC[8] _10403_/C vssd1 vssd1 vccd1 vccd1 _10779_/D sky130_fd_sc_hd__and3_1
XFILLER_0_61_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11383_ _11758_/A _11383_/B vssd1 vssd1 vccd1 vccd1 _11385_/B sky130_fd_sc_hd__xnor2_1
X_13122_ hold294/X _12789_/B _13121_/X _12790_/A vssd1 vssd1 vccd1 vccd1 _13123_/B
+ sky130_fd_sc_hd__a22o_1
X_10334_ _10334_/A _10334_/B vssd1 vssd1 vccd1 vccd1 _10338_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_103_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13053_ _06986_/B _12818_/B hold163/X vssd1 vssd1 vccd1 vccd1 _13329_/D sky130_fd_sc_hd__a21boi_1
X_10265_ reg1_val[7] curr_PC[7] vssd1 vssd1 vccd1 vccd1 _10266_/B sky130_fd_sc_hd__nand2_1
XANTENNA__11387__A _11564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10196_ _10195_/A _10195_/B _10195_/C vssd1 vssd1 vccd1 vccd1 _10197_/B sky130_fd_sc_hd__a21oi_1
X_12004_ _12005_/A _12005_/B vssd1 vssd1 vccd1 vccd1 _12081_/B sky130_fd_sc_hd__nor2_1
XANTENNA__08581__B1 _08038_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12906_ hold291/A hold35/X vssd1 vssd1 vccd1 vccd1 _12907_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_88_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12837_ hold9/X _12848_/B _12836_/Y _13210_/A vssd1 vssd1 vccd1 vccd1 hold10/A sky130_fd_sc_hd__o211a_1
XFILLER_0_69_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12768_ _12768_/A _12768_/B _12768_/C vssd1 vssd1 vccd1 vccd1 _12769_/B sky130_fd_sc_hd__and3_2
X_11719_ _10774_/Y _11718_/Y _12244_/S vssd1 vssd1 vccd1 vccd1 _11719_/X sky130_fd_sc_hd__mux2_1
X_12699_ _12699_/A _12705_/A vssd1 vssd1 vccd1 vccd1 _12701_/C sky130_fd_sc_hd__nand2_1
XANTENNA__10443__A1 _10589_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10443__B2 _07208_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10746__A2 _10782_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07611__A2 _10570_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08930_ _08930_/A _08930_/B vssd1 vssd1 vccd1 vccd1 _08932_/A sky130_fd_sc_hd__xnor2_4
X_08861_ _08861_/A _08861_/B vssd1 vssd1 vccd1 vccd1 _08863_/B sky130_fd_sc_hd__xnor2_4
X_07812_ _07759_/A _07759_/B _07759_/C vssd1 vssd1 vccd1 vccd1 _07814_/B sky130_fd_sc_hd__a21oi_1
X_08792_ _08729_/Y _08736_/B _08734_/Y vssd1 vssd1 vccd1 vccd1 _08793_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_74_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07743_ _07744_/B _07744_/A vssd1 vssd1 vccd1 vccd1 _08013_/B sky130_fd_sc_hd__and2b_1
XANTENNA__13017__A _13214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06838__B _06838_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout179_A _09423_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07674_ _07674_/A _07674_/B vssd1 vssd1 vccd1 vccd1 _08942_/A sky130_fd_sc_hd__xnor2_4
X_06625_ _07343_/B reg1_val[28] vssd1 vssd1 vccd1 vccd1 _06625_/X sky130_fd_sc_hd__and2b_1
XANTENNA__12408__C1 _12407_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09413_ _09413_/A _09413_/B vssd1 vssd1 vccd1 vccd1 _09465_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_90_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11760__A _11908_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09344_ _09344_/A _09344_/B vssd1 vssd1 vccd1 vccd1 _09345_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_75_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09275_ _07075_/Y _11653_/A _08752_/B _12820_/A vssd1 vssd1 vccd1 vccd1 _09276_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_7_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10434__A1 _10664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10434__B2 _10567_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08226_ _08284_/A _08284_/B _08222_/X vssd1 vssd1 vccd1 vccd1 _08238_/B sky130_fd_sc_hd__o21ai_2
XFILLER_0_7_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10095__B _10096_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08157_ _08158_/A _08158_/B vssd1 vssd1 vccd1 vccd1 _08157_/X sky130_fd_sc_hd__or2_1
X_07108_ fanout30/X _12798_/A _07688_/B _09423_/B2 vssd1 vssd1 vccd1 vccd1 _07109_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_101_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08088_ _08739_/A1 _08744_/A2 _08564_/B _08436_/A vssd1 vssd1 vccd1 vccd1 _08089_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_100_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07039_ _11987_/A _07039_/B vssd1 vssd1 vccd1 vccd1 _07041_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_100_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10050_ _11470_/A _10050_/B vssd1 vssd1 vccd1 vccd1 _10054_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__07118__A1 _12626_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06748__B _07095_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10952_ _11076_/D _10952_/B vssd1 vssd1 vccd1 vccd1 _10954_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_97_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06877__B1 _09168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10673__A1 _07087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10883_ _10883_/A vssd1 vssd1 vccd1 vccd1 _10883_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_66_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10673__B2 fanout66/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12622_ reg1_val[27] curr_PC[27] _12622_/S vssd1 vssd1 vccd1 vccd1 _12623_/B sky130_fd_sc_hd__mux2_1
XANTENNA__08618__A1 _08671_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08618__B2 _08646_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09815__B1 _09163_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12553_ reg1_val[16] curr_PC[16] _12622_/S vssd1 vssd1 vccd1 vccd1 _12554_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_93_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11504_ _11504_/A _11504_/B vssd1 vssd1 vccd1 vccd1 _11506_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_102_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12484_ _12654_/B _12485_/B vssd1 vssd1 vccd1 vccd1 _12495_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_80_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11435_ _11435_/A vssd1 vssd1 vccd1 vccd1 _11435_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_1_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11366_ _12317_/A _11366_/B vssd1 vssd1 vccd1 vccd1 _11369_/A sky130_fd_sc_hd__xnor2_1
X_13105_ _13245_/A _13105_/B vssd1 vssd1 vccd1 vccd1 _13350_/D sky130_fd_sc_hd__and2_1
XANTENNA__06801__B1 _06799_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11297_ _11297_/A _11297_/B vssd1 vssd1 vccd1 vccd1 _11310_/A sky130_fd_sc_hd__xnor2_1
X_10317_ _10169_/B _10169_/C _10169_/A vssd1 vssd1 vccd1 vccd1 _10326_/A sky130_fd_sc_hd__a21boi_1
X_10248_ _09662_/X _09667_/X _10248_/S vssd1 vssd1 vccd1 vccd1 _10248_/X sky130_fd_sc_hd__mux2_1
X_13036_ hold5/X _12788_/A _13236_/B hold148/X _13109_/A vssd1 vssd1 vccd1 vccd1 hold149/A
+ sky130_fd_sc_hd__o221a_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06939__A _12423_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10179_ _10178_/B _10178_/C _10178_/A vssd1 vssd1 vccd1 vccd1 _10195_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_88_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07390_ _07396_/B _07396_/A vssd1 vssd1 vccd1 vccd1 _07390_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09060_ _09060_/A _09065_/B vssd1 vssd1 vccd1 vccd1 _09061_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_60_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08011_ _07783_/A _07783_/B _07782_/A vssd1 vssd1 vccd1 vccd1 _08016_/A sky130_fd_sc_hd__a21o_2
XANTENNA__07832__A2 _09609_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09585__A2 _11751_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09962_ _06782_/Y _09816_/X _06784_/B vssd1 vssd1 vccd1 vccd1 _09962_/X sky130_fd_sc_hd__o21a_1
X_08913_ _09053_/A _09056_/B _09058_/A _08085_/X _08023_/X vssd1 vssd1 vccd1 vccd1
+ _09060_/A sky130_fd_sc_hd__a32o_2
XFILLER_0_0_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout296_A _06578_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09893_ _09567_/B fanout13/X fanout6/X _07192_/Y vssd1 vssd1 vccd1 vccd1 _09894_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07899__A2 _07087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08844_ _08844_/A _08844_/B vssd1 vssd1 vccd1 vccd1 _08845_/C sky130_fd_sc_hd__and2_1
X_08775_ _08775_/A _08775_/B vssd1 vssd1 vccd1 vccd1 _08778_/A sky130_fd_sc_hd__xnor2_2
X_07726_ _08742_/A _07726_/B vssd1 vssd1 vccd1 vccd1 _07835_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__10655__A1 _11707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13181__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07657_ _07655_/Y _07703_/B _07652_/Y vssd1 vssd1 vccd1 vccd1 _07664_/B sky130_fd_sc_hd__a21oi_1
X_06608_ _06702_/A _12703_/B vssd1 vssd1 vccd1 vccd1 _06608_/Y sky130_fd_sc_hd__nor2_1
X_07588_ _07589_/A _07589_/B vssd1 vssd1 vccd1 vccd1 _07588_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_48_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09327_ _09117_/X _09119_/X _09330_/S vssd1 vssd1 vccd1 vccd1 _09327_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_62_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10818__B _12316_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10958__A2 _10797_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09258_ _09379_/B _09258_/B _09258_/C vssd1 vssd1 vccd1 vccd1 _09260_/B sky130_fd_sc_hd__and3_1
XFILLER_0_106_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09189_ _11142_/S _09187_/X _09188_/X vssd1 vssd1 vccd1 vccd1 dest_val[0] sky130_fd_sc_hd__o21ai_4
X_08209_ _08210_/A _08210_/B vssd1 vssd1 vccd1 vccd1 _08209_/X sky130_fd_sc_hd__and2_1
XANTENNA__09576__A2 _10167_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11220_ _11107_/B _11107_/C _11792_/A vssd1 vssd1 vccd1 vccd1 _11221_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__08304__A _08752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11649__B _11649_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11151_ _11303_/B _11151_/B vssd1 vssd1 vccd1 vccd1 _11191_/A sky130_fd_sc_hd__nor2_1
X_10102_ _10617_/A _10102_/B vssd1 vssd1 vccd1 vccd1 _10275_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__07339__B2 _09236_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07339__A1 _09444_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11082_ _10956_/A _10956_/B _10953_/Y vssd1 vssd1 vccd1 vccd1 _11085_/A sky130_fd_sc_hd__a21bo_1
X_10033_ _07510_/A _12366_/B _10148_/A vssd1 vssd1 vccd1 vccd1 _10036_/B sky130_fd_sc_hd__a21oi_1
X_11984_ _10780_/A _11980_/X _11981_/X _11983_/Y vssd1 vssd1 vccd1 vccd1 dest_val[23]
+ sky130_fd_sc_hd__a22o_4
XFILLER_0_105_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07511__A1 _12798_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11843__B1 fanout4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10935_ _10935_/A _10935_/B _10935_/C vssd1 vssd1 vccd1 vccd1 _10938_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_85_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07511__B2 _08671_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10866_ _10866_/A vssd1 vssd1 vccd1 vccd1 _10866_/Y sky130_fd_sc_hd__inv_2
XPHY_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12605_ _12605_/A _12605_/B _12605_/C _12605_/D vssd1 vssd1 vccd1 vccd1 _12607_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_0_94_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07275__B1 fanout66/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10797_ _11065_/A _10797_/B vssd1 vssd1 vccd1 vccd1 _10799_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_124_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12536_ _12537_/A _12537_/B _12537_/C vssd1 vssd1 vccd1 vccd1 _12544_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_53_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06941__B _09343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_max_cap261_A _09593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12467_ _12467_/A _12467_/B _12467_/C vssd1 vssd1 vccd1 vccd1 _12468_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_34_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11418_ _11511_/A _11511_/B vssd1 vssd1 vccd1 vccd1 _11606_/A sky130_fd_sc_hd__or2_2
X_12398_ hold298/A _11341_/B _12396_/X _09837_/A vssd1 vssd1 vccd1 vccd1 _12398_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__11374__A2 _12150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11349_ _09152_/Y _11247_/X _11347_/Y _11348_/X vssd1 vssd1 vccd1 vccd1 _11349_/X
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__07042__A3 _09351_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_load_slew214_A _09594_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08527__B1 _08727_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13019_ _13214_/A hold170/X vssd1 vssd1 vccd1 vccd1 hold171/A sky130_fd_sc_hd__and2_1
X_06890_ _12790_/A _12791_/B vssd1 vssd1 vccd1 vccd1 _06890_/Y sky130_fd_sc_hd__nor2_4
XFILLER_0_55_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11294__B _12214_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08560_ _08560_/A _08560_/B vssd1 vssd1 vccd1 vccd1 _08567_/B sky130_fd_sc_hd__xnor2_1
X_07511_ _12798_/A fanout9/A fanout5/X _08671_/B2 vssd1 vssd1 vccd1 vccd1 _07512_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_76_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08491_ _09018_/A _08491_/B vssd1 vssd1 vccd1 vccd1 _09017_/A sky130_fd_sc_hd__or2_1
XANTENNA__11834__B1 fanout12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07442_ fanout23/X _12808_/A _12810_/A _11171_/A vssd1 vssd1 vccd1 vccd1 _07443_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_71_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout18 _12852_/A vssd1 vssd1 vccd1 vccd1 _09568_/A sky130_fd_sc_hd__clkbuf_4
Xfanout29 fanout30/X vssd1 vssd1 vccd1 vccd1 fanout29/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_92_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07373_ _07374_/A _07374_/B vssd1 vssd1 vccd1 vccd1 _07579_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_9_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09112_ _09110_/X _09111_/X _09330_/S vssd1 vssd1 vccd1 vccd1 _09112_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_44_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07012__B _11172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout211_A _09898_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09043_ _09043_/A _09043_/B _08836_/Y _09042_/B vssd1 vssd1 vccd1 vccd1 _09043_/X
+ sky130_fd_sc_hd__or4bb_1
XFILLER_0_111_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout309_A _12341_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07018__B1 _12798_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmax_cap151 _11164_/A vssd1 vssd1 vccd1 vccd1 _10949_/A sky130_fd_sc_hd__buf_6
XANTENNA__11365__A2 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08230__A2 _08798_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10573__B1 _11269_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09945_ _09945_/A _09945_/B vssd1 vssd1 vccd1 vccd1 _09946_/B sky130_fd_sc_hd__xor2_4
XANTENNA__12314__A1 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13176__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09876_ _11261_/A _09876_/B vssd1 vssd1 vccd1 vccd1 _09878_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__12314__B2 fanout12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11485__A _12210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08827_ _08775_/A _08773_/Y _08772_/Y vssd1 vssd1 vccd1 vccd1 _08829_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_95_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08758_ _11564_/A _08758_/B vssd1 vssd1 vccd1 vccd1 _08759_/B sky130_fd_sc_hd__xnor2_1
XTAP_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08689_ _08689_/A _08689_/B _08689_/C vssd1 vssd1 vccd1 vccd1 _08690_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07709_ _12804_/A _07087_/A _07087_/B _08752_/B _09768_/A1 vssd1 vssd1 vccd1 vccd1
+ _07710_/B sky130_fd_sc_hd__o32a_1
XTAP_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10720_ _10720_/A _10720_/B vssd1 vssd1 vccd1 vccd1 _10725_/A sky130_fd_sc_hd__nand2_1
XTAP_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07203__A _10449_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13042__A2 _12788_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10651_ _10119_/S _09977_/Y _09181_/X vssd1 vssd1 vccd1 vccd1 _10651_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_63_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13370_ _13371_/CLK _13370_/D vssd1 vssd1 vccd1 vccd1 hold265/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10582_ _11261_/A _10582_/B vssd1 vssd1 vccd1 vccd1 _10583_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_106_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12321_ _12322_/B _12321_/B vssd1 vssd1 vccd1 vccd1 _12373_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_35_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06761__B _07080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12252_ _07144_/A _11343_/B _09354_/B _06606_/B _12455_/S vssd1 vssd1 vccd1 vccd1
+ _12252_/X sky130_fd_sc_hd__o221a_1
XANTENNA__09549__A2 fanout99/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08757__B1 _09396_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11203_ _11203_/A _11203_/B vssd1 vssd1 vccd1 vccd1 _11205_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_102_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12183_ reg1_val[26] curr_PC[26] vssd1 vssd1 vccd1 vccd1 _12184_/B sky130_fd_sc_hd__nand2_1
XANTENNA__10564__B1 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11134_ _10119_/S _09339_/X _09181_/X vssd1 vssd1 vccd1 vccd1 _11443_/B sky130_fd_sc_hd__o21a_1
X_11065_ _11065_/A _12412_/B vssd1 vssd1 vccd1 vccd1 _11069_/A sky130_fd_sc_hd__or2_1
X_10016_ _10016_/A _10016_/B vssd1 vssd1 vccd1 vccd1 _10019_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_116_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11967_ _12434_/B1 _12043_/B hold192/A vssd1 vssd1 vccd1 vccd1 _11969_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_86_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10918_ _11269_/A _10918_/B vssd1 vssd1 vccd1 vccd1 _10922_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_128_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11898_ _11892_/Y _11893_/X _11897_/X _11890_/X vssd1 vssd1 vccd1 vccd1 _11898_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_86_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10849_ _10850_/B _10850_/A vssd1 vssd1 vccd1 vccd1 _10849_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__06952__A _10710_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12519_ _12680_/B _12520_/B vssd1 vssd1 vccd1 vccd1 _12530_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_82_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12673__B _12673_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06671__B _12654_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08460__A2 _08732_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10555__B1 _11171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout219 _13213_/A2 vssd1 vssd1 vccd1 vccd1 _13006_/B1 sky130_fd_sc_hd__buf_4
Xfanout208 _09155_/X vssd1 vssd1 vccd1 vccd1 _12403_/A1 sky130_fd_sc_hd__clkbuf_4
X_07991_ _07991_/A _07991_/B vssd1 vssd1 vccd1 vccd1 _07997_/A sky130_fd_sc_hd__or2_1
X_06942_ reg1_val[4] reg1_val[5] reg1_val[6] _07160_/B vssd1 vssd1 vccd1 vccd1 _07182_/B
+ sky130_fd_sc_hd__or4_1
X_09730_ _09730_/A _09730_/B vssd1 vssd1 vccd1 vccd1 _09732_/C sky130_fd_sc_hd__xor2_1
X_06873_ _11332_/A _06873_/B _06873_/C _06873_/D vssd1 vssd1 vccd1 vccd1 _06874_/C
+ sky130_fd_sc_hd__or4_1
X_09661_ _09659_/X _09660_/X _10250_/S vssd1 vssd1 vccd1 vccd1 _09661_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_96_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08612_ _08612_/A _08612_/B vssd1 vssd1 vccd1 vccd1 _08613_/B sky130_fd_sc_hd__and2_1
XFILLER_0_82_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09592_ _09593_/A _09593_/B vssd1 vssd1 vccd1 vccd1 _09592_/X sky130_fd_sc_hd__or2_1
X_08543_ _08543_/A _08543_/B _08543_/C vssd1 vssd1 vccd1 vccd1 _08544_/B sky130_fd_sc_hd__nand3_1
XANTENNA__13025__A _13242_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout259_A _09442_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout161_A _08979_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11283__A1 fanout27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07023__A _12341_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08474_ _08474_/A _08474_/B _08474_/C vssd1 vssd1 vccd1 vccd1 _08474_/X sky130_fd_sc_hd__and3_1
XFILLER_0_65_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11283__B2 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13024__A2 _06892_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07425_ _07426_/A _07426_/B vssd1 vssd1 vccd1 vccd1 _07425_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__09228__A1 _12826_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09228__B2 _12828_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07239__B1 _12844_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07356_ _07355_/B _07356_/B vssd1 vssd1 vccd1 vccd1 _07357_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_45_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09779__A2 _11653_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11035__B2 fanout27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11035__A1 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07287_ _07290_/A _07290_/B vssd1 vssd1 vccd1 vccd1 _07292_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_5_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06581__B _06581_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09026_ _09026_/A _09026_/B vssd1 vssd1 vccd1 vccd1 _09027_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__10794__B1 _07282_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08739__B1 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold251 hold251/A vssd1 vssd1 vccd1 vccd1 hold251/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold262 hold262/A vssd1 vssd1 vccd1 vccd1 hold262/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold240 hold240/A vssd1 vssd1 vccd1 vccd1 hold240/X sky130_fd_sc_hd__buf_1
XFILLER_0_41_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold284 hold284/A vssd1 vssd1 vccd1 vccd1 hold284/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold295 hold295/A vssd1 vssd1 vccd1 vccd1 hold295/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold273 hold273/A vssd1 vssd1 vccd1 vccd1 hold273/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07693__A _09716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09928_ _09928_/A _09928_/B vssd1 vssd1 vccd1 vccd1 _09929_/B sky130_fd_sc_hd__nor2_2
XANTENNA_fanout74_A fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09703__A2 _09699_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07714__A1 _10148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09859_ _11180_/A _09859_/B vssd1 vssd1 vccd1 vccd1 _09863_/A sky130_fd_sc_hd__xnor2_1
X_12870_ hold254/X hold41/X vssd1 vssd1 vccd1 vccd1 _13206_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__07714__B2 _07089_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11821_ _11142_/S _11817_/X _11820_/X vssd1 vssd1 vccd1 vccd1 dest_val[21] sky130_fd_sc_hd__o21ai_4
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10559__A _12076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11752_ _11754_/A _11754_/B vssd1 vssd1 vccd1 vccd1 _11753_/A sky130_fd_sc_hd__or2_1
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10703_ _10844_/B _10702_/B _10702_/C vssd1 vssd1 vccd1 vccd1 _10704_/B sky130_fd_sc_hd__o21ai_1
X_11683_ _11772_/A _11683_/B vssd1 vssd1 vccd1 vccd1 _11685_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_125_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11026__A1 _12254_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10634_ _10513_/A _10510_/Y _10512_/B vssd1 vssd1 vccd1 vccd1 _10636_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_36_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13353_ _13355_/CLK _13353_/D vssd1 vssd1 vccd1 vccd1 hold242/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12304_ hold195/A _12304_/B vssd1 vssd1 vccd1 vccd1 _12355_/B sky130_fd_sc_hd__or2_1
X_10565_ _10959_/A _10565_/B vssd1 vssd1 vccd1 vccd1 _10566_/B sky130_fd_sc_hd__xnor2_2
X_13284_ _13285_/CLK _13284_/D vssd1 vssd1 vccd1 vccd1 hold248/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10496_ _10496_/A _10617_/A _10741_/A _10741_/B vssd1 vssd1 vccd1 vccd1 _10496_/X
+ sky130_fd_sc_hd__or4_1
XANTENNA__07650__B1 _08436_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12235_ _06846_/A _12234_/Y _11624_/A vssd1 vssd1 vccd1 vccd1 _12235_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__10537__B1 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12166_ _11870_/B _12165_/X _12164_/Y vssd1 vssd1 vccd1 vccd1 _12167_/B sky130_fd_sc_hd__o21ai_1
X_11117_ _11117_/A _11117_/B vssd1 vssd1 vccd1 vccd1 _11117_/X sky130_fd_sc_hd__xor2_1
XANTENNA__12829__A2 _12830_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06631__A_N _07169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12097_ _11945_/Y _12228_/A _12095_/X vssd1 vssd1 vccd1 vccd1 _12097_/X sky130_fd_sc_hd__a21o_1
X_11048_ _11048_/A _11048_/B vssd1 vssd1 vccd1 vccd1 _11049_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_127_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12668__B _12669_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12999_ _13013_/A hold178/X vssd1 vssd1 vccd1 vccd1 hold179/A sky130_fd_sc_hd__and2_1
XANTENNA__11349__A1_N _09152_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07210_ _07210_/A _07210_/B vssd1 vssd1 vccd1 vccd1 _07210_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__07778__A _07833_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08190_ _08189_/A _08242_/A _08200_/A vssd1 vssd1 vccd1 vccd1 _08190_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_0_125_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07141_ _07142_/B _07142_/C _07142_/D vssd1 vssd1 vccd1 vccd1 _07141_/X sky130_fd_sc_hd__and3_1
XFILLER_0_82_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07072_ _11271_/A _07072_/B vssd1 vssd1 vccd1 vccd1 _07072_/X sky130_fd_sc_hd__and2_1
XFILLER_0_23_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07944__B2 _08432_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07944__A1 _10537_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11740__A2 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07974_ _07974_/A _08890_/A vssd1 vssd1 vccd1 vccd1 _08027_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09697__A1 _09156_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06925_ instruction[6] instruction[5] vssd1 vssd1 vccd1 vccd1 _09157_/B sky130_fd_sc_hd__or2_2
X_09713_ _12808_/A fanout16/X _07282_/B _12810_/A vssd1 vssd1 vccd1 vccd1 _09714_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_93_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06856_ _12176_/A _06855_/X _06841_/X vssd1 vssd1 vccd1 vccd1 _12233_/B sky130_fd_sc_hd__a21o_1
X_09644_ _09644_/A _09644_/B vssd1 vssd1 vccd1 vccd1 _09647_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_96_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06787_ _06596_/A _06695_/A _12644_/B _06785_/X vssd1 vssd1 vccd1 vccd1 _06787_/X
+ sky130_fd_sc_hd__a31o_1
X_09575_ _09575_/A _09575_/B vssd1 vssd1 vccd1 vccd1 _09578_/A sky130_fd_sc_hd__nor2_1
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09449__B2 _09745_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09449__A1 _10418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08526_ _08530_/A _08530_/B vssd1 vssd1 vccd1 vccd1 _08526_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_38_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08457_ _08457_/A _08457_/B vssd1 vssd1 vccd1 vccd1 _08459_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_37_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07408_ _07409_/A _07409_/B vssd1 vssd1 vccd1 vccd1 _07460_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__07688__A _08752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08388_ _07885_/B _08732_/A2 _09440_/B1 _08721_/B1 vssd1 vssd1 vccd1 vccd1 _08389_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11559__A2 _12214_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10767__A0 _09527_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07339_ _09444_/A _12848_/A _10941_/B _09236_/B2 vssd1 vssd1 vccd1 vccd1 _07340_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09082__C1 _11707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10350_ _10194_/A _10193_/B _10193_/A vssd1 vssd1 vccd1 vccd1 _10352_/B sky130_fd_sc_hd__o21ba_1
XFILLER_0_33_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09009_ _10625_/B _10625_/C _10748_/C _09009_/D vssd1 vssd1 vccd1 vccd1 _10999_/B
+ sky130_fd_sc_hd__and4_1
X_10281_ _07087_/X _10574_/B _10575_/B fanout66/X vssd1 vssd1 vccd1 vccd1 _10282_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_14_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12020_ _11863_/A _11942_/A _11944_/B vssd1 vssd1 vccd1 vccd1 _12021_/A sky130_fd_sc_hd__a21oi_2
XANTENNA__10829__B1_N _10707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12922_ _12907_/B _13110_/B _12905_/X vssd1 vssd1 vccd1 vccd1 _13115_/A sky130_fd_sc_hd__a21o_1
XANTENNA__11673__A _11673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12853_ hold31/X _12856_/B _12852_/Y _13128_/A vssd1 vssd1 vccd1 vccd1 hold32/A sky130_fd_sc_hd__o211a_1
X_12784_ hold166/X hold172/X hold63/X vssd1 vssd1 vccd1 vccd1 _12784_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_95_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11804_ _11886_/A _10651_/Y _11803_/Y _06924_/X vssd1 vssd1 vccd1 vccd1 _11804_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12444__A0 _12626_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08112__A1 _10537_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11735_ curr_PC[19] _11734_/C curr_PC[20] vssd1 vssd1 vccd1 vccd1 _11736_/C sky130_fd_sc_hd__a21oi_1
XFILLER_0_56_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08112__B2 _08432_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08663__A2 _07752_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09860__B2 fanout30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11666_ _12317_/A _11666_/B vssd1 vssd1 vccd1 vccd1 _11670_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__11955__C1 _12423_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10617_ _10617_/A _10741_/A _10741_/B _10739_/A vssd1 vssd1 vccd1 vccd1 _10617_/X
+ sky130_fd_sc_hd__or4_2
XFILLER_0_52_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11597_ _11598_/A _11598_/B vssd1 vssd1 vccd1 vccd1 _11697_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_122_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13336_ _13340_/CLK hold125/X vssd1 vssd1 vccd1 vccd1 hold123/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10548_ _10549_/A _10549_/B vssd1 vssd1 vccd1 vccd1 _10720_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_122_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13267_ _13365_/CLK hold18/X vssd1 vssd1 vccd1 vccd1 hold17/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13172__B2 _13246_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12218_ _12219_/A _12219_/B vssd1 vssd1 vccd1 vccd1 _12277_/A sky130_fd_sc_hd__and2_1
XFILLER_0_20_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10479_ _10290_/A _10290_/B _10293_/A vssd1 vssd1 vccd1 vccd1 _10484_/A sky130_fd_sc_hd__o21ai_2
X_13198_ _13198_/A _13198_/B vssd1 vssd1 vccd1 vccd1 _13198_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12149_ fanout56/X fanout9/X fanout4/X _12213_/A vssd1 vssd1 vccd1 vccd1 _12214_/C
+ sky130_fd_sc_hd__o22ai_2
XANTENNA__09679__A1 _12244_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06710_ _06988_/A reg1_val[15] vssd1 vssd1 vccd1 vccd1 _06710_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_47_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07690_ _07691_/A _07691_/B vssd1 vssd1 vccd1 vccd1 _07986_/A sky130_fd_sc_hd__and2_1
XANTENNA__13227__A2 _12789_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06641_ _06695_/A _12669_/B vssd1 vssd1 vccd1 vccd1 _06641_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_2_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06572_ _06572_/A vssd1 vssd1 vccd1 vccd1 _06572_/Y sky130_fd_sc_hd__inv_2
X_09360_ _09350_/A _12402_/A0 _09354_/X _09358_/X _09359_/X vssd1 vssd1 vccd1 vccd1
+ _09361_/D sky130_fd_sc_hd__o2111a_1
XANTENNA__08103__A1 _08038_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09291_ _09291_/A _09291_/B vssd1 vssd1 vccd1 vccd1 _09292_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__07004__C _09351_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08311_ _08315_/A _08315_/B vssd1 vssd1 vccd1 vccd1 _08311_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_19_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08103__B2 _08730_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_13 reg1_val[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10997__B1 _12290_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08242_ _08242_/A _08242_/B vssd1 vssd1 vccd1 vccd1 _08244_/B sky130_fd_sc_hd__and2_1
XFILLER_0_117_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_46 reg1_val[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_35 reg2_val[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_24 reg2_val[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_57 reg1_val[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10461__A2 _12214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout124_A _12826_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_423 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08173_ _08741_/B2 _08727_/B1 _12820_/A _08727_/A2 vssd1 vssd1 vccd1 vccd1 _08174_/B
+ sky130_fd_sc_hd__o22a_1
X_07124_ _12626_/A _09343_/A _07200_/A vssd1 vssd1 vccd1 vccd1 _07125_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_88_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07055_ _07629_/A _07629_/B _07040_/Y vssd1 vssd1 vccd1 vccd1 _07057_/B sky130_fd_sc_hd__a21o_1
XANTENNA__11758__A _11758_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07955__B _09396_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11174__B1 _12213_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09662__S _09666_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07957_ _07956_/B _07956_/C _11564_/A vssd1 vssd1 vccd1 vccd1 _08030_/B sky130_fd_sc_hd__a21o_1
X_06908_ instruction[13] _06884_/Y _06907_/X _06694_/B vssd1 vssd1 vccd1 vccd1 reg1_idx[2]
+ sky130_fd_sc_hd__o211a_4
XANTENNA__12269__A3 _07263_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07888_ _07889_/B _07889_/C _07889_/A vssd1 vssd1 vccd1 vccd1 _07890_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__13218__A2 _12789_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06839_ reg1_val[28] _07343_/B vssd1 vssd1 vccd1 vccd1 _06839_/Y sky130_fd_sc_hd__nand2_1
X_09627_ _09628_/A _09628_/B vssd1 vssd1 vccd1 vccd1 _09629_/A sky130_fd_sc_hd__and2_1
X_09558_ _09558_/A _09558_/B _09558_/C vssd1 vssd1 vccd1 vccd1 _09559_/B sky130_fd_sc_hd__and3_1
XANTENNA__09898__A _09898_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08578__A_N _08584_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08509_ _08546_/A _08546_/B vssd1 vssd1 vccd1 vccd1 _08547_/A sky130_fd_sc_hd__nor2_1
XANTENNA_fanout37_A _07263_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09489_ _09953_/B _09489_/B vssd1 vssd1 vccd1 vccd1 _09542_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_65_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11520_ _11519_/A _11649_/C _12290_/A vssd1 vssd1 vccd1 vccd1 _11520_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_92_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11451_ _11450_/B _11544_/B _13300_/Q vssd1 vssd1 vccd1 vccd1 _11451_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_108_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10402_ _12290_/A _10372_/Y _10373_/X _10401_/X vssd1 vssd1 vccd1 vccd1 _10402_/X
+ sky130_fd_sc_hd__o31a_1
XANTENNA__07605__B1 _10567_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11382_ _11653_/A fanout56/X _12316_/A _08752_/B vssd1 vssd1 vccd1 vccd1 _11383_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_21_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13121_ hold242/X _13120_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13121_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_103_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10333_ _10334_/A _10334_/B vssd1 vssd1 vccd1 vccd1 _10454_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11668__A _12073_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09358__B1 _06939_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10572__A _11269_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13052_ hold152/X _12791_/A _13080_/B1 hold121/X _13113_/A vssd1 vssd1 vccd1 vccd1
+ hold163/A sky130_fd_sc_hd__o221a_1
X_10264_ reg1_val[7] curr_PC[7] vssd1 vssd1 vccd1 vccd1 _10264_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__11165__B1 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10195_ _10195_/A _10195_/B _10195_/C vssd1 vssd1 vccd1 vccd1 _10197_/A sky130_fd_sc_hd__and3_1
X_12003_ _12081_/A _12003_/B vssd1 vssd1 vccd1 vccd1 _12005_/B sky130_fd_sc_hd__or2_1
XANTENNA__08581__A1 _08730_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08581__B2 _09768_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12499__A _12664_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13209__A2 _13213_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12905_ hold35/X hold291/A vssd1 vssd1 vccd1 vccd1 _12905_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_88_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12836_ _12836_/A _12848_/B vssd1 vssd1 vccd1 vccd1 _12836_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_75_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09601__A _12264_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13090__B1 _06892_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13123__A _13128_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12767_ _12768_/B _12768_/C _12768_/A vssd1 vssd1 vccd1 vccd1 _12773_/B sky130_fd_sc_hd__a21oi_2
XANTENNA__11640__A1 _07210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11718_ _11718_/A _11718_/B vssd1 vssd1 vccd1 vccd1 _11718_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_84_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12698_ reg1_val[14] _12698_/B vssd1 vssd1 vccd1 vccd1 _12705_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_44_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10443__A2 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07121__A _12626_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11649_ _11649_/A _11649_/B _11649_/C _11649_/D vssd1 vssd1 vccd1 vccd1 _11650_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_0_24_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13319_ _13343_/CLK _13319_/D vssd1 vssd1 vccd1 vccd1 hold79/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06960__A _07080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11156__B1 _11766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08860_ _08861_/B _08861_/A vssd1 vssd1 vccd1 vccd1 _08860_/X sky130_fd_sc_hd__and2b_1
X_07811_ _07811_/A _07811_/B vssd1 vssd1 vccd1 vccd1 _07816_/A sky130_fd_sc_hd__xor2_1
X_08791_ _08743_/A _08743_/B _08748_/A vssd1 vssd1 vccd1 vccd1 _08795_/A sky130_fd_sc_hd__o21ba_1
X_07742_ _08013_/A _07742_/B vssd1 vssd1 vccd1 vccd1 _07744_/B sky130_fd_sc_hd__or2_1
XFILLER_0_74_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07673_ _07675_/A _07675_/B vssd1 vssd1 vccd1 vccd1 _07676_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_94_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06624_ reg2_val[28] _06720_/B _06703_/B1 _06623_/Y vssd1 vssd1 vccd1 vccd1 _07343_/B
+ sky130_fd_sc_hd__o2bb2a_4
X_09412_ _09413_/A _09413_/B vssd1 vssd1 vccd1 vccd1 _09633_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_87_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09343_ _09343_/A curr_PC[1] vssd1 vssd1 vccd1 vccd1 _09344_/B sky130_fd_sc_hd__or2_1
XFILLER_0_59_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08088__B1 _08564_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout241_A _09147_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11631__A1 _12394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09274_ _09272_/X _09274_/B vssd1 vssd1 vccd1 vccd1 _09277_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_47_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10434__A2 _10797_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08225_ _08225_/A _08225_/B vssd1 vssd1 vccd1 vccd1 _08284_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_15_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08156_ _08724_/A _08156_/B vssd1 vssd1 vccd1 vccd1 _08158_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__07063__A1 _07095_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07107_ _07107_/A _07107_/B vssd1 vssd1 vccd1 vccd1 _07309_/A sky130_fd_sc_hd__or2_2
XFILLER_0_31_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08087_ _08742_/A _08087_/B vssd1 vssd1 vccd1 vccd1 _08146_/A sky130_fd_sc_hd__xnor2_1
X_07038_ _12804_/A _10574_/A _09768_/A1 _10575_/A vssd1 vssd1 vccd1 vccd1 _07039_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_3_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08797__A _11385_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08989_ _08989_/A _08989_/B vssd1 vssd1 vccd1 vccd1 _09961_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__07118__A2 _09343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10951_ _10950_/A _10950_/B _10950_/C vssd1 vssd1 vccd1 vccd1 _10952_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_98_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10673__A2 _07087_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12621_ _12618_/B _12620_/B _12618_/A vssd1 vssd1 vccd1 vccd1 _12624_/A sky130_fd_sc_hd__o21ba_2
X_10882_ _10252_/S _09681_/X _10881_/X vssd1 vssd1 vccd1 vccd1 _10883_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_78_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09421__A _12798_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08618__A2 _09238_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10567__A _10567_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12552_ _12556_/B _12552_/B vssd1 vssd1 vccd1 vccd1 new_PC[15] sky130_fd_sc_hd__and2_4
XFILLER_0_93_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07826__B1 _08721_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08037__A _08733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12483_ reg1_val[6] curr_PC[6] _12622_/S vssd1 vssd1 vccd1 vccd1 _12485_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11503_ _11503_/A _11503_/B vssd1 vssd1 vccd1 vccd1 _11506_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_124_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11434_ _06707_/B _11329_/X _06705_/X vssd1 vssd1 vccd1 vccd1 _11435_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_80_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09579__B1 _10570_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11386__B1 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10506__S _12388_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11365_ _11751_/A fanout15/X fanout36/X _11766_/A vssd1 vssd1 vccd1 vccd1 _11366_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__13127__B2 _12790_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13104_ hold284/X _06892_/B _13103_/X _06572_/A vssd1 vssd1 vccd1 vccd1 _13105_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11138__B1 _11137_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11296_ _11297_/A _11297_/B vssd1 vssd1 vccd1 vccd1 _11296_/X sky130_fd_sc_hd__and2b_1
X_10316_ _10190_/A _10190_/B _10187_/A vssd1 vssd1 vccd1 vccd1 _10328_/A sky130_fd_sc_hd__o21ba_1
XFILLER_0_119_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13035_ hold5/X _13236_/B _09897_/A _13087_/B2 _13034_/Y vssd1 vssd1 vccd1 vccd1
+ hold6/A sky130_fd_sc_hd__o221a_1
X_10247_ _09660_/X _09663_/X _10250_/S vssd1 vssd1 vccd1 vccd1 _10247_/X sky130_fd_sc_hd__mux2_1
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10178_ _10178_/A _10178_/B _10178_/C vssd1 vssd1 vccd1 vccd1 _10195_/A sky130_fd_sc_hd__or3_1
XFILLER_0_28_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13118__A _13128_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12819_ hold45/X _12818_/B _12818_/Y _13245_/A vssd1 vssd1 vccd1 vccd1 hold46/A sky130_fd_sc_hd__o211a_1
XANTENNA__06674__B _07135_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08010_ _07847_/A _07847_/B _07845_/Y vssd1 vssd1 vccd1 vccd1 _08017_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__07786__A _08733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09961_ _09961_/A _09961_/B vssd1 vssd1 vccd1 vccd1 _09961_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_40_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08912_ _08912_/A _08912_/B vssd1 vssd1 vccd1 vccd1 _09065_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09892_ _10076_/B _09892_/B vssd1 vssd1 vccd1 vccd1 _09929_/A sky130_fd_sc_hd__or2_2
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout191_A _09111_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07899__A3 _07087_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08843_ _08752_/A _09614_/A _08046_/A _08811_/A vssd1 vssd1 vccd1 vccd1 _08844_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_0_109_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout289_A _06771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08774_ _08774_/A _08774_/B vssd1 vssd1 vccd1 vccd1 _08775_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07725_ _08741_/A2 _11472_/A _11558_/A _08617_/B vssd1 vssd1 vccd1 vccd1 _07726_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__06865__A _12626_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09241__A _09441_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07656_ _07656_/A _07656_/B vssd1 vssd1 vccd1 vccd1 _07703_/B sky130_fd_sc_hd__xor2_1
X_06607_ instruction[40] _06634_/B vssd1 vssd1 vccd1 vccd1 _12703_/B sky130_fd_sc_hd__and2_4
XFILLER_0_94_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07587_ _07571_/A _07571_/B _07574_/A vssd1 vssd1 vccd1 vccd1 _07589_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_47_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09326_ _09116_/X _09142_/X _09351_/B vssd1 vssd1 vccd1 vccd1 _09326_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_48_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09257_ _09257_/A _09257_/B vssd1 vssd1 vccd1 vccd1 _09258_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08208_ _08208_/A _08208_/B vssd1 vssd1 vccd1 vccd1 _08210_/B sky130_fd_sc_hd__xnor2_1
X_09188_ curr_PC[0] _10780_/A vssd1 vssd1 vccd1 vccd1 _09188_/X sky130_fd_sc_hd__or2_1
XFILLER_0_62_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11649__C _11649_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08233__B1 _07955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08139_ _08139_/A _08139_/B vssd1 vssd1 vccd1 vccd1 _08213_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_113_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08304__B _08304_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11150_ _11150_/A _11150_/B vssd1 vssd1 vccd1 vccd1 _11151_/B sky130_fd_sc_hd__and2_1
XFILLER_0_101_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10101_ _09489_/B _10097_/X _10100_/Y vssd1 vssd1 vccd1 vccd1 _10102_/B sky130_fd_sc_hd__o21a_1
XANTENNA__07339__A2 _12848_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11081_ _11081_/A _11081_/B vssd1 vssd1 vccd1 vccd1 _11086_/A sky130_fd_sc_hd__nand2_1
X_10032_ _10032_/A vssd1 vssd1 vccd1 vccd1 _10042_/A sky130_fd_sc_hd__inv_2
Xclkbuf_4_4_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13299_/CLK sky130_fd_sc_hd__clkbuf_8
X_11983_ _12448_/S _12058_/B vssd1 vssd1 vccd1 vccd1 _11983_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_86_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07511__A2 fanout9/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11843__B2 _11923_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11843__A1 _11989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10934_ _10938_/A vssd1 vssd1 vccd1 vccd1 _11076_/A sky130_fd_sc_hd__inv_2
XFILLER_0_39_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10865_ _10613_/X _10735_/X _10736_/X vssd1 vssd1 vccd1 vccd1 _10866_/A sky130_fd_sc_hd__a21oi_1
XPHY_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12604_ _12623_/A _12604_/B vssd1 vssd1 vccd1 vccd1 _12608_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_121_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12535_ _12544_/A _12535_/B vssd1 vssd1 vccd1 vccd1 _12537_/C sky130_fd_sc_hd__nand2_1
XANTENNA__07275__A1 _11653_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10796_ _07510_/A _12366_/B _07178_/Y vssd1 vssd1 vccd1 vccd1 _10799_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_26_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08472__B1 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07275__B2 _10413_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12466_ _12467_/A _12467_/B _12467_/C vssd1 vssd1 vccd1 vccd1 _12474_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_81_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11359__B1 _11142_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12397_ _11341_/B _12396_/X hold298/A vssd1 vssd1 vccd1 vccd1 _12397_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_105_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11417_ _11417_/A _11417_/B _11417_/C vssd1 vssd1 vccd1 vccd1 _11511_/B sky130_fd_sc_hd__and3_1
X_11348_ hold174/A _11450_/B _11449_/B _11968_/B1 vssd1 vssd1 vccd1 vccd1 _11348_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_39_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06786__B1 _06785_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12308__C1 _12404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08527__A1 _08723_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11279_ _12073_/A _11279_/B vssd1 vssd1 vccd1 vccd1 _11280_/B sky130_fd_sc_hd__xnor2_1
X_13018_ hold169/X _13213_/B2 _13213_/A2 _13312_/Q vssd1 vssd1 vccd1 vccd1 hold170/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08527__B2 _12808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07510_ _07510_/A _12366_/B vssd1 vssd1 vccd1 vccd1 fanout5/A sky130_fd_sc_hd__and2_1
XFILLER_0_71_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08490_ _09018_/A _08491_/B vssd1 vssd1 vccd1 vccd1 _08490_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__11834__A1 fanout24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11834__B2 _07819_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout19 _07154_/X vssd1 vssd1 vccd1 vccd1 _12852_/A sky130_fd_sc_hd__buf_4
X_07441_ _09548_/A _07441_/B vssd1 vssd1 vccd1 vccd1 _07445_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_29_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07372_ _07174_/A _07174_/B _07172_/Y vssd1 vssd1 vccd1 vccd1 _07374_/B sky130_fd_sc_hd__a21o_1
X_09111_ reg1_val[8] reg1_val[23] _09111_/S vssd1 vssd1 vccd1 vccd1 _09111_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_91_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_112 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07012__C _07013_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09042_ _09042_/A _09042_/B vssd1 vssd1 vccd1 vccd1 _09042_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_103_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07018__B2 _07688_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07018__A1 _08671_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11471__A2_N fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10022__B1 _10022_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11766__A _11766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09944_ _09945_/A _09945_/B vssd1 vssd1 vccd1 vccd1 _09944_/X sky130_fd_sc_hd__and2_1
XFILLER_0_0_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09715__B1 _10818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09875_ _11294_/A _07087_/A _07087_/B fanout66/X _10418_/A vssd1 vssd1 vccd1 vccd1
+ _09876_/B sky130_fd_sc_hd__o32a_1
XANTENNA__12314__A2 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08826_ _08826_/A _08826_/B vssd1 vssd1 vccd1 vccd1 _08829_/A sky130_fd_sc_hd__xnor2_2
X_08757_ _08798_/B2 _09609_/B _09396_/B _07821_/A vssd1 vssd1 vccd1 vccd1 _08758_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08688_ _08670_/B _08987_/B _08668_/X vssd1 vssd1 vccd1 vccd1 _08989_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_67_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07708_ _11385_/A _07708_/B vssd1 vssd1 vccd1 vccd1 _07712_/A sky130_fd_sc_hd__xnor2_1
XTAP_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07639_ _12076_/A _07639_/B vssd1 vssd1 vccd1 vccd1 _07642_/A sky130_fd_sc_hd__xnor2_1
X_10650_ _10642_/Y _10643_/X _10648_/X _10649_/Y vssd1 vssd1 vccd1 vccd1 _10650_/X
+ sky130_fd_sc_hd__o211a_1
X_09309_ _09190_/X _09542_/B _12290_/A vssd1 vssd1 vccd1 vccd1 _09309_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_35_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10581_ fanout66/X fanout48/X _10930_/B _07087_/X vssd1 vssd1 vccd1 vccd1 _10582_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_91_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12320_ _12320_/A _12320_/B vssd1 vssd1 vccd1 vccd1 _12322_/B sky130_fd_sc_hd__or2_1
XFILLER_0_106_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12251_ _06606_/B _09158_/Y _09154_/Y vssd1 vssd1 vccd1 vccd1 _12251_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_44_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08757__B2 _07821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08757__A1 _08798_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10013__B1 _10570_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11202_ _11203_/A _11203_/B vssd1 vssd1 vccd1 vccd1 _11311_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_102_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12182_ reg1_val[26] curr_PC[26] vssd1 vssd1 vccd1 vccd1 _12182_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_31_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10564__A1 _10818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10564__B2 _10664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11133_ _11128_/Y _11129_/X _11132_/Y _11126_/X vssd1 vssd1 vccd1 vccd1 _11133_/X
+ sky130_fd_sc_hd__o211a_1
X_11064_ _12261_/A _11064_/B vssd1 vssd1 vccd1 vccd1 _11070_/A sky130_fd_sc_hd__xnor2_1
X_10015_ _10016_/A _10016_/B vssd1 vssd1 vccd1 vccd1 _10015_/X sky130_fd_sc_hd__or2_1
XFILLER_0_116_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12069__A1 _11989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11966_ hold225/A _11966_/B vssd1 vssd1 vccd1 vccd1 _12043_/B sky130_fd_sc_hd__or2_1
XANTENNA__11816__A1 _11624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13018__B1 _13213_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10917_ _10570_/A _12150_/A fanout59/X _10571_/A vssd1 vssd1 vccd1 vccd1 _10918_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_128_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11897_ _10113_/A _10516_/Y _10528_/Y _12254_/A1 _11896_/X vssd1 vssd1 vccd1 vccd1
+ _11897_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_128_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10848_ _10848_/A _10848_/B vssd1 vssd1 vccd1 vccd1 _10850_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_26_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10779_ curr_PC[9] curr_PC[10] curr_PC[11] _10779_/D vssd1 vssd1 vccd1 vccd1 _10906_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_0_54_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06952__B _06954_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11044__A2 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12518_ reg1_val[11] curr_PC[11] _12622_/S vssd1 vssd1 vccd1 vccd1 _12520_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_26_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12449_ _12629_/B _12450_/B vssd1 vssd1 vccd1 vccd1 _12460_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_2_724 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10555__A1 _10418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10555__B2 _09745_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout209 _09081_/X vssd1 vssd1 vccd1 vccd1 _12290_/A sky130_fd_sc_hd__buf_4
X_07990_ _07990_/A _07990_/B vssd1 vssd1 vccd1 vccd1 _07991_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_1_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06941_ _12626_/A _09343_/A reg1_val[2] reg1_val[3] vssd1 vssd1 vccd1 vccd1 _07160_/B
+ sky130_fd_sc_hd__or4_2
XFILLER_0_5_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09660_ _09314_/X _09322_/X _09666_/S vssd1 vssd1 vccd1 vccd1 _09660_/X sky130_fd_sc_hd__mux2_1
X_06872_ _06872_/A _06872_/B vssd1 vssd1 vccd1 vccd1 _06873_/D sky130_fd_sc_hd__nand2_1
XANTENNA__07184__B1 _07200_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08611_ _08611_/A _08611_/B vssd1 vssd1 vccd1 vccd1 _08625_/A sky130_fd_sc_hd__xnor2_2
X_09591_ _09898_/A _09591_/B vssd1 vssd1 vccd1 vccd1 _09593_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08542_ _08543_/B _08543_/C _08543_/A vssd1 vssd1 vccd1 vccd1 _08542_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__12210__A _12210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08473_ _10444_/A _08473_/B vssd1 vssd1 vccd1 vccd1 _08474_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_49_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11283__A2 _11847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07424_ _09441_/A _07424_/B vssd1 vssd1 vccd1 vccd1 _07426_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_15_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07023__B _07064_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09228__A2 fanout69/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07239__B2 _09444_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07239__A1 _12846_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07355_ _07356_/B _07355_/B vssd1 vssd1 vccd1 vccd1 _07357_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__11035__A2 _11558_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10243__B1 _11624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07286_ _09442_/A _07286_/B vssd1 vssd1 vccd1 vccd1 _07290_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_45_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09025_ _08426_/A _08426_/B _09020_/X _09024_/X vssd1 vssd1 vccd1 vccd1 _09026_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10794__B2 _11294_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10794__A1 _11146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08739__B2 _08436_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08739__A1 _08739_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_362 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold252 hold252/A vssd1 vssd1 vccd1 vccd1 hold252/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold230 hold232/X vssd1 vssd1 vccd1 vccd1 hold230/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold241 hold241/A vssd1 vssd1 vccd1 vccd1 hold241/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold263 hold263/A vssd1 vssd1 vccd1 vccd1 hold263/X sky130_fd_sc_hd__buf_1
Xhold285 hold285/A vssd1 vssd1 vccd1 vccd1 hold285/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold274 hold274/A vssd1 vssd1 vccd1 vccd1 hold274/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold296 hold296/A vssd1 vssd1 vccd1 vccd1 hold296/X sky130_fd_sc_hd__dlygate4sd3_1
X_09927_ _09927_/A _09927_/B vssd1 vssd1 vccd1 vccd1 _09928_/B sky130_fd_sc_hd__and2_1
XANTENNA__07714__A2 _09609_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09858_ _11065_/A _10574_/A _10575_/A _11146_/A vssd1 vssd1 vccd1 vccd1 _09859_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07175__B1 _08732_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13248__B1 _13242_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09789_ _09789_/A _09789_/B vssd1 vssd1 vccd1 vccd1 _09790_/B sky130_fd_sc_hd__nand2_1
X_08809_ _08809_/A _08809_/B vssd1 vssd1 vccd1 vccd1 _08811_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_68_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11820_ _12448_/S _11820_/B _11982_/C vssd1 vssd1 vccd1 vccd1 _11820_/X sky130_fd_sc_hd__or3_1
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11751_ _11751_/A _12214_/B _11661_/A vssd1 vssd1 vccd1 vccd1 _11754_/B sky130_fd_sc_hd__or3b_1
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10702_ _10844_/B _10702_/B _10702_/C vssd1 vssd1 vccd1 vccd1 _10704_/A sky130_fd_sc_hd__or3_1
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11682_ _11682_/A _11682_/B _11682_/C vssd1 vssd1 vccd1 vccd1 _11683_/B sky130_fd_sc_hd__and3_1
XFILLER_0_126_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11026__A2 _11012_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10633_ reg1_val[10] curr_PC[10] vssd1 vssd1 vccd1 vccd1 _10636_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_48_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10575__A _10575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13352_ _13355_/CLK _13352_/D vssd1 vssd1 vccd1 vccd1 hold258/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10564_ _10818_/A _10797_/B fanout5/X _10664_/A vssd1 vssd1 vccd1 vccd1 _10565_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_23_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12303_ hold266/A _11341_/B _12352_/B _12302_/Y _09837_/A vssd1 vssd1 vccd1 vccd1
+ _12303_/X sky130_fd_sc_hd__a311o_1
XANTENNA__06989__B1 _10948_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13283_ _13285_/CLK _13283_/D vssd1 vssd1 vccd1 vccd1 hold290/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12790__A _12790_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10495_ _10741_/A _10233_/X _10741_/B _10494_/X vssd1 vssd1 vccd1 vccd1 _10499_/A
+ sky130_fd_sc_hd__o31a_1
XANTENNA__07650__A1 _07149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07650__B2 _12067_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12234_ _12423_/A _12195_/S _12176_/Y _12233_/Y vssd1 vssd1 vccd1 vccd1 _12234_/Y
+ sky130_fd_sc_hd__o31ai_1
XFILLER_0_32_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10537__B2 _10706_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10537__A1 _10537_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12165_ _12165_/A _12165_/B _12281_/A vssd1 vssd1 vccd1 vccd1 _12165_/X sky130_fd_sc_hd__or3_1
X_11116_ _11009_/A _11009_/B _11007_/B vssd1 vssd1 vccd1 vccd1 _11117_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_127_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12096_ _12165_/B _12162_/A vssd1 vssd1 vccd1 vccd1 _12228_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_36_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11047_ _11048_/A _11048_/B vssd1 vssd1 vccd1 vccd1 _11196_/A sky130_fd_sc_hd__nor2_1
X_12998_ hold200/A _13004_/A2 _13006_/B1 hold177/X vssd1 vssd1 vccd1 vccd1 hold178/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12965__A _13214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11949_ _12165_/B _11949_/B vssd1 vssd1 vccd1 vccd1 _11985_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__06963__A _06963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06682__B _07210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07140_ _07169_/A _07140_/B _07140_/C vssd1 vssd1 vccd1 vccd1 _07142_/D sky130_fd_sc_hd__and3_1
XFILLER_0_55_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10776__A1 _09172_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07071_ _11163_/A _07071_/B _07071_/C _07071_/D vssd1 vssd1 vccd1 vccd1 _07072_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_2_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07944__A2 _08739_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09712_ _09597_/A _09597_/B _09595_/Y vssd1 vssd1 vccd1 vccd1 _09726_/A sky130_fd_sc_hd__a21o_2
X_07973_ _07974_/A _07973_/B _07973_/C vssd1 vssd1 vccd1 vccd1 _08890_/A sky130_fd_sc_hd__nand3_1
XANTENNA__07157__B1 _07200_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06924_ instruction[6] instruction[5] _09165_/A vssd1 vssd1 vccd1 vccd1 _06924_/X
+ sky130_fd_sc_hd__or3_4
X_06855_ _12110_/A _06854_/X _06842_/X vssd1 vssd1 vccd1 vccd1 _06855_/X sky130_fd_sc_hd__a21o_1
X_09643_ _09643_/A _09643_/B vssd1 vssd1 vccd1 vccd1 _09644_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_117_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09574_ _09573_/A _09573_/B _09573_/C vssd1 vssd1 vccd1 vccd1 _09575_/B sky130_fd_sc_hd__a21oi_1
X_06786_ _06596_/A _06695_/A _12644_/B _06785_/X vssd1 vssd1 vccd1 vccd1 _07044_/A
+ sky130_fd_sc_hd__a31oi_4
XFILLER_0_89_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08525_ _08681_/A _08525_/B vssd1 vssd1 vccd1 vccd1 _08530_/B sky130_fd_sc_hd__xnor2_1
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09449__A2 fanout69/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08456_ _08456_/A _08456_/B vssd1 vssd1 vccd1 vccd1 _08459_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_80_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07407_ _07485_/A _07407_/B vssd1 vssd1 vccd1 vccd1 _07409_/B sky130_fd_sc_hd__xnor2_1
X_08387_ _08387_/A _08387_/B vssd1 vssd1 vccd1 vccd1 _08419_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_46_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07688__B _07688_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07338_ _07338_/A vssd1 vssd1 vccd1 vccd1 _07363_/A sky130_fd_sc_hd__inv_2
XFILLER_0_18_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10767__A1 _09354_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07269_ _07269_/A _07269_/B vssd1 vssd1 vccd1 vccd1 _07672_/A sky130_fd_sc_hd__xnor2_2
X_09008_ _09008_/A _09008_/B vssd1 vssd1 vccd1 vccd1 _09009_/D sky130_fd_sc_hd__xnor2_1
X_10280_ _11470_/A _10280_/B vssd1 vssd1 vccd1 vccd1 _10284_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_13_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12921_ _12910_/B _13106_/B _12908_/X vssd1 vssd1 vccd1 vccd1 _13110_/B sky130_fd_sc_hd__a21o_1
XANTENNA__09424__A _12264_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06767__B _07036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12852_ _12852_/A _12856_/B vssd1 vssd1 vccd1 vccd1 _12852_/Y sky130_fd_sc_hd__nand2_1
X_12783_ hold172/X hold63/X vssd1 vssd1 vccd1 vccd1 _12783_/Y sky130_fd_sc_hd__nand2_1
X_11803_ _11886_/A _11803_/B vssd1 vssd1 vccd1 vccd1 _11803_/Y sky130_fd_sc_hd__nor2_1
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11734_ curr_PC[19] curr_PC[20] _11734_/C vssd1 vssd1 vccd1 vccd1 _11819_/B sky130_fd_sc_hd__and3_1
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08112__A2 _08723_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09860__A2 _10664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11665_ _11923_/A fanout15/X fanout36/X _11989_/A vssd1 vssd1 vccd1 vccd1 _11666_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_126_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10616_ _10741_/B _10739_/A vssd1 vssd1 vccd1 vccd1 _10616_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_37_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10207__B1 _10574_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11596_ _11596_/A _11596_/B vssd1 vssd1 vccd1 vccd1 _11598_/B sky130_fd_sc_hd__xnor2_1
X_13335_ _13340_/CLK _13335_/D vssd1 vssd1 vccd1 vccd1 hold130/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10547_ _10433_/Y _10440_/B _10438_/Y vssd1 vssd1 vccd1 vccd1 _10549_/B sky130_fd_sc_hd__a21bo_1
X_13266_ _13384_/CLK hold14/X vssd1 vssd1 vccd1 vccd1 hold13/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06977__A3 _06994_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10478_ _10353_/A _10353_/B _10351_/Y vssd1 vssd1 vccd1 vccd1 _10485_/A sky130_fd_sc_hd__a21o_1
XANTENNA__13172__A2 _06890_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08503__A _09433_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12217_ _12217_/A _12217_/B vssd1 vssd1 vccd1 vccd1 _12219_/B sky130_fd_sc_hd__xnor2_1
X_13197_ _12872_/X _13197_/B vssd1 vssd1 vccd1 vccd1 _13198_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_20_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12148_ _12148_/A _12148_/B vssd1 vssd1 vccd1 vccd1 _12153_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__06958__A _11118_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12079_ _12145_/B _12079_/B vssd1 vssd1 vccd1 vccd1 _12081_/C sky130_fd_sc_hd__nor2_1
XANTENNA__09679__A2 _09672_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12679__B _12680_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06640_ instruction[34] _06694_/B vssd1 vssd1 vccd1 vccd1 _12669_/B sky130_fd_sc_hd__and2_4
XFILLER_0_63_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06571_ hold296/X vssd1 vssd1 vccd1 vccd1 _06571_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_59_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09290_ _07516_/Y _07520_/A _09291_/B vssd1 vssd1 vccd1 vccd1 _09290_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_47_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08310_ _08731_/A _08310_/B vssd1 vssd1 vccd1 vccd1 _08315_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_19_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10446__B1 _10706_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08103__A2 _11472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_14 reg1_val[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08241_ _08241_/A _08241_/B vssd1 vssd1 vccd1 vccd1 _08242_/B sky130_fd_sc_hd__nand2_1
XANTENNA_47 reg1_val[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12199__B1 _12190_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_25 reg2_val[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_36 _09699_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_58 reg1_val[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08172_ _08178_/A _08178_/B vssd1 vssd1 vccd1 vccd1 _08172_/X sky130_fd_sc_hd__and2_1
XFILLER_0_27_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07123_ _09343_/A _07123_/B vssd1 vssd1 vccd1 vccd1 _07123_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10943__A _11470_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07054_ _09716_/A _07054_/B vssd1 vssd1 vccd1 vccd1 _07629_/B sky130_fd_sc_hd__xnor2_2
XANTENNA_fanout117_A _08741_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11174__A1 _07087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11174__B2 fanout66/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07956_ _11564_/A _07956_/B _07956_/C vssd1 vssd1 vccd1 vccd1 _08030_/A sky130_fd_sc_hd__nand3_1
X_06907_ instruction[20] _06921_/B vssd1 vssd1 vccd1 vccd1 _06907_/X sky130_fd_sc_hd__or2_1
XANTENNA__12269__A4 _12412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07887_ _07886_/B _07886_/C _11385_/A vssd1 vssd1 vccd1 vccd1 _07889_/C sky130_fd_sc_hd__a21o_1
X_06838_ _06838_/A _06838_/B vssd1 vssd1 vccd1 vccd1 _06838_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__07550__B1 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09626_ _09626_/A _09626_/B vssd1 vssd1 vccd1 vccd1 _09628_/B sky130_fd_sc_hd__xnor2_1
X_06769_ _06769_/A _06769_/B vssd1 vssd1 vccd1 vccd1 _10109_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_78_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09557_ _09558_/A _09558_/B _09558_/C vssd1 vssd1 vccd1 vccd1 _09559_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_77_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08508_ _08508_/A _08508_/B vssd1 vssd1 vccd1 vccd1 _08546_/B sky130_fd_sc_hd__xor2_1
X_09488_ _09069_/B _09485_/X _09486_/X _09487_/X vssd1 vssd1 vccd1 vccd1 _09489_/B
+ sky130_fd_sc_hd__o211a_2
XANTENNA__07699__A _08731_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08439_ _08681_/A _08439_/B _08439_/C vssd1 vssd1 vccd1 vccd1 _08442_/B sky130_fd_sc_hd__and3_1
XFILLER_0_65_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11450_ _13300_/Q _11450_/B _11544_/B vssd1 vssd1 vccd1 vccd1 _11450_/X sky130_fd_sc_hd__and3_1
XFILLER_0_104_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10401_ _10374_/Y _10375_/X _10379_/X _10400_/X vssd1 vssd1 vccd1 vccd1 _10401_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__07605__A1 _10664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07605__B2 fanout69/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08802__B1 _09396_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11381_ _11381_/A _11381_/B vssd1 vssd1 vccd1 vccd1 _11396_/A sky130_fd_sc_hd__xor2_1
X_13120_ _13120_/A _13120_/B vssd1 vssd1 vccd1 vccd1 _13120_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_61_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10332_ _11673_/A _10332_/B vssd1 vssd1 vccd1 vccd1 _10334_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_21_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13051_ _10707_/A _12798_/B hold153/X vssd1 vssd1 vccd1 vccd1 hold154/A sky130_fd_sc_hd__a21boi_1
X_10263_ _10133_/A _10130_/Y _10132_/B vssd1 vssd1 vccd1 vccd1 _10267_/A sky130_fd_sc_hd__o21a_1
XANTENNA__11165__A1 _10941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11165__B2 fanout94/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12002_ _12002_/A _12002_/B vssd1 vssd1 vccd1 vccd1 _12003_/B sky130_fd_sc_hd__nor2_1
X_10194_ _10194_/A _10194_/B vssd1 vssd1 vccd1 vccd1 _10195_/C sky130_fd_sc_hd__xor2_1
XANTENNA__08581__A2 _12808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12904_ hold258/X hold90/X vssd1 vssd1 vccd1 vccd1 _13114_/B sky130_fd_sc_hd__nand2b_1
XTAP_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12835_ hold15/X _12848_/B _12834_/Y _13214_/A vssd1 vssd1 vccd1 vccd1 hold16/A sky130_fd_sc_hd__o211a_1
XTAP_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13090__A1 _06572_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12766_ _12766_/A _12766_/B _12766_/C vssd1 vssd1 vccd1 vccd1 _12768_/C sky130_fd_sc_hd__or3_1
XFILLER_0_126_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11640__A2 _11343_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11717_ _11627_/A _11629_/B _11627_/B vssd1 vssd1 vccd1 vccd1 _11718_/B sky130_fd_sc_hd__a21boi_1
XFILLER_0_84_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12697_ reg1_val[14] _12698_/B vssd1 vssd1 vccd1 vccd1 _12699_/A sky130_fd_sc_hd__or2_1
XFILLER_0_114_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11648_ _12448_/S _11645_/X _11646_/X _11647_/Y vssd1 vssd1 vccd1 vccd1 dest_val[19]
+ sky130_fd_sc_hd__a22o_4
XFILLER_0_4_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11579_ _11578_/B _11579_/B vssd1 vssd1 vccd1 vccd1 _11580_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_24_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13318_ _13343_/CLK hold58/X vssd1 vssd1 vccd1 vccd1 hold57/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06960__B _07036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13249_ _13384_/CLK _13249_/D vssd1 vssd1 vccd1 vccd1 hold65/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11156__B2 fanout27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11156__A1 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10903__A1 _09152_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10903__B2 _09172_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07810_ _07810_/A _07810_/B vssd1 vssd1 vccd1 vccd1 _07818_/A sky130_fd_sc_hd__xnor2_1
X_08790_ _08779_/A _08779_/B _08777_/X vssd1 vssd1 vccd1 vccd1 _08835_/A sky130_fd_sc_hd__a21o_2
X_07741_ _07741_/A _07741_/B _07741_/C vssd1 vssd1 vccd1 vccd1 _07742_/B sky130_fd_sc_hd__and3_1
XFILLER_0_35_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11459__A2 _11649_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07672_ _07672_/A _07672_/B vssd1 vssd1 vccd1 vccd1 _07675_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_94_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06623_ _06702_/A _12692_/B vssd1 vssd1 vccd1 vccd1 _06623_/Y sky130_fd_sc_hd__nor2_1
X_09411_ _09411_/A _09411_/B vssd1 vssd1 vccd1 vccd1 _09413_/B sky130_fd_sc_hd__xor2_1
XANTENNA__12408__A1 _11876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09342_ _09343_/A curr_PC[1] vssd1 vssd1 vccd1 vccd1 _09344_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_59_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08088__A1 _08739_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13081__A1 _07263_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08088__B2 _08436_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09273_ _09273_/A _09273_/B _09273_/C _09273_/D vssd1 vssd1 vccd1 vccd1 _09274_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_0_7_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07031__B _10422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08224_ _08742_/A _08224_/B vssd1 vssd1 vccd1 vccd1 _08284_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_31_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08155_ fanout75/X _07752_/B _07955_/A _08304_/B vssd1 vssd1 vccd1 vccd1 _08156_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_15_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07106_ _07671_/A _07671_/B vssd1 vssd1 vccd1 vccd1 _07107_/B sky130_fd_sc_hd__and2b_1
XANTENNA__07063__A2 _07089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08086_ fanout99/X _08741_/A2 _08617_/B _12818_/A vssd1 vssd1 vccd1 vccd1 _08087_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_15_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07037_ _10422_/A _07037_/B vssd1 vssd1 vccd1 vccd1 _09400_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_30_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12344__B1 _11624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08988_ _08988_/A _08988_/B vssd1 vssd1 vccd1 vccd1 _09960_/B sky130_fd_sc_hd__nor2_1
XANTENNA__07771__B1 _08739_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07939_ _08060_/A _08060_/B _07935_/Y vssd1 vssd1 vccd1 vccd1 _08072_/A sky130_fd_sc_hd__a21o_1
XANTENNA__07523__B1 _10413_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10950_ _10950_/A _10950_/B _10950_/C vssd1 vssd1 vccd1 vccd1 _11076_/D sky130_fd_sc_hd__and3_1
X_10881_ _11231_/S _09823_/X _10880_/X _11233_/S vssd1 vssd1 vccd1 vccd1 _10881_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09609_ _11294_/A _09609_/B vssd1 vssd1 vccd1 vccd1 _09611_/B sky130_fd_sc_hd__or2_1
X_12620_ _12620_/A _12620_/B vssd1 vssd1 vccd1 vccd1 new_PC[26] sky130_fd_sc_hd__xnor2_4
XANTENNA__09421__B _12316_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10673__A3 fanout48/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10567__B _12316_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12551_ _12551_/A _12551_/B _12551_/C vssd1 vssd1 vccd1 vccd1 _12552_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_81_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07826__A1 fanout69/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07826__B2 _08216_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12482_ _12488_/B _12482_/B vssd1 vssd1 vccd1 vccd1 new_PC[5] sky130_fd_sc_hd__and2_4
XFILLER_0_81_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11502_ _11503_/A _11503_/B vssd1 vssd1 vccd1 vccd1 _11603_/A sky130_fd_sc_hd__and2_1
XFILLER_0_124_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09579__A1 _10445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09579__B2 _10706_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11433_ _09027_/C _11431_/X _11432_/X vssd1 vssd1 vccd1 vccd1 _11433_/Y sky130_fd_sc_hd__a21boi_1
XANTENNA__09149__A _12626_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11386__B2 _09396_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11386__A1 _09609_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11364_ _12261_/A _11364_/B vssd1 vssd1 vccd1 vccd1 _11371_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__13127__A2 _12789_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13103_ hold240/X _13102_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13103_/X sky130_fd_sc_hd__mux2_1
XANTENNA__11138__A1 _11876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11295_ _11295_/A _11295_/B vssd1 vssd1 vccd1 vccd1 _11297_/B sky130_fd_sc_hd__xnor2_1
X_10315_ _10471_/B _10315_/B vssd1 vssd1 vccd1 vccd1 _10342_/A sky130_fd_sc_hd__or2_1
XFILLER_0_21_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10246_ _10252_/S _10245_/X _09181_/X vssd1 vssd1 vccd1 vccd1 _10246_/X sky130_fd_sc_hd__o21a_1
X_13034_ hold80/A _06572_/A rst vssd1 vssd1 vccd1 vccd1 _13034_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__07892__A _08724_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_4_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10897__A0 _09527_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10177_ _10292_/B _10176_/B _10159_/Y vssd1 vssd1 vccd1 vccd1 _10178_/C sky130_fd_sc_hd__o21ba_1
XFILLER_0_44_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12818_ _12818_/A _12818_/B vssd1 vssd1 vccd1 vccd1 _12818_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__13063__A1 _07833_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12749_ _12749_/A _12749_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[24] sky130_fd_sc_hd__xnor2_4
XFILLER_0_121_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12692__B _12692_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06690__B _06691_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10493__A _10493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09960_ _10748_/A _09960_/B vssd1 vssd1 vccd1 vccd1 _09961_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_40_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08911_ _08912_/A _08912_/B vssd1 vssd1 vccd1 vccd1 _09058_/A sky130_fd_sc_hd__xor2_1
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09891_ _09890_/B _09891_/B vssd1 vssd1 vccd1 vccd1 _09892_/B sky130_fd_sc_hd__and2b_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12213__A _12213_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08842_ _08034_/A _08034_/B _08034_/C vssd1 vssd1 vccd1 vccd1 _08845_/B sky130_fd_sc_hd__o21ai_1
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08773_ _08774_/A _08774_/B vssd1 vssd1 vccd1 vccd1 _08773_/Y sky130_fd_sc_hd__nand2_1
XANTENNA_fanout184_A _08671_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07724_ _07727_/A _07727_/B vssd1 vssd1 vccd1 vccd1 _07724_/X sky130_fd_sc_hd__or2_1
XFILLER_0_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07655_ _07703_/A vssd1 vssd1 vccd1 vccd1 _07655_/Y sky130_fd_sc_hd__inv_2
XANTENNA__06865__B _09351_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06606_ _06606_/A _06606_/B vssd1 vssd1 vccd1 vccd1 _06846_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_79_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10668__A _10959_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07586_ _07567_/A _07567_/B _07565_/Y vssd1 vssd1 vccd1 vccd1 _07589_/A sky130_fd_sc_hd__a21oi_4
XFILLER_0_48_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12801__A1 _09598_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09325_ _09317_/X _09324_/X _11231_/S vssd1 vssd1 vccd1 vccd1 _09325_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_118_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09256_ _09256_/A _09256_/B vssd1 vssd1 vccd1 vccd1 _09257_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_106_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08207_ _08207_/A _08207_/B vssd1 vssd1 vccd1 vccd1 _08208_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_105_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09187_ _08673_/A _09186_/X _11343_/B vssd1 vssd1 vccd1 vccd1 _09187_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_50_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09430__B1 _08507_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08233__A1 _10537_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08233__B2 _08432_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08138_ _08138_/A _08138_/B vssd1 vssd1 vccd1 vccd1 _08139_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_113_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08069_ _08069_/A _08069_/B vssd1 vssd1 vccd1 vccd1 _08874_/B sky130_fd_sc_hd__xnor2_2
X_10100_ _10100_/A _10100_/B vssd1 vssd1 vccd1 vccd1 _10100_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_fanout97_A _07075_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11080_ _10967_/A _10967_/C _10967_/B vssd1 vssd1 vccd1 vccd1 _11090_/A sky130_fd_sc_hd__a21bo_1
X_10031_ _12138_/A _10031_/B vssd1 vssd1 vccd1 vccd1 _10032_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__07217__A _10165_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11982_ curr_PC[22] curr_PC[23] _11982_/C vssd1 vssd1 vccd1 vccd1 _12058_/B sky130_fd_sc_hd__and3_1
XANTENNA__06775__B _06960_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10933_ _10935_/B _10935_/C _10935_/A vssd1 vssd1 vccd1 vccd1 _10938_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11843__A2 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10864_ _10864_/A _10864_/B vssd1 vssd1 vccd1 vccd1 _10870_/C sky130_fd_sc_hd__or2_1
XPHY_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12603_ reg1_val[24] curr_PC[24] _12622_/S vssd1 vssd1 vccd1 vccd1 _12604_/B sky130_fd_sc_hd__mux2_2
X_10795_ _10928_/A _10795_/B vssd1 vssd1 vccd1 vccd1 _10800_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_26_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12534_ _12692_/B _12534_/B vssd1 vssd1 vccd1 vccd1 _12535_/B sky130_fd_sc_hd__or2_1
XFILLER_0_93_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08472__A1 _08673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07275__A2 _12810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08472__B2 _08798_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10517__S _11886_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12465_ _12474_/A _12465_/B vssd1 vssd1 vccd1 vccd1 _12467_/C sky130_fd_sc_hd__nand2_1
X_12396_ hold268/A _12396_/B vssd1 vssd1 vccd1 vccd1 _12396_/X sky130_fd_sc_hd__or2_1
XFILLER_0_62_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11416_ _11417_/A _11417_/B _11417_/C vssd1 vssd1 vccd1 vccd1 _11416_/X sky130_fd_sc_hd__a21o_1
X_11347_ _11450_/B _11449_/B hold174/A vssd1 vssd1 vccd1 vccd1 _11347_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_111_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08527__A2 _08661_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11278_ _07819_/B _11989_/A _11923_/A fanout24/X vssd1 vssd1 vccd1 vccd1 _11279_/B
+ sky130_fd_sc_hd__o22a_1
X_13017_ _13214_/A hold196/X vssd1 vssd1 vccd1 vccd1 _13311_/D sky130_fd_sc_hd__and2_1
X_10229_ _10231_/A _10231_/B vssd1 vssd1 vccd1 vccd1 _10229_/X sky130_fd_sc_hd__or2_1
Xhold1 hold1/A vssd1 vssd1 vccd1 vccd1 hold1/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07127__A _09442_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06966__A _11020_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09342__A _09343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11834__A2 _12316_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07440_ _09423_/B2 fanout16/X _07282_/B _12802_/A vssd1 vssd1 vccd1 vccd1 _07441_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_71_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07371_ _07570_/S _07371_/B vssd1 vssd1 vccd1 vccd1 _07378_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_57_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09110_ reg1_val[9] reg1_val[22] _09111_/S vssd1 vssd1 vccd1 vccd1 _09110_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_72_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07797__A _08740_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09041_ _08836_/Y _08867_/X _08868_/X vssd1 vssd1 vccd1 vccd1 _09041_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_115_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07018__A2 fanout30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10022__B2 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10022__A1 _09568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09943_ _09943_/A _09943_/B vssd1 vssd1 vccd1 vccd1 _09945_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__11766__B _12214_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09715__A1 fanout23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09715__B2 _07819_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09874_ _11470_/A _09874_/B vssd1 vssd1 vccd1 vccd1 _09878_/A sky130_fd_sc_hd__xnor2_4
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07037__A _10422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08825_ _08825_/A _08825_/B vssd1 vssd1 vccd1 vccd1 _08826_/B sky130_fd_sc_hd__xor2_2
X_08756_ _08756_/A _08756_/B vssd1 vssd1 vccd1 vccd1 _08759_/A sky130_fd_sc_hd__nor2_1
XTAP_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08687_ _08984_/A _08982_/A _08686_/X _08684_/Y vssd1 vssd1 vccd1 vccd1 _08987_/B
+ sky130_fd_sc_hd__o22a_1
X_07707_ fanout69/X _10413_/A _10567_/A _08216_/B vssd1 vssd1 vccd1 vccd1 _07708_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08151__B1 _08723_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13027__A1 _09593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07638_ _12794_/A fanout30/X _07688_/B _08671_/B2 vssd1 vssd1 vccd1 vccd1 _07639_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_82_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07569_ _07569_/A _07569_/B vssd1 vssd1 vccd1 vccd1 _07571_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_48_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09308_ _09953_/A _09308_/B vssd1 vssd1 vccd1 vccd1 _09542_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout12_A _12854_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10580_ _10578_/X _10580_/B vssd1 vssd1 vccd1 vccd1 _10583_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_90_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09239_ _07154_/A _07154_/B _09440_/B1 vssd1 vssd1 vccd1 vccd1 _09241_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_51_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12250_ hold195/A _12434_/B1 _12304_/B _12401_/B1 vssd1 vssd1 vccd1 vccd1 _12250_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_106_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12181_ _12112_/Y _12114_/X _12115_/X vssd1 vssd1 vccd1 vccd1 _12185_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__08757__A2 _09609_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11201_ _11201_/A _11201_/B vssd1 vssd1 vccd1 vccd1 _11203_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__10013__A1 _10948_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10013__B2 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11132_ _06981_/A _12404_/A _11131_/Y vssd1 vssd1 vccd1 vccd1 _11132_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__10564__A2 _10797_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11063_ _11294_/A fanout9/X fanout4/X _11146_/A vssd1 vssd1 vccd1 vccd1 _11064_/B
+ sky130_fd_sc_hd__o22a_1
X_10014_ _11163_/A _10014_/B vssd1 vssd1 vccd1 vccd1 _10016_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__12788__A _12788_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08390__B1 _08038_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12069__A2 _12214_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11965_ _10398_/Y _11964_/Y _12244_/S vssd1 vssd1 vccd1 vccd1 _11965_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_98_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10916_ _10916_/A _10916_/B vssd1 vssd1 vccd1 vccd1 _10967_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__06705__A_N _11343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11896_ _07135_/B _11343_/B _11895_/X _06662_/B vssd1 vssd1 vccd1 vccd1 _11896_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_39_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10847_ _10725_/A _10725_/B _10723_/X vssd1 vssd1 vccd1 vccd1 _10848_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_109_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09101__S _09108_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10778_ curr_PC[9] curr_PC[10] _10779_/D curr_PC[11] vssd1 vssd1 vccd1 vccd1 _10778_/X
+ sky130_fd_sc_hd__a31o_1
X_12517_ _12523_/B _12517_/B vssd1 vssd1 vccd1 vccd1 new_PC[10] sky130_fd_sc_hd__and2_4
XFILLER_0_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12448_ _09343_/A curr_PC[1] _12448_/S vssd1 vssd1 vccd1 vccd1 _12450_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_54_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10004__A1 _07035_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12379_ _12380_/B _12413_/A _12377_/Y _12378_/X vssd1 vssd1 vccd1 vccd1 _12379_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_2_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10555__A2 fanout23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06940_ reg1_val[31] _12341_/A vssd1 vssd1 vccd1 vccd1 _06940_/X sky130_fd_sc_hd__and2_1
XFILLER_0_5_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06871_ _08680_/A _06865_/Y _10378_/A _09527_/A _09350_/A vssd1 vssd1 vccd1 vccd1
+ _06872_/B sky130_fd_sc_hd__o2111a_1
XFILLER_0_66_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08610_ _08697_/A _08697_/B vssd1 vssd1 vccd1 vccd1 _08699_/A sky130_fd_sc_hd__or2_1
XFILLER_0_66_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09590_ _09238_/B _12854_/A fanout7/X _07167_/Y vssd1 vssd1 vccd1 vccd1 _09591_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_89_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08541_ _08570_/B _08570_/A vssd1 vssd1 vccd1 vccd1 _08543_/C sky130_fd_sc_hd__nand2b_1
XANTENNA__11268__B1 fanout12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08472_ _08673_/A fanout87/X fanout82/X _08798_/B2 vssd1 vssd1 vccd1 vccd1 _08473_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_92_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07423_ _12846_/A _09238_/B _09440_/B1 _12848_/A vssd1 vssd1 vccd1 vccd1 _07424_/B
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_9_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07023__C _09147_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout147_A _12804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07239__A2 _09236_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07354_ _07485_/A _07354_/B vssd1 vssd1 vccd1 vccd1 _07355_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_17_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07320__A _09716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07285_ _07149_/A fanout59/X _08436_/B _12214_/A vssd1 vssd1 vccd1 vccd1 _07286_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_33_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09024_ _08426_/A _08426_/B _08708_/X vssd1 vssd1 vccd1 vccd1 _09024_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_31_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10794__A2 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold220 hold220/A vssd1 vssd1 vccd1 vccd1 hold220/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08739__A2 fanout87/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold253 hold253/A vssd1 vssd1 vccd1 vccd1 hold253/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold231 hold231/A vssd1 vssd1 vccd1 vccd1 hold231/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold242 hold242/A vssd1 vssd1 vccd1 vccd1 hold242/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold275 hold275/A vssd1 vssd1 vccd1 vccd1 hold275/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold264 hold264/A vssd1 vssd1 vccd1 vccd1 hold264/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold286 hold286/A vssd1 vssd1 vccd1 vccd1 hold286/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold297 hold297/A vssd1 vssd1 vccd1 vccd1 hold297/X sky130_fd_sc_hd__dlygate4sd3_1
X_09926_ _09927_/A _09927_/B vssd1 vssd1 vccd1 vccd1 _09928_/A sky130_fd_sc_hd__nor2_1
X_09857_ _09765_/A _09765_/B _09763_/X vssd1 vssd1 vccd1 vccd1 _09871_/A sky130_fd_sc_hd__a21oi_4
XANTENNA__07175__B2 _10445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07175__A1 _11294_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09788_ _09789_/A _09789_/B vssd1 vssd1 vccd1 vccd1 _09788_/Y sky130_fd_sc_hd__nor2_1
X_08808_ _08808_/A _08808_/B vssd1 vssd1 vccd1 vccd1 _08813_/A sky130_fd_sc_hd__nor2_1
XANTENNA__06728__A_N _07074_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08739_ _08739_/A1 fanout87/X fanout82/X _08436_/A vssd1 vssd1 vccd1 vccd1 _08740_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11750_ _11750_/A _11750_/B vssd1 vssd1 vccd1 vccd1 _11754_/A sky130_fd_sc_hd__xor2_1
XANTENNA__08124__B1 _11472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10701_ _10701_/A _10701_/B vssd1 vssd1 vccd1 vccd1 _10702_/C sky130_fd_sc_hd__xnor2_1
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11681_ _11682_/A _11682_/B _11682_/C vssd1 vssd1 vccd1 vccd1 _11772_/A sky130_fd_sc_hd__a21oi_1
X_10632_ reg1_val[10] curr_PC[10] vssd1 vssd1 vccd1 vccd1 _10632_/X sky130_fd_sc_hd__and2_1
XANTENNA__07065__B1_N _06963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10575__B _10575_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_693 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13351_ _13357_/CLK _13351_/D vssd1 vssd1 vccd1 vccd1 hold291/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10563_ _10452_/A _10451_/B _10449_/X vssd1 vssd1 vccd1 vccd1 _10566_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_11_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12302_ _11341_/B _12352_/B hold266/A vssd1 vssd1 vccd1 vccd1 _12302_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__06989__A1 _12822_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06989__B2 _12824_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13282_ _13378_/CLK _13282_/D vssd1 vssd1 vccd1 vccd1 hold86/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07650__A2 _12214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10494_ _10229_/X _10861_/C _10861_/D vssd1 vssd1 vccd1 vccd1 _10494_/X sky130_fd_sc_hd__a21bo_1
X_12233_ _12341_/A _12233_/B vssd1 vssd1 vccd1 vccd1 _12233_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__10537__A2 _09568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12164_ _12164_/A vssd1 vssd1 vccd1 vccd1 _12164_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_31_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11115_ _11115_/A _11115_/B vssd1 vssd1 vccd1 vccd1 _11117_/A sky130_fd_sc_hd__nand2_1
X_12095_ _11944_/A _12017_/X _12019_/B vssd1 vssd1 vccd1 vccd1 _12095_/X sky130_fd_sc_hd__o21a_1
X_11046_ _11046_/A _11046_/B vssd1 vssd1 vccd1 vccd1 _11048_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_127_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07405__A _10707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12997_ _13013_/A hold201/X vssd1 vssd1 vccd1 vccd1 hold202/A sky130_fd_sc_hd__and2_1
XFILLER_0_98_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11948_ _11613_/B _11787_/B _11946_/Y _11947_/X vssd1 vssd1 vccd1 vccd1 _11949_/B
+ sky130_fd_sc_hd__o31a_1
X_11879_ _11877_/X _11878_/X _12341_/A vssd1 vssd1 vccd1 vccd1 _11880_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_86_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06963__B _07100_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07140__A _07169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07070_ _07071_/B _07071_/C _07071_/D _11163_/A vssd1 vssd1 vccd1 vccd1 _11271_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_14_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09711_ _09639_/A _09639_/B _09640_/Y vssd1 vssd1 vccd1 vccd1 _09805_/A sky130_fd_sc_hd__o21ai_4
X_07972_ _07972_/A _07972_/B vssd1 vssd1 vccd1 vccd1 _07973_/C sky130_fd_sc_hd__and2_1
X_06923_ instruction[6] instruction[5] _09165_/A vssd1 vssd1 vccd1 vccd1 _06923_/Y
+ sky130_fd_sc_hd__nor3_2
XFILLER_0_93_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06854_ _06648_/D _06836_/B _06843_/X vssd1 vssd1 vccd1 vccd1 _06854_/X sky130_fd_sc_hd__a21o_1
X_09642_ _09643_/A _09643_/B vssd1 vssd1 vccd1 vccd1 _09642_/X sky130_fd_sc_hd__and2_1
XFILLER_0_93_86 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06785_ reg2_val[3] _06799_/B vssd1 vssd1 vccd1 vccd1 _06785_/X sky130_fd_sc_hd__and2_2
X_09573_ _09573_/A _09573_/B _09573_/C vssd1 vssd1 vccd1 vccd1 _09575_/A sky130_fd_sc_hd__and3_1
XANTENNA__07315__A _11987_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout264_A _12455_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08524_ _08730_/A1 _08739_/A1 _08038_/A _08721_/B1 vssd1 vssd1 vccd1 vccd1 _08525_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08455_ _08710_/A _08710_/B vssd1 vssd1 vccd1 vccd1 _08711_/A sky130_fd_sc_hd__or2_1
XFILLER_0_92_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07406_ _12822_/A _10941_/A _08216_/B _12824_/A vssd1 vssd1 vccd1 vccd1 _07407_/B
+ sky130_fd_sc_hd__o22a_1
X_08386_ _08422_/A _08422_/B vssd1 vssd1 vccd1 vccd1 _08386_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_46_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07337_ _07337_/A _07337_/B vssd1 vssd1 vccd1 vccd1 _07338_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_73_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07268_ _07268_/A _07268_/B vssd1 vssd1 vccd1 vccd1 _07269_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_5_360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07199_ reg1_val[9] _07199_/B vssd1 vssd1 vccd1 vccd1 _07199_/Y sky130_fd_sc_hd__xnor2_1
X_09007_ _10625_/B _10625_/C _10748_/C vssd1 vssd1 vccd1 vccd1 _09007_/X sky130_fd_sc_hd__and3_1
XFILLER_0_14_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09909_ _09910_/A _09910_/B vssd1 vssd1 vccd1 vccd1 _09911_/A sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_4_9_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12920_ _13101_/B _13102_/A _12911_/X vssd1 vssd1 vccd1 vccd1 _13106_/B sky130_fd_sc_hd__a21o_1
XANTENNA__10152__B1 _11171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12851_ _12264_/A _13087_/B2 hold141/X _13128_/A vssd1 vssd1 vccd1 vccd1 _13279_/D
+ sky130_fd_sc_hd__o211a_1
X_11802_ _11802_/A _11802_/B vssd1 vssd1 vccd1 vccd1 _11803_/B sky130_fd_sc_hd__xnor2_1
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12782_ _12782_/A _12782_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[31] sky130_fd_sc_hd__xnor2_4
XFILLER_0_95_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06659__B1 _06771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11733_ _11705_/X _11707_/Y _11709_/X _09163_/X _11732_/X vssd1 vssd1 vccd1 vccd1
+ _11733_/X sky130_fd_sc_hd__o221a_1
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11664_ _11664_/A _11664_/B vssd1 vssd1 vccd1 vccd1 _11677_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_52_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10615_ _10615_/A _10615_/B vssd1 vssd1 vccd1 vccd1 _11102_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__10207__A1 _07087_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10207__B2 fanout66/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11595_ _11596_/B _11596_/A vssd1 vssd1 vccd1 vccd1 _11693_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_24_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13334_ _13340_/CLK _13334_/D vssd1 vssd1 vccd1 vccd1 hold99/A sky130_fd_sc_hd__dfxtp_1
X_10546_ _10546_/A _10546_/B vssd1 vssd1 vccd1 vccd1 _10549_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_24_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13265_ _13383_/CLK hold24/X vssd1 vssd1 vccd1 vccd1 hold23/A sky130_fd_sc_hd__dfxtp_1
X_10477_ _10346_/A _10346_/B _10345_/A vssd1 vssd1 vccd1 vccd1 _10487_/A sky130_fd_sc_hd__a21o_1
X_12216_ _12217_/B vssd1 vssd1 vccd1 vccd1 _12216_/Y sky130_fd_sc_hd__inv_2
X_13196_ _13214_/A hold247/X vssd1 vssd1 vccd1 vccd1 _13369_/D sky130_fd_sc_hd__and2_1
XFILLER_0_20_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12147_ _12148_/A _12148_/B vssd1 vssd1 vccd1 vccd1 _12147_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_20_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10772__A1_N _06963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09615__A _11987_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12078_ _12078_/A _12078_/B vssd1 vssd1 vccd1 vccd1 _12079_/B sky130_fd_sc_hd__nor2_1
X_11029_ curr_PC[13] _11139_/C vssd1 vssd1 vccd1 vccd1 _11029_/X sky130_fd_sc_hd__or2_1
XANTENNA__07135__A _07194_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06570_ hold57/X vssd1 vssd1 vccd1 vccd1 _06570_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_86_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10446__A1 _07154_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10997__A2 _10996_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08240_ _08240_/A _08240_/B vssd1 vssd1 vccd1 vccd1 _08244_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_28_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12199__A1 _06924_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_48 reg1_val[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_26 reg2_val[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_37 _10270_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_15 reg1_val[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08171_ _11385_/A _08171_/B vssd1 vssd1 vccd1 vccd1 _08178_/B sky130_fd_sc_hd__xnor2_1
XANTENNA_59 reg2_val[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07122_ _09343_/A _07123_/B vssd1 vssd1 vccd1 vccd1 _09593_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_7_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07053_ _09423_/B2 fanout23/X _12802_/A _11171_/A vssd1 vssd1 vccd1 vccd1 _07054_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_30_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_439 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11174__A2 _07087_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07955_ _07955_/A _09396_/B vssd1 vssd1 vccd1 vccd1 _07956_/C sky130_fd_sc_hd__or2_1
XFILLER_0_128_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06906_ instruction[12] _06884_/Y _06905_/X _06694_/B vssd1 vssd1 vccd1 vccd1 reg1_idx[1]
+ sky130_fd_sc_hd__o211a_4
XANTENNA__06889__B1 _09170_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09625_ _09626_/A _09626_/B vssd1 vssd1 vccd1 vccd1 _09625_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_37_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07886_ _11385_/A _07886_/B _07886_/C vssd1 vssd1 vccd1 vccd1 _07889_/B sky130_fd_sc_hd__nand3_1
X_06837_ reg1_val[30] _07345_/A vssd1 vssd1 vccd1 vccd1 _06837_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__07550__B2 _12794_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07550__A1 _08671_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06768_ reg1_val[6] _07036_/A vssd1 vssd1 vccd1 vccd1 _06769_/B sky130_fd_sc_hd__and2_1
X_09556_ _09556_/A _09556_/B vssd1 vssd1 vccd1 vccd1 _09558_/C sky130_fd_sc_hd__xnor2_1
X_06699_ reg1_val[17] _07130_/A vssd1 vssd1 vccd1 vccd1 _06700_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_93_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08507_ _08673_/A _08507_/B vssd1 vssd1 vccd1 vccd1 _08546_/A sky130_fd_sc_hd__or2_1
X_09487_ _09706_/A _09487_/B _09487_/C _09953_/A vssd1 vssd1 vccd1 vccd1 _09487_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_92_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08438_ _08439_/B _08439_/C _08731_/A vssd1 vssd1 vccd1 vccd1 _08442_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_19_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08369_ _08387_/A _08366_/Y _08368_/A vssd1 vssd1 vccd1 vccd1 _08376_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_34_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10400_ _12254_/A1 _10387_/Y _10388_/X _06924_/X _10399_/X vssd1 vssd1 vccd1 vccd1
+ _10400_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_73_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07605__A2 fanout94/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08802__B2 _07752_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08802__A1 _07821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11380_ _12073_/A _11380_/B vssd1 vssd1 vccd1 vccd1 _11381_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_103_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10331_ _11065_/A _07688_/B _10963_/A fanout29/X vssd1 vssd1 vccd1 vccd1 _10332_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_21_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10262_ _10254_/Y _10255_/X _10261_/X vssd1 vssd1 vccd1 vccd1 _10262_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_104_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13050_ hold164/A _12788_/A _13236_/B hold152/X _13113_/A vssd1 vssd1 vccd1 vccd1
+ hold153/A sky130_fd_sc_hd__o221a_1
XANTENNA__11165__A2 fanout12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12001_ _12002_/A _12002_/B vssd1 vssd1 vccd1 vccd1 _12081_/A sky130_fd_sc_hd__and2_1
X_10193_ _10193_/A _10193_/B vssd1 vssd1 vccd1 vccd1 _10194_/B sky130_fd_sc_hd__or2_1
XFILLER_0_108_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06778__B _06799_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08318__B1 _08617_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12903_ hold90/X hold258/X vssd1 vssd1 vccd1 vccd1 _12903_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_17_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12834_ _12834_/A _12848_/B vssd1 vssd1 vccd1 vccd1 _12834_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__09818__B1 _11624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09170__A _09170_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12765_ _12782_/A _12765_/B vssd1 vssd1 vccd1 vccd1 _12768_/B sky130_fd_sc_hd__nand2_1
X_11716_ _11716_/A _11716_/B vssd1 vssd1 vccd1 vccd1 _11718_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_84_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12696_ _12701_/B _12696_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[13] sky130_fd_sc_hd__and2_4
X_11647_ curr_PC[19] _11734_/C _12448_/S vssd1 vssd1 vccd1 vccd1 _11647_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_4_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11578_ _11579_/B _11578_/B vssd1 vssd1 vccd1 vccd1 _11580_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13317_ _13343_/CLK hold106/X vssd1 vssd1 vccd1 vccd1 hold296/A sky130_fd_sc_hd__dfxtp_1
X_10529_ _12254_/A1 _10516_/Y _10528_/Y _10113_/A _10527_/X vssd1 vssd1 vccd1 vccd1
+ _10529_/X sky130_fd_sc_hd__o221a_1
XANTENNA__06960__C _06960_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13248_ hold160/X _12789_/C _13242_/A vssd1 vssd1 vccd1 vccd1 hold161/A sky130_fd_sc_hd__o21a_1
XFILLER_0_58_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11156__A2 _11751_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13179_ _12878_/X _13179_/B vssd1 vssd1 vccd1 vccd1 _13180_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_110_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07740_ _07741_/B _07741_/C _07741_/A vssd1 vssd1 vccd1 vccd1 _08013_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__08309__B1 _08038_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11459__A3 _11649_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07671_ _07671_/A _07671_/B vssd1 vssd1 vccd1 vccd1 _07675_/A sky130_fd_sc_hd__xor2_1
X_06622_ instruction[38] _06634_/B vssd1 vssd1 vccd1 vccd1 _12692_/B sky130_fd_sc_hd__and2_4
XFILLER_0_90_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09410_ _09411_/A _09411_/B vssd1 vssd1 vccd1 vccd1 _09633_/A sky130_fd_sc_hd__nand2_1
X_09341_ _09341_/A vssd1 vssd1 vccd1 vccd1 _09341_/Y sky130_fd_sc_hd__inv_2
XANTENNA__08088__A2 _08744_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13081__A2 _13087_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12813__C1 _13128_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09272_ _09273_/A _09273_/B _09273_/C _09273_/D vssd1 vssd1 vccd1 vccd1 _09272_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_35_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07031__C _07037_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08223_ _08739_/A1 _08741_/A2 _08617_/B _08436_/A vssd1 vssd1 vccd1 vccd1 _08224_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_16_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08154_ _08740_/A _08154_/B vssd1 vssd1 vccd1 vccd1 _08158_/A sky130_fd_sc_hd__xnor2_2
X_08085_ _08912_/A _08912_/B _08910_/A vssd1 vssd1 vccd1 vccd1 _08085_/X sky130_fd_sc_hd__a21bo_1
X_07105_ _07093_/A _07093_/B _07637_/A vssd1 vssd1 vccd1 vccd1 _07671_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_31_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08796__B1 _08216_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07036_ _07036_/A _07036_/B vssd1 vssd1 vccd1 vccd1 _07036_/X sky130_fd_sc_hd__xor2_4
XFILLER_0_30_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08987_ _08987_/A _08987_/B vssd1 vssd1 vccd1 vccd1 _08988_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07771__B2 _08216_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07771__A1 fanout69/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07938_ _07938_/A _07938_/B vssd1 vssd1 vccd1 vccd1 _08060_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_97_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07523__A1 _10574_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07869_ _08733_/A _07869_/B vssd1 vssd1 vccd1 vccd1 _07876_/A sky130_fd_sc_hd__xnor2_1
X_10880_ _11118_/A _10880_/B vssd1 vssd1 vccd1 vccd1 _10880_/X sky130_fd_sc_hd__or2_1
X_09608_ _09389_/A _09389_/B _09386_/A vssd1 vssd1 vccd1 vccd1 _09626_/A sky130_fd_sc_hd__o21a_1
XANTENNA__07523__B2 _10575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout42_A _12834_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09539_ curr_PC[0] curr_PC[1] curr_PC[2] vssd1 vssd1 vccd1 vccd1 _09701_/B sky130_fd_sc_hd__and3_1
XFILLER_0_66_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12550_ _12551_/A _12551_/B _12551_/C vssd1 vssd1 vccd1 vccd1 _12556_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_65_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07826__A2 _07885_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12481_ _12481_/A _12481_/B _12481_/C vssd1 vssd1 vccd1 vccd1 _12482_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_81_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11501_ _11501_/A _11501_/B vssd1 vssd1 vccd1 vccd1 _11503_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10830__A1 _10707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09579__A2 _11847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11432_ _09027_/C _11431_/X _11876_/A vssd1 vssd1 vccd1 vccd1 _11432_/X sky130_fd_sc_hd__o21a_1
XANTENNA__11386__A2 fanout12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13102_ _13102_/A _13102_/B vssd1 vssd1 vccd1 vccd1 _13102_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_104_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11363_ _11558_/A fanout9/X fanout4/X _11472_/A vssd1 vssd1 vccd1 vccd1 _11364_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06801__A3 _12634_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10314_ _10314_/A _10314_/B vssd1 vssd1 vccd1 vccd1 _10315_/B sky130_fd_sc_hd__nor2_1
X_11294_ _11294_/A _12214_/B vssd1 vssd1 vccd1 vccd1 _11295_/B sky130_fd_sc_hd__or2_1
XFILLER_0_21_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10245_ _11010_/S _09145_/X _09179_/B vssd1 vssd1 vccd1 vccd1 _10245_/X sky130_fd_sc_hd__o21a_1
X_13033_ _07164_/B _12798_/B hold81/X vssd1 vssd1 vccd1 vccd1 _13319_/D sky130_fd_sc_hd__a21oi_1
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10897__A1 _09354_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07211__B1 _08507_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10176_ _10292_/B _10176_/B _10159_/Y vssd1 vssd1 vccd1 vccd1 _10178_/B sky130_fd_sc_hd__nor3b_1
Xfanout190 _09127_/S vssd1 vssd1 vccd1 vccd1 _10113_/A sky130_fd_sc_hd__buf_4
XANTENNA__10649__A1 _07100_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12817_ hold37/X _12818_/B _12816_/Y _13245_/A vssd1 vssd1 vccd1 vccd1 hold38/A sky130_fd_sc_hd__o211a_1
XANTENNA__09104__S _09108_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13063__A2 _13087_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12748_ _12749_/A _12749_/B vssd1 vssd1 vccd1 vccd1 _12754_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_127_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12679_ reg1_val[11] _12680_/B vssd1 vssd1 vccd1 vccd1 _12681_/A sky130_fd_sc_hd__or2_1
XFILLER_0_44_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10493__B _10493_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08910_ _08910_/A _08910_/B vssd1 vssd1 vccd1 vccd1 _09056_/B sky130_fd_sc_hd__and2_1
X_09890_ _09891_/B _09890_/B vssd1 vssd1 vccd1 vccd1 _10076_/B sky130_fd_sc_hd__and2b_1
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08841_ _09033_/A _08839_/X _08840_/Y _09043_/B vssd1 vssd1 vccd1 vccd1 _09040_/A
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_0_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12213__B _12214_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08772_ _08774_/A _08774_/B vssd1 vssd1 vccd1 vccd1 _08772_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__10014__A _11163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07723_ _08745_/A _07723_/B vssd1 vssd1 vccd1 vccd1 _07727_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__10949__A _10949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout177_A _09444_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07654_ _08728_/A _07654_/B vssd1 vssd1 vccd1 vccd1 _07703_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06605_ _06606_/B vssd1 vssd1 vccd1 vccd1 _06605_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_67_409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07585_ _07581_/A _07581_/B _07580_/A vssd1 vssd1 vccd1 vccd1 _07590_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_118_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09324_ _09320_/X _09323_/X _09503_/S vssd1 vssd1 vccd1 vccd1 _09324_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_75_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09255_ _09256_/B _09256_/A vssd1 vssd1 vccd1 vccd1 _09255_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_47_188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08206_ _08207_/A _08207_/B vssd1 vssd1 vccd1 vccd1 _08206_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_121_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09186_ instruction[5] _06853_/X _09168_/A _09185_/Y vssd1 vssd1 vccd1 vccd1 _09186_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_43_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08154__A _08740_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09430__A1 _12840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09430__B2 _12842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08233__A2 _07752_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08137_ _11564_/A _08137_/B vssd1 vssd1 vccd1 vccd1 _08138_/B sky130_fd_sc_hd__xnor2_2
X_08068_ _08848_/A _08848_/B _08061_/X vssd1 vssd1 vccd1 vccd1 _08874_/A sky130_fd_sc_hd__a21o_1
XANTENNA__11719__S _12244_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07019_ _11673_/A _07019_/B vssd1 vssd1 vccd1 vccd1 _07041_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__12404__A _12404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09194__B1 _07282_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10030_ _10413_/A fanout16/X _07282_/B _10567_/A vssd1 vssd1 vccd1 vccd1 _10031_/B
+ sky130_fd_sc_hd__o22a_1
X_11981_ curr_PC[21] curr_PC[22] _11819_/B curr_PC[23] vssd1 vssd1 vccd1 vccd1 _11981_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__11828__B1 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10932_ _10931_/B _10931_/C _12073_/A vssd1 vssd1 vccd1 vccd1 _10935_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_86_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13045__A2 _12830_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10863_ _09810_/A _09810_/B _10368_/X _10864_/B vssd1 vssd1 vccd1 vccd1 _10870_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_38_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12602_ _12605_/D _12602_/B vssd1 vssd1 vccd1 vccd1 new_PC[23] sky130_fd_sc_hd__xnor2_4
XFILLER_0_94_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10794_ _11146_/A fanout15/X _07282_/B _11294_/A vssd1 vssd1 vccd1 vccd1 _10795_/B
+ sky130_fd_sc_hd__o22a_1
XPHY_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12533_ _12692_/B _12534_/B vssd1 vssd1 vccd1 vccd1 _12544_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_54_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08472__A2 fanout87/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12464_ _12639_/B _12464_/B vssd1 vssd1 vccd1 vccd1 _12465_/B sky130_fd_sc_hd__or2_1
XFILLER_0_81_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12395_ _12394_/A _12393_/X _12394_/Y _06923_/Y vssd1 vssd1 vccd1 vccd1 _12395_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_34_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11415_ _11417_/A _11417_/B _11417_/C vssd1 vssd1 vccd1 vccd1 _11511_/A sky130_fd_sc_hd__a21oi_2
X_11346_ hold183/A _11346_/B vssd1 vssd1 vccd1 vccd1 _11449_/B sky130_fd_sc_hd__or2_1
XFILLER_0_111_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13016_ hold195/X _13016_/A2 _13016_/B1 hold169/X vssd1 vssd1 vccd1 vccd1 hold196/A
+ sky130_fd_sc_hd__a22o_1
X_11277_ _12317_/A _11277_/B vssd1 vssd1 vccd1 vccd1 _11281_/B sky130_fd_sc_hd__xnor2_1
X_10228_ _10228_/A _10228_/B vssd1 vssd1 vccd1 vccd1 _10231_/B sky130_fd_sc_hd__xnor2_4
Xhold2 hold2/A vssd1 vssd1 vccd1 vccd1 hold2/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10159_ _10159_/A _10159_/B vssd1 vssd1 vccd1 vccd1 _10159_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_55_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06966__B _07074_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13036__A2 _12788_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12244__A0 _09821_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07370_ _07371_/B vssd1 vssd1 vccd1 vccd1 _07370_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_57_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_528 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09040_ _09040_/A _09042_/B vssd1 vssd1 vccd1 vccd1 _11875_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10558__B1 _07688_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10009__A _10448_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07423__B1 _09440_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10022__A2 _10167_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09942_ _09943_/B _09943_/A vssd1 vssd1 vccd1 vccd1 _09942_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_0_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout294_A _06578_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09715__A2 _10664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09873_ _10941_/A _11751_/A _11766_/A fanout94/X vssd1 vssd1 vccd1 vccd1 _09874_/B
+ sky130_fd_sc_hd__o22a_2
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07037__B _07037_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08824_ _08825_/A _08825_/B vssd1 vssd1 vccd1 vccd1 _08824_/Y sky130_fd_sc_hd__nor2_1
X_08755_ _08754_/B _08755_/B vssd1 vssd1 vccd1 vccd1 _08756_/B sky130_fd_sc_hd__and2b_1
X_07706_ _07808_/A _07706_/B vssd1 vssd1 vccd1 vccd1 _07718_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__10679__A _11269_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08686_ _09445_/A _08677_/X _08685_/A vssd1 vssd1 vccd1 vccd1 _08686_/X sky130_fd_sc_hd__o21ba_1
XANTENNA__08151__A1 _10537_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07637_ _07637_/A _07637_/B vssd1 vssd1 vccd1 vccd1 _07666_/A sky130_fd_sc_hd__and2_1
XANTENNA__08151__B2 _08432_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12235__B1 _11624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07568_ _07568_/A _07568_/B vssd1 vssd1 vccd1 vccd1 _07569_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_48_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09307_ _09307_/A _09307_/B vssd1 vssd1 vccd1 vccd1 _09308_/B sky130_fd_sc_hd__and2_1
XFILLER_0_63_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07499_ _07499_/A _07499_/B vssd1 vssd1 vccd1 vccd1 _07500_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_63_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09238_ _10941_/B _09238_/B vssd1 vssd1 vccd1 vccd1 _09241_/B sky130_fd_sc_hd__or2_1
XFILLER_0_35_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09169_ _09170_/A _09170_/B vssd1 vssd1 vccd1 vccd1 _09169_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_90_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12180_ _12180_/A _12180_/B vssd1 vssd1 vccd1 vccd1 _12180_/X sky130_fd_sc_hd__or2_1
XFILLER_0_9_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11200_ _11201_/A _11201_/B vssd1 vssd1 vccd1 vccd1 _11311_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__10013__A2 _10571_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11131_ _12307_/B1 _11130_/X _06719_/B vssd1 vssd1 vccd1 vccd1 _11131_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_8_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07228__A _08584_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11062_ _11196_/B _11062_/B vssd1 vssd1 vccd1 vccd1 _11072_/A sky130_fd_sc_hd__or2_1
X_10013_ _10948_/B2 _10571_/B _10570_/B fanout74/X vssd1 vssd1 vccd1 vccd1 _10014_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07193__A2 _07220_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09443__A _09593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10589__A _10589_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11964_ _11964_/A _11964_/B vssd1 vssd1 vccd1 vccd1 _11964_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__09162__B _09170_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11895_ _11894_/A _09527_/B _11894_/Y _12307_/B1 vssd1 vssd1 vccd1 vccd1 _11895_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_58_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10915_ _10916_/A _10916_/B vssd1 vssd1 vccd1 vccd1 _11081_/B sky130_fd_sc_hd__nand2b_1
X_10846_ _10846_/A _10846_/B vssd1 vssd1 vccd1 vccd1 _10848_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10777_ _11876_/A _10748_/X _10749_/Y _10776_/X _10747_/X vssd1 vssd1 vccd1 vccd1
+ _10777_/X sky130_fd_sc_hd__a311o_1
XFILLER_0_27_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12516_ _12516_/A _12516_/B _12516_/C vssd1 vssd1 vccd1 vccd1 _12517_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_81_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07653__B1 _11923_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12447_ _12453_/A _12447_/B vssd1 vssd1 vccd1 vccd1 new_PC[0] sky130_fd_sc_hd__and2_4
XFILLER_0_35_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10004__A2 _12264_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12378_ _12276_/X _12328_/A _12330_/B vssd1 vssd1 vccd1 vccd1 _12378_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_22_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11329_ _11224_/A _11222_/X _11244_/S vssd1 vssd1 vccd1 vccd1 _11329_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_5_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07138__A _07140_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06870_ _10109_/A _09964_/A _06870_/C _09686_/B vssd1 vssd1 vccd1 vccd1 _06872_/A
+ sky130_fd_sc_hd__and4b_1
XANTENNA__12698__B _12698_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08540_ _08540_/A _08540_/B vssd1 vssd1 vccd1 vccd1 _08570_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_49_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11268__A1 _10570_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11268__B2 _10571_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08471_ _08442_/A _08442_/B _08442_/C vssd1 vssd1 vccd1 vccd1 _08474_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_49_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09499__S _09666_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07422_ _09442_/A _07422_/B vssd1 vssd1 vccd1 vccd1 _07426_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_9_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07353_ _12822_/A fanout94/X _07178_/Y fanout69/X vssd1 vssd1 vccd1 vccd1 _07354_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_9_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07284_ _09441_/A _07284_/B vssd1 vssd1 vccd1 vccd1 _07290_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09023_ _09023_/A _09023_/B vssd1 vssd1 vccd1 vccd1 _11328_/C sky130_fd_sc_hd__xnor2_1
Xhold210 hold210/A vssd1 vssd1 vccd1 vccd1 hold210/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11728__C1 _12307_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold232 hold232/A vssd1 vssd1 vccd1 vccd1 hold232/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold221 hold221/A vssd1 vssd1 vccd1 vccd1 hold221/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold243 hold243/A vssd1 vssd1 vccd1 vccd1 hold243/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08432__A _08673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold276 hold276/A vssd1 vssd1 vccd1 vccd1 hold276/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold254 hold254/A vssd1 vssd1 vccd1 vccd1 hold254/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold287 hold287/A vssd1 vssd1 vccd1 vccd1 hold287/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold265 hold265/A vssd1 vssd1 vccd1 vccd1 hold265/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold298 hold298/A vssd1 vssd1 vccd1 vccd1 hold298/X sky130_fd_sc_hd__dlygate4sd3_1
X_09925_ _10056_/B _09925_/B vssd1 vssd1 vccd1 vccd1 _09927_/B sky130_fd_sc_hd__or2_1
X_09856_ _09800_/A _09800_/B _09801_/Y vssd1 vssd1 vccd1 vccd1 _09946_/A sky130_fd_sc_hd__a21bo_2
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07175__A2 _10706_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08807_ _08058_/B _08807_/B vssd1 vssd1 vccd1 vccd1 _08808_/B sky130_fd_sc_hd__and2b_1
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09787_ _09787_/A _09787_/B vssd1 vssd1 vccd1 vccd1 _09789_/B sky130_fd_sc_hd__xnor2_1
X_06999_ reg1_val[24] reg1_val[25] _07254_/C vssd1 vssd1 vccd1 vccd1 _06999_/X sky130_fd_sc_hd__or3_1
X_08738_ _08738_/A _08738_/B vssd1 vssd1 vccd1 vccd1 _08749_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__10202__A _11269_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08124__A1 _11367_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08669_ _08667_/B _08669_/B vssd1 vssd1 vccd1 vccd1 _08670_/B sky130_fd_sc_hd__and2b_1
XANTENNA__08124__B2 _08730_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12208__B1 fanout4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10700_ _10700_/A _10700_/B vssd1 vssd1 vccd1 vccd1 _10701_/B sky130_fd_sc_hd__xor2_1
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11680_ _11564_/A _11564_/B _11569_/A vssd1 vssd1 vccd1 vccd1 _11682_/C sky130_fd_sc_hd__o21a_1
X_10631_ reg1_val[10] curr_PC[10] vssd1 vssd1 vccd1 vccd1 _10636_/A sky130_fd_sc_hd__or2_1
XFILLER_0_63_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13350_ _13383_/CLK _13350_/D vssd1 vssd1 vccd1 vccd1 hold284/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10562_ _10562_/A _10562_/B vssd1 vssd1 vccd1 vccd1 _10586_/A sky130_fd_sc_hd__or2_2
XFILLER_0_24_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12301_ hold256/A _12301_/B vssd1 vssd1 vccd1 vccd1 _12352_/B sky130_fd_sc_hd__or2_1
X_13281_ _13378_/CLK hold12/X vssd1 vssd1 vccd1 vccd1 hold11/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06989__A2 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12232_ _12205_/Y _12286_/B _12231_/Y vssd1 vssd1 vccd1 vccd1 _12232_/Y sky130_fd_sc_hd__a21oi_1
X_10493_ _10493_/A _10493_/B vssd1 vssd1 vccd1 vccd1 _10739_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_32_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12163_ _12021_/Y _12281_/A _12161_/Y vssd1 vssd1 vccd1 vccd1 _12164_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__10942__B1 fanout94/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11114_ reg1_val[14] curr_PC[14] vssd1 vssd1 vccd1 vccd1 _11115_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_102_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12094_ _12094_/A _12094_/B vssd1 vssd1 vccd1 vccd1 _12226_/A sky130_fd_sc_hd__nand2_2
X_11045_ _11046_/A _11046_/B vssd1 vssd1 vccd1 vccd1 _11150_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_127_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12996_ _13300_/Q _13004_/A2 _13006_/B1 hold200/X vssd1 vssd1 vccd1 vccd1 hold201/A
+ sky130_fd_sc_hd__a22o_1
X_11947_ _11784_/Y _11946_/Y _11945_/Y vssd1 vssd1 vccd1 vccd1 _11947_/X sky130_fd_sc_hd__o21ba_1
XANTENNA__06963__C _07095_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11878_ _11797_/A _11795_/X _06829_/Y vssd1 vssd1 vccd1 vccd1 _11878_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_55_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10829_ _06971_/B fanout6/X _10707_/A vssd1 vssd1 vccd1 vccd1 _10829_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_39_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07140__B _07140_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10630__C1 _09156_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08051__B1 _08617_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07971_ _07903_/A _07903_/C _07913_/A vssd1 vssd1 vccd1 vccd1 _07972_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_10_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06922_ instruction[22] _06884_/Y _06921_/X _06694_/B vssd1 vssd1 vccd1 vccd1 reg2_idx[4]
+ sky130_fd_sc_hd__o211a_4
X_09710_ _09644_/A _09644_/B _09642_/X vssd1 vssd1 vccd1 vccd1 _09808_/A sky130_fd_sc_hd__a21oi_4
XANTENNA__09083__A _12388_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06853_ instruction[6] _06853_/B _06853_/C _06852_/Y vssd1 vssd1 vccd1 vccd1 _06853_/X
+ sky130_fd_sc_hd__or4b_1
X_09641_ _09641_/A _09641_/B vssd1 vssd1 vccd1 vccd1 _09643_/B sky130_fd_sc_hd__xnor2_4
X_06784_ _06782_/Y _06784_/B vssd1 vssd1 vccd1 vccd1 _06870_/C sky130_fd_sc_hd__nand2b_2
XANTENNA__11118__A _11118_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09572_ _10444_/A _09572_/B vssd1 vssd1 vccd1 vccd1 _09573_/C sky130_fd_sc_hd__xnor2_1
X_08523_ _08733_/A _08523_/B vssd1 vssd1 vccd1 vccd1 _08530_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_26_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08454_ _08454_/A _08454_/B vssd1 vssd1 vccd1 vccd1 _08710_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07331__A _09433_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07405_ _10707_/A _07405_/B vssd1 vssd1 vccd1 vccd1 _07409_/A sky130_fd_sc_hd__xnor2_1
X_08385_ _08385_/A _08385_/B vssd1 vssd1 vccd1 vccd1 _08422_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_46_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07336_ _08584_/A _07336_/B vssd1 vssd1 vccd1 vccd1 _07337_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_61_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07617__B1 _10963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07267_ _07267_/A _07267_/B _07267_/C vssd1 vssd1 vccd1 vccd1 _07268_/B sky130_fd_sc_hd__nor3_1
X_09006_ _09006_/A _09006_/B vssd1 vssd1 vccd1 vccd1 _10748_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_33_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07198_ reg1_val[8] _07200_/A _07215_/B vssd1 vssd1 vccd1 vccd1 _07199_/B sky130_fd_sc_hd__a21o_1
XANTENNA__08162__A _08752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10924__B1 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout72_A _09614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09908_ _09908_/A _09908_/B vssd1 vssd1 vccd1 vccd1 _09910_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__12412__A _12412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09839_ _09673_/X _09674_/Y _09676_/Y vssd1 vssd1 vccd1 vccd1 _09843_/A sky130_fd_sc_hd__o21a_1
XANTENNA__07506__A _09351_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10152__A1 _11065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10152__B2 _11146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12850_ hold140/X _12856_/B vssd1 vssd1 vccd1 vccd1 hold141/A sky130_fd_sc_hd__or2_1
X_11801_ _11718_/A _11718_/B _11716_/B vssd1 vssd1 vccd1 vccd1 _11802_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_68_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09721__A _11673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12781_ reg1_val[31] _12781_/B vssd1 vssd1 vccd1 vccd1 _12782_/B sky130_fd_sc_hd__xnor2_2
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11732_ _06924_/X _11719_/X _11731_/X _11713_/X vssd1 vssd1 vccd1 vccd1 _11732_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11663_ _11663_/A _11663_/B vssd1 vssd1 vccd1 vccd1 _11664_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10614_ _10615_/A _10615_/B vssd1 vssd1 vccd1 vccd1 _10614_/X sky130_fd_sc_hd__and2_1
XANTENNA__10207__A2 _11472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13333_ _13340_/CLK hold94/X vssd1 vssd1 vccd1 vccd1 hold92/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11594_ _11594_/A _11594_/B vssd1 vssd1 vccd1 vccd1 _11596_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_106_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10545_ _11163_/A _10545_/B vssd1 vssd1 vccd1 vccd1 _10546_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_121_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13157__B2 _13246_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13264_ _13383_/CLK hold44/X vssd1 vssd1 vccd1 vccd1 hold43/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09168__A _09168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10476_ _10476_/A _10476_/B vssd1 vssd1 vccd1 vccd1 _10489_/A sky130_fd_sc_hd__xnor2_4
X_13195_ hold246/X _13213_/A2 _13194_/X _13213_/B2 vssd1 vssd1 vccd1 vccd1 hold247/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12215_ _12213_/A _12213_/Y _12215_/S vssd1 vssd1 vccd1 vccd1 _12217_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_20_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12146_ _12146_/A _12146_/B vssd1 vssd1 vccd1 vccd1 _12148_/B sky130_fd_sc_hd__and2_1
XFILLER_0_20_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12077_ _12078_/A _12078_/B vssd1 vssd1 vccd1 vccd1 _12145_/B sky130_fd_sc_hd__and2_1
XANTENNA__09107__S _09108_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06958__C _09669_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07416__A _09445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11028_ _11876_/A _10999_/X _11000_/Y _11027_/X _10998_/X vssd1 vssd1 vccd1 vccd1
+ _11028_/X sky130_fd_sc_hd__a311o_1
XFILLER_0_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13093__A0 hold260/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12979_ _13013_/A hold233/X vssd1 vssd1 vccd1 vccd1 _13292_/D sky130_fd_sc_hd__and2_1
XFILLER_0_86_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10446__A2 _07154_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07151__A _07343_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_38 instruction[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_27 reg2_val[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_16 reg1_val[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08170_ _08752_/A fanout69/X _08216_/B _08798_/B2 vssd1 vssd1 vccd1 vccd1 _08171_/B
+ sky130_fd_sc_hd__o22a_1
X_07121_ _12626_/A reg1_val[31] instruction[7] vssd1 vssd1 vccd1 vccd1 _07123_/B sky130_fd_sc_hd__and3_2
XANTENNA_49 reg1_val[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06990__A _11163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07052_ _11987_/A _11987_/B vssd1 vssd1 vccd1 vccd1 _07052_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_0_100_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09806__A _09808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11174__A3 _12150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07954_ _07099_/A _07099_/B _07752_/B vssd1 vssd1 vccd1 vccd1 _07956_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06905_ instruction[19] _06921_/B vssd1 vssd1 vccd1 vccd1 _06905_/X sky130_fd_sc_hd__or2_1
XANTENNA__10134__A1 _12244_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07885_ _08216_/B _07885_/B vssd1 vssd1 vccd1 vccd1 _07886_/C sky130_fd_sc_hd__or2_1
XANTENNA__06889__A1 _06771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06836_ _06874_/A _06836_/B vssd1 vssd1 vccd1 vccd1 _06853_/B sky130_fd_sc_hd__and2b_1
X_09624_ _09624_/A _09624_/B vssd1 vssd1 vccd1 vccd1 _09626_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_97_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07550__A2 fanout9/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13084__B1 _06892_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06767_ reg1_val[6] _07036_/A vssd1 vssd1 vccd1 vccd1 _06767_/X sky130_fd_sc_hd__or2_1
X_09555_ _11673_/A _09555_/B vssd1 vssd1 vccd1 vccd1 _09556_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__10687__A _11180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06698_ _07130_/A reg1_val[17] vssd1 vssd1 vccd1 vccd1 _06698_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_93_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08506_ _08506_/A _08506_/B vssd1 vssd1 vccd1 vccd1 _08519_/A sky130_fd_sc_hd__xor2_1
X_09486_ _07683_/X _09300_/X _09301_/X vssd1 vssd1 vccd1 vccd1 _09486_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_65_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08437_ _07067_/A _07067_/B _08730_/A1 vssd1 vssd1 vccd1 vccd1 _08439_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08368_ _08368_/A _08368_/B vssd1 vssd1 vccd1 vccd1 _08387_/B sky130_fd_sc_hd__and2_1
XFILLER_0_34_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07319_ _12804_/A fanout23/X _11171_/A _09768_/A1 vssd1 vssd1 vccd1 vccd1 _07320_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_61_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08299_ _08300_/A _08300_/B vssd1 vssd1 vccd1 vccd1 _08342_/A sky130_fd_sc_hd__or2_1
XANTENNA__08263__B1 _08038_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08802__A2 _09609_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10330_ _11180_/A _10330_/B vssd1 vssd1 vccd1 vccd1 _10334_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_5_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10261_ _06867_/B _12402_/A0 _10259_/X _10260_/X vssd1 vssd1 vccd1 vccd1 _10261_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_14_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12000_ _12210_/A _12000_/B vssd1 vssd1 vccd1 vccd1 _12002_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__09716__A _09716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10192_ _10192_/A _10192_/B _10192_/C vssd1 vssd1 vccd1 vccd1 _10193_/B sky130_fd_sc_hd__and3_1
XANTENNA__08318__A1 _07885_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07236__A _09441_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08318__B2 _08721_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12902_ hold242/X hold51/X vssd1 vssd1 vccd1 vccd1 _13119_/B sky130_fd_sc_hd__nand2b_1
XTAP_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12833_ hold21/X _12856_/B _12832_/Y _13235_/A vssd1 vssd1 vccd1 vccd1 hold22/A sky130_fd_sc_hd__o211a_1
XTAP_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12764_ _12764_/A _12773_/A vssd1 vssd1 vccd1 vccd1 _12768_/A sky130_fd_sc_hd__or2_1
X_11715_ reg1_val[20] curr_PC[20] vssd1 vssd1 vccd1 vccd1 _11716_/B sky130_fd_sc_hd__nand2_1
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12695_ _12695_/A _12695_/B _12695_/C vssd1 vssd1 vccd1 vccd1 _12696_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_37_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11646_ curr_PC[19] _11734_/C vssd1 vssd1 vccd1 vccd1 _11646_/X sky130_fd_sc_hd__or2_1
XFILLER_0_25_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12317__A _12317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11577_ _12210_/A _11577_/B vssd1 vssd1 vccd1 vccd1 _11578_/B sky130_fd_sc_hd__xnor2_1
X_13316_ _13380_/CLK _13316_/D vssd1 vssd1 vccd1 vccd1 hold111/A sky130_fd_sc_hd__dfxtp_1
X_10528_ _10119_/S _10118_/X _09181_/X vssd1 vssd1 vccd1 vccd1 _10528_/Y sky130_fd_sc_hd__o21ai_2
XANTENNA__06960__D _09147_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13247_ hold53/X hold167/A _13246_/X _13242_/A vssd1 vssd1 vccd1 vccd1 hold54/A sky130_fd_sc_hd__o211a_1
XFILLER_0_12_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10459_ _10459_/A _10459_/B vssd1 vssd1 vccd1 vccd1 _10460_/B sky130_fd_sc_hd__nand2_1
X_13178_ _13235_/A hold264/X vssd1 vssd1 vccd1 vccd1 _13365_/D sky130_fd_sc_hd__and2_1
XFILLER_0_20_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12129_ _09111_/S _10119_/X _12128_/X vssd1 vssd1 vccd1 vccd1 _12129_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_0_74_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08309__B2 _12820_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08309__A1 _08730_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07670_ _08944_/A _08944_/B _07635_/X vssd1 vssd1 vccd1 vccd1 _07678_/B sky130_fd_sc_hd__a21oi_4
X_06621_ _06621_/A _06621_/B vssd1 vssd1 vccd1 vccd1 _06621_/Y sky130_fd_sc_hd__nand2_1
X_09340_ _09325_/X _09339_/X _10119_/S vssd1 vssd1 vccd1 vccd1 _09341_/A sky130_fd_sc_hd__mux2_1
XANTENNA__09080__B _09170_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09271_ _09270_/B _09270_/C _11987_/A vssd1 vssd1 vccd1 vccd1 _09273_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08222_ _08225_/A _08225_/B vssd1 vssd1 vccd1 vccd1 _08222_/X sky130_fd_sc_hd__or2_1
XFILLER_0_7_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout122_A _06971_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08153_ _07885_/B fanout87/X fanout82/X _08721_/B1 vssd1 vssd1 vccd1 vccd1 _08154_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_15_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08084_ _08909_/A _08909_/B vssd1 vssd1 vccd1 vccd1 _08910_/A sky130_fd_sc_hd__or2_1
X_07104_ _07636_/A _07636_/B vssd1 vssd1 vccd1 vccd1 _07637_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_43_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08796__A1 _07955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08796__B2 _07896_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07035_ _07036_/A _07036_/B vssd1 vssd1 vccd1 vccd1 _07035_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_0_3_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08986_ _09656_/B _09656_/C vssd1 vssd1 vccd1 vccd1 _08988_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07771__A2 _08721_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07046__A_N _11172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07937_ _08598_/A _07937_/B vssd1 vssd1 vccd1 vccd1 _08060_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__07523__A2 _12810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07868_ _08732_/A2 _11472_/A _11558_/A _08656_/B vssd1 vssd1 vccd1 vccd1 _07869_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_3_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06819_ _10752_/A _06818_/X _06734_/X vssd1 vssd1 vccd1 vccd1 _06819_/X sky130_fd_sc_hd__o21ba_1
X_09607_ _09607_/A _09607_/B vssd1 vssd1 vccd1 vccd1 _09628_/A sky130_fd_sc_hd__xor2_1
X_07799_ _08304_/B _08436_/A vssd1 vssd1 vccd1 vccd1 _07800_/C sky130_fd_sc_hd__nor2_1
X_09538_ _09491_/X _09493_/X _09533_/X _09537_/X _06881_/X vssd1 vssd1 vccd1 vccd1
+ _09538_/X sky130_fd_sc_hd__a41o_2
XANTENNA_fanout35_A _07504_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09469_ _09469_/A _09469_/B vssd1 vssd1 vccd1 vccd1 _09474_/A sky130_fd_sc_hd__or2_4
X_11500_ _11501_/A _11501_/B vssd1 vssd1 vccd1 vccd1 _11599_/B sky130_fd_sc_hd__and2b_1
XANTENNA_fanout1_A fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12480_ _12481_/A _12481_/B _12481_/C vssd1 vssd1 vccd1 vccd1 _12488_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_80_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11431_ _11328_/B _11328_/C _11792_/A vssd1 vssd1 vccd1 vccd1 _11431_/X sky130_fd_sc_hd__a21o_1
XANTENNA__09984__B1 _06939_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11362_ _11304_/A _11304_/B _11306_/B _11307_/X vssd1 vssd1 vccd1 vccd1 _11414_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_22_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13101_ _12911_/X _13101_/B vssd1 vssd1 vccd1 vccd1 _13102_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__11791__B1 _12290_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10313_ _10314_/A _10314_/B vssd1 vssd1 vccd1 vccd1 _10471_/B sky130_fd_sc_hd__and2_1
XANTENNA__10880__A _11118_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11293_ _11293_/A _11293_/B vssd1 vssd1 vccd1 vccd1 _11295_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_21_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13032_ _06570_/Y _06572_/A _06892_/B hold80/X rst vssd1 vssd1 vccd1 vccd1 hold81/A
+ sky130_fd_sc_hd__a221o_1
X_10244_ _06867_/B _10242_/X _10243_/Y vssd1 vssd1 vccd1 vccd1 _10270_/C sky130_fd_sc_hd__o21a_1
XANTENNA__09736__B1 _11923_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07211__B2 _12832_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07211__A1 _10589_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10175_ _10174_/B _10174_/C _10174_/A vssd1 vssd1 vccd1 vccd1 _10176_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout191 _09111_/S vssd1 vssd1 vccd1 vccd1 _09108_/S sky130_fd_sc_hd__clkbuf_8
Xfanout180 _07043_/Y vssd1 vssd1 vccd1 vccd1 _09423_/B2 sky130_fd_sc_hd__buf_8
XANTENNA__10649__A2 _12404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12816_ _12816_/A _12818_/B vssd1 vssd1 vccd1 vccd1 _12816_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_84_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_112 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08475__B1 _08038_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12747_ _12728_/B _12746_/X _12741_/B _07254_/C vssd1 vssd1 vccd1 vccd1 _12749_/B
+ sky130_fd_sc_hd__a2bb2o_2
XANTENNA__08525__A _08681_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12678_ _12683_/B _12678_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[10] sky130_fd_sc_hd__and2_4
XANTENNA__09120__S _09142_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11629_ _11629_/A _11629_/B vssd1 vssd1 vccd1 vccd1 _11629_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_65_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11886__A _11886_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06699__B _07130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11534__B1 _11886_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08840_ _08838_/A _08838_/B _08786_/Y vssd1 vssd1 vccd1 vccd1 _08840_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_0_20_270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08771_ _08120_/A _08120_/B _08118_/X vssd1 vssd1 vccd1 vccd1 _08774_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_18_60 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07722_ _10927_/A1 _10167_/A1 _10022_/B1 _11367_/A vssd1 vssd1 vccd1 vccd1 _07723_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11837__A1 _07033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07653_ _08727_/B1 _11989_/A _11923_/A _08727_/A2 vssd1 vssd1 vccd1 vccd1 _07654_/B
+ sky130_fd_sc_hd__o22a_1
X_06604_ _07144_/A reg1_val[27] vssd1 vssd1 vccd1 vccd1 _06606_/B sky130_fd_sc_hd__nand2b_2
X_09323_ _09321_/X _09322_/X _09663_/S vssd1 vssd1 vccd1 vccd1 _09323_/X sky130_fd_sc_hd__mux2_1
X_07584_ _07582_/A _07575_/Y _07583_/X vssd1 vssd1 vccd1 vccd1 _07595_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_34_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09254_ _12412_/B _09254_/B vssd1 vssd1 vccd1 vccd1 _09256_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_8_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09185_ _06861_/Y _06939_/B _09082_/X _09184_/X vssd1 vssd1 vccd1 vccd1 _09185_/Y
+ sky130_fd_sc_hd__a211oi_1
XANTENNA__08218__B1 _08656_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08205_ _08207_/A _08207_/B vssd1 vssd1 vccd1 vccd1 _08205_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_28_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08136_ _08752_/A _09609_/B _09396_/B _08798_/B2 vssd1 vssd1 vccd1 vccd1 _08137_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09430__A2 _10589_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08067_ _08067_/A _08067_/B vssd1 vssd1 vccd1 vccd1 _08848_/B sky130_fd_sc_hd__xnor2_4
X_07018_ _08671_/B2 fanout30/X _12798_/A _07688_/B vssd1 vssd1 vccd1 vccd1 _07019_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_101_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09194__B2 _12804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09194__A1 _12802_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08969_ _08971_/A _08971_/B vssd1 vssd1 vccd1 vccd1 _09487_/B sky130_fd_sc_hd__nor2_1
X_11980_ _11707_/A _11950_/Y _11951_/Y _11979_/X vssd1 vssd1 vccd1 vccd1 _11980_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__11828__B2 fanout27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11828__A1 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10931_ _12073_/A _10931_/B _10931_/C vssd1 vssd1 vccd1 vccd1 _10935_/B sky130_fd_sc_hd__nand3_1
XANTENNA__11036__A _12210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10862_ _10862_/A vssd1 vssd1 vccd1 vccd1 _10864_/B sky130_fd_sc_hd__inv_2
XPHY_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12601_ _12593_/B _12598_/B _12591_/X vssd1 vssd1 vccd1 vccd1 _12602_/B sky130_fd_sc_hd__a21o_1
X_10793_ _10793_/A _10793_/B vssd1 vssd1 vccd1 vccd1 _10802_/A sky130_fd_sc_hd__xor2_1
XPHY_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12532_ reg1_val[13] curr_PC[13] _12586_/S vssd1 vssd1 vccd1 vccd1 _12534_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_94_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12463_ _12639_/B _12464_/B vssd1 vssd1 vccd1 vccd1 _12474_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_53_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11414_ _11414_/A _11414_/B vssd1 vssd1 vccd1 vccd1 _11417_/C sky130_fd_sc_hd__xnor2_2
XFILLER_0_111_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12394_ _12394_/A _12394_/B vssd1 vssd1 vccd1 vccd1 _12394_/Y sky130_fd_sc_hd__nand2_1
X_11345_ _09167_/Y _11340_/X _11341_/Y _11344_/X vssd1 vssd1 vccd1 vccd1 _11345_/X
+ sky130_fd_sc_hd__a31o_2
XANTENNA__06786__A3 _12644_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12308__A2 _11973_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11276_ _10574_/B fanout15/X fanout36/X _11751_/A vssd1 vssd1 vccd1 vccd1 _11277_/B
+ sky130_fd_sc_hd__o22a_1
X_13015_ _13214_/A hold224/X vssd1 vssd1 vccd1 vccd1 _13310_/D sky130_fd_sc_hd__and2_1
XFILLER_0_120_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10227_ _10227_/A _10227_/B vssd1 vssd1 vccd1 vccd1 _10228_/B sky130_fd_sc_hd__xor2_4
Xhold3 hold3/A vssd1 vssd1 vccd1 vccd1 hold3/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09904__A _10710_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10158_ _10159_/B vssd1 vssd1 vccd1 vccd1 _10158_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_55_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10089_ _10090_/B _10090_/A vssd1 vssd1 vccd1 vccd1 _10089_/X sky130_fd_sc_hd__and2b_1
XANTENNA__07424__A _09441_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10785__A _11470_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_746 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10558__A1 _11146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10558__B2 _11294_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12505__A _12669_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07423__B2 _12848_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07423__A1 _12846_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08620__A0 _09433_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09941_ _09941_/A _09941_/B vssd1 vssd1 vccd1 vccd1 _09943_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_40_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09872_ _09722_/A _09722_/B _09719_/A vssd1 vssd1 vccd1 vccd1 _09885_/A sky130_fd_sc_hd__o21ai_4
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08823_ _08759_/A _08759_/B _08756_/A vssd1 vssd1 vccd1 vccd1 _08825_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_29_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08754_ _08755_/B _08754_/B vssd1 vssd1 vccd1 vccd1 _08756_/A sky130_fd_sc_hd__and2b_1
X_07705_ _12210_/A _07705_/B vssd1 vssd1 vccd1 vccd1 _07706_/B sky130_fd_sc_hd__xnor2_1
XTAP_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08685_ _08685_/A _08685_/B vssd1 vssd1 vccd1 vccd1 _08982_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__08151__A2 _07896_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07636_ _07636_/A _07636_/B vssd1 vssd1 vccd1 vccd1 _07637_/B sky130_fd_sc_hd__or2_1
X_07567_ _07567_/A _07567_/B vssd1 vssd1 vccd1 vccd1 _07582_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_48_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06892__B _06892_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09306_ _09066_/A _09066_/B _09072_/Y _09649_/B _09706_/A vssd1 vssd1 vccd1 vccd1
+ _09307_/B sky130_fd_sc_hd__a2111o_1
X_07498_ _07499_/A _07499_/B vssd1 vssd1 vccd1 vccd1 _07498_/X sky130_fd_sc_hd__and2_1
X_09237_ _09594_/A _09237_/B vssd1 vssd1 vccd1 vccd1 _09237_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_36_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08165__A _08752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09168_ _09168_/A _09170_/A vssd1 vssd1 vccd1 vccd1 _09168_/X sky130_fd_sc_hd__or2_1
XFILLER_0_121_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09099_ _09091_/X _09098_/X _10248_/S vssd1 vssd1 vccd1 vccd1 _09099_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_31_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08119_ _08119_/A _08119_/B vssd1 vssd1 vccd1 vccd1 _08120_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_16_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11130_ _09527_/B _09354_/B _11130_/S vssd1 vssd1 vccd1 vccd1 _11130_/X sky130_fd_sc_hd__mux2_1
XANTENNA__07509__A _12138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11061_ _11061_/A _11061_/B vssd1 vssd1 vccd1 vccd1 _11062_/B sky130_fd_sc_hd__nor2_1
XANTENNA__11973__B _11973_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12710__A2 _12703_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10012_ _10710_/A _10012_/B vssd1 vssd1 vccd1 vccd1 _10016_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__12150__A _12150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10589__B fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11963_ _11883_/A _11885_/B _11883_/B vssd1 vssd1 vccd1 vccd1 _11964_/B sky130_fd_sc_hd__a21boi_1
XFILLER_0_86_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11894_ _11894_/A _11973_/B vssd1 vssd1 vccd1 vccd1 _11894_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_58_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10914_ _11081_/A _10914_/B vssd1 vssd1 vccd1 vccd1 _10916_/B sky130_fd_sc_hd__and2_1
X_10845_ _10843_/X _10845_/B vssd1 vssd1 vccd1 vccd1 _10846_/B sky130_fd_sc_hd__and2b_1
XANTENNA__10237__B1 _12290_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10776_ _09172_/B _10763_/Y _10775_/Y _10753_/X vssd1 vssd1 vccd1 vccd1 _10776_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_82_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07102__B1 _10567_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12515_ _12516_/A _12516_/B _12516_/C vssd1 vssd1 vccd1 vccd1 _12523_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_82_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07653__A1 _08727_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07653__B2 _08727_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12446_ _12626_/B _12446_/B vssd1 vssd1 vccd1 vccd1 _12447_/B sky130_fd_sc_hd__or2_1
XFILLER_0_35_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08803__A _11564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08602__B1 _09568_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12377_ _12164_/Y _12281_/B _12283_/Y vssd1 vssd1 vccd1 vccd1 _12377_/Y sky130_fd_sc_hd__o21ai_1
X_11328_ _11792_/A _11328_/B _11328_/C vssd1 vssd1 vccd1 vccd1 _11328_/X sky130_fd_sc_hd__or3_1
XFILLER_0_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11259_ _11908_/A _11259_/B vssd1 vssd1 vccd1 vccd1 _11263_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_89_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07154__A _07154_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11268__A2 _12316_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07341__B1 _12844_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08470_ _08483_/A _08483_/B vssd1 vssd1 vccd1 vccd1 _08485_/A sky130_fd_sc_hd__nand2b_1
X_07421_ _08436_/B _12854_/A fanout7/X _07149_/A vssd1 vssd1 vccd1 vccd1 _07422_/B
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_15_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07352_ _10707_/A _07352_/B vssd1 vssd1 vccd1 vccd1 _07356_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07283_ _09238_/B fanout48/X _10570_/B _09440_/B1 vssd1 vssd1 vccd1 vccd1 _07284_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_31_60 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09022_ _11107_/B _11107_/C _11221_/A vssd1 vssd1 vccd1 vccd1 _11328_/B sky130_fd_sc_hd__and3_1
XFILLER_0_31_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold211 hold211/A vssd1 vssd1 vccd1 vccd1 hold211/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold200 hold200/A vssd1 vssd1 vccd1 vccd1 hold200/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_4_3_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13376_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold222 hold222/A vssd1 vssd1 vccd1 vccd1 hold222/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold233 hold233/A vssd1 vssd1 vccd1 vccd1 hold233/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout202_A _12830_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold244 hold244/A vssd1 vssd1 vccd1 vccd1 hold244/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09528__B hold260/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07329__A _10710_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08432__B _08432_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold277 hold277/A vssd1 vssd1 vccd1 vccd1 hold277/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold266 hold266/A vssd1 vssd1 vccd1 vccd1 hold266/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold255 hold255/A vssd1 vssd1 vccd1 vccd1 hold255/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold288 hold288/A vssd1 vssd1 vccd1 vccd1 hold288/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold299 hold299/A vssd1 vssd1 vccd1 vccd1 hold299/X sky130_fd_sc_hd__dlygate4sd3_1
X_09924_ _09923_/A _09923_/B _09923_/C vssd1 vssd1 vccd1 vccd1 _09925_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09855_ _09805_/A _09805_/B _09803_/X vssd1 vssd1 vccd1 vccd1 _09949_/A sky130_fd_sc_hd__a21oi_4
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08806_ _08853_/B _08806_/B vssd1 vssd1 vccd1 vccd1 _08815_/A sky130_fd_sc_hd__or2_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07064__A _12423_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09786_ _09786_/A _09786_/B vssd1 vssd1 vccd1 vccd1 _09787_/B sky130_fd_sc_hd__xor2_2
X_06998_ reg1_val[23] _06998_/B _12726_/B vssd1 vssd1 vccd1 vccd1 _07254_/C sky130_fd_sc_hd__or3_4
X_08737_ _08738_/A _08738_/B vssd1 vssd1 vccd1 vccd1 _08737_/X sky130_fd_sc_hd__and2b_1
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08668_ _08683_/A _08683_/B _08669_/B vssd1 vssd1 vccd1 vccd1 _08668_/X sky130_fd_sc_hd__or3_1
XANTENNA__08124__A2 _08038_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07619_ _10445_/A _11065_/A _11146_/A _10706_/B2 vssd1 vssd1 vccd1 vccd1 _07620_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12208__A1 _12316_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10630_ _10629_/A _10629_/B _10629_/Y _09156_/Y vssd1 vssd1 vccd1 vccd1 _10630_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08599_ _08646_/B2 _08732_/A2 _09440_/B1 _09423_/B2 vssd1 vssd1 vccd1 vccd1 _08600_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_49_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12208__B2 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10561_ _10560_/B _10561_/B vssd1 vssd1 vccd1 vccd1 _10562_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_24_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13280_ _13365_/CLK hold32/X vssd1 vssd1 vccd1 vccd1 hold31/A sky130_fd_sc_hd__dfxtp_1
X_12300_ _12429_/B _12298_/Y _12299_/Y _06924_/X vssd1 vssd1 vccd1 vccd1 _12300_/X
+ sky130_fd_sc_hd__a211o_1
X_10492_ _10493_/A _10493_/B vssd1 vssd1 vccd1 vccd1 _10492_/X sky130_fd_sc_hd__and2b_1
X_12231_ _12205_/Y _12286_/B _11707_/A vssd1 vssd1 vccd1 vccd1 _12231_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_32_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12162_ _12162_/A _12226_/A vssd1 vssd1 vccd1 vccd1 _12281_/A sky130_fd_sc_hd__or2_1
XANTENNA__10942__A1 _07154_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11113_ reg1_val[14] curr_PC[14] vssd1 vssd1 vccd1 vccd1 _11115_/A sky130_fd_sc_hd__or2_1
X_12093_ _12093_/A _12093_/B _12093_/C vssd1 vssd1 vccd1 vccd1 _12094_/B sky130_fd_sc_hd__nand3_1
X_11044_ _06985_/A fanout8/X _11043_/X vssd1 vssd1 vccd1 vccd1 _11046_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_36_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12995_ _13013_/A hold175/X vssd1 vssd1 vccd1 vccd1 hold176/A sky130_fd_sc_hd__and2_1
XFILLER_0_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11946_ _12098_/A _12098_/B vssd1 vssd1 vccd1 vccd1 _11946_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_86_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_48 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11877_ _11797_/A _11794_/X _11811_/S vssd1 vssd1 vccd1 vccd1 _11877_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_74_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06963__D _07089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10828_ _11164_/A _10828_/B vssd1 vssd1 vccd1 vccd1 _10961_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_125_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10759_ _10759_/A _11886_/A _10757_/X vssd1 vssd1 vccd1 vccd1 _10759_/X sky130_fd_sc_hd__or3b_1
XFILLER_0_82_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10782__B _10782_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12429_ reg1_val[30] _12429_/B _12429_/C vssd1 vssd1 vccd1 vccd1 _12430_/B sky130_fd_sc_hd__and3_1
XFILLER_0_23_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07149__A _07149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08051__B2 _08732_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08051__A1 _08741_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07970_ _07969_/A _07969_/B _07969_/C vssd1 vssd1 vccd1 vccd1 _07973_/B sky130_fd_sc_hd__o21ai_1
X_06921_ instruction[29] _06921_/B vssd1 vssd1 vccd1 vccd1 _06921_/X sky130_fd_sc_hd__or2_1
XANTENNA__06988__A _06988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06852_ reg1_val[31] _07420_/A vssd1 vssd1 vccd1 vccd1 _06852_/Y sky130_fd_sc_hd__nand2_1
X_09640_ _09641_/B _09641_/A vssd1 vssd1 vccd1 vccd1 _09640_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_117_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06783_ reg1_val[4] _10252_/S vssd1 vssd1 vccd1 vccd1 _06784_/B sky130_fd_sc_hd__nand2_1
XANTENNA__12438__B2 _09152_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09571_ _10571_/B _10589_/A _08507_/B fanout51/X vssd1 vssd1 vccd1 vccd1 _09572_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_89_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08522_ _12802_/A _09238_/B _09440_/B1 _07896_/A vssd1 vssd1 vccd1 vccd1 _08523_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_77_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07314__B1 _12810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08453_ _08451_/A _08451_/B _08452_/Y vssd1 vssd1 vccd1 vccd1 _08710_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__07612__A _11269_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07404_ _10445_/A _12830_/A _12832_/A _10706_/B2 vssd1 vssd1 vccd1 vccd1 _07405_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout152_A _10707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08384_ _08384_/A _08384_/B vssd1 vssd1 vccd1 vccd1 _08422_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_116_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07335_ _12838_/A _10022_/B1 _12836_/A _10167_/A1 vssd1 vssd1 vccd1 vccd1 _07336_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07617__B2 _10948_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07617__A1 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07266_ _07267_/A _07267_/B _07267_/C vssd1 vssd1 vccd1 vccd1 _07268_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_33_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09005_ _09000_/A _09004_/Y _08590_/B vssd1 vssd1 vccd1 vccd1 _09006_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07197_ reg1_val[7] _07182_/B _07200_/A vssd1 vssd1 vccd1 vccd1 _07215_/B sky130_fd_sc_hd__o21a_1
XANTENNA__08162__B _09396_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10924__A1 _11653_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10924__B2 fanout66/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09907_ _09908_/A _09908_/B vssd1 vssd1 vccd1 vccd1 _09907_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_6_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12412__B _12412_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09838_ _11233_/S _11343_/B _09354_/B _06784_/B _09837_/X vssd1 vssd1 vccd1 vccd1
+ _09838_/X sky130_fd_sc_hd__o221a_1
XANTENNA__07506__B _12264_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10152__A2 fanout23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09769_ _12264_/B _09769_/B vssd1 vssd1 vccd1 vccd1 _09771_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_96_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11800_ _11800_/A _11800_/B vssd1 vssd1 vccd1 vccd1 _11802_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_68_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09845__A2 _09527_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07522__A _07522_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12780_ _12777_/A _12779_/B _12777_/B vssd1 vssd1 vccd1 vccd1 _12781_/B sky130_fd_sc_hd__a21bo_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11731_ _11725_/Y _11726_/X _11730_/X _11723_/X vssd1 vssd1 vccd1 vccd1 _11731_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_96_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11662_ _11663_/A _11663_/B vssd1 vssd1 vccd1 vccd1 _11664_/A sky130_fd_sc_hd__or2_1
XFILLER_0_22_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10613_ _10615_/A _10615_/B vssd1 vssd1 vccd1 vccd1 _10613_/X sky130_fd_sc_hd__or2_1
X_11593_ _11594_/A _11594_/B vssd1 vssd1 vccd1 vccd1 _11693_/A sky130_fd_sc_hd__or2_1
X_13332_ _13340_/CLK hold139/X vssd1 vssd1 vccd1 vccd1 hold137/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10544_ fanout74/X fanout59/X fanout56/X _10948_/B2 vssd1 vssd1 vccd1 vccd1 _10545_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08353__A _08745_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13157__A2 _06892_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13263_ _13357_/CLK hold46/X vssd1 vssd1 vccd1 vccd1 hold45/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09168__B _09170_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07509__C_N _07508_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12365__B1 _12316_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10475_ _10603_/B _10475_/B vssd1 vssd1 vccd1 vccd1 _10476_/B sky130_fd_sc_hd__nor2_2
X_13194_ hold252/A _13193_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13194_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_122_668 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12214_ _12214_/A _12214_/B _12214_/C vssd1 vssd1 vccd1 vccd1 _12215_/S sky130_fd_sc_hd__or3_1
XFILLER_0_121_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12145_ _12145_/A _12145_/B _12145_/C vssd1 vssd1 vccd1 vccd1 _12146_/B sky130_fd_sc_hd__or3_1
XFILLER_0_20_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12117__B1 _12244_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12076_ _12076_/A _12076_/B vssd1 vssd1 vccd1 vccd1 _12078_/B sky130_fd_sc_hd__xnor2_1
X_11027_ _09156_/Y _11003_/Y _11004_/X _11013_/X _11026_/Y vssd1 vssd1 vccd1 vccd1
+ _11027_/X sky130_fd_sc_hd__a311o_1
XANTENNA__09533__A1 _12423_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07135__C _07223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12978_ hold220/X _13004_/A2 _13006_/B1 hold230/X vssd1 vssd1 vccd1 vccd1 hold233/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09123__S _09142_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08528__A _08598_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11929_ _11929_/A _11929_/B vssd1 vssd1 vccd1 vccd1 _11931_/C sky130_fd_sc_hd__xnor2_1
XANTENNA_39 instruction[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_28 reg2_val[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_17 reg1_val[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07120_ reg1_val[3] _07120_/B vssd1 vssd1 vccd1 vccd1 _07120_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_55_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07051_ _08632_/A _08632_/B vssd1 vssd1 vccd1 vccd1 _09766_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_70_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09221__B1 _10022_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12513__A _12673_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09806__B _09808_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07953_ _07962_/B _07962_/A vssd1 vssd1 vccd1 vccd1 _07953_/X sky130_fd_sc_hd__and2b_1
X_06904_ instruction[11] _06884_/Y _06903_/X _06694_/B vssd1 vssd1 vccd1 vccd1 reg1_idx[0]
+ sky130_fd_sc_hd__o211a_4
XANTENNA__10134__A2 _09172_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07884_ _11271_/A _07072_/B _09768_/A1 vssd1 vssd1 vccd1 vccd1 _07886_/B sky130_fd_sc_hd__a21o_2
X_06835_ _06874_/B _06827_/Y _06834_/Y vssd1 vssd1 vccd1 vccd1 _06836_/B sky130_fd_sc_hd__o21ai_1
X_09623_ _09429_/A _09426_/Y _09428_/A vssd1 vssd1 vccd1 vccd1 _09624_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__07535__B1 _10413_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06766_ reg1_val[6] _07036_/A vssd1 vssd1 vccd1 vccd1 _06769_/A sky130_fd_sc_hd__nor2_1
XANTENNA__07342__A _09441_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09554_ fanout30/X _07089_/Y _10413_/A _07688_/B vssd1 vssd1 vccd1 vccd1 _09555_/B
+ sky130_fd_sc_hd__o22a_1
X_06697_ reg1_val[17] _07130_/A vssd1 vssd1 vccd1 vccd1 _06697_/X sky130_fd_sc_hd__and2_1
XFILLER_0_77_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08505_ _08506_/A _08506_/B vssd1 vssd1 vccd1 vccd1 _08505_/X sky130_fd_sc_hd__and2_1
X_09485_ _09706_/A _09485_/B _09649_/B _09953_/A vssd1 vssd1 vccd1 vccd1 _09485_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_53_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_13_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08436_ _08436_/A _08436_/B vssd1 vssd1 vccd1 vccd1 _08439_/B sky130_fd_sc_hd__or2_1
XFILLER_0_65_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08367_ _10949_/A _08414_/A vssd1 vssd1 vccd1 vccd1 _08368_/B sky130_fd_sc_hd__or2_1
XFILLER_0_18_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07318_ _07573_/A _07318_/B vssd1 vssd1 vccd1 vccd1 _07322_/A sky130_fd_sc_hd__or2_1
XFILLER_0_116_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08298_ _08298_/A _08298_/B vssd1 vssd1 vccd1 vccd1 _08300_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__08263__A1 _08730_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08263__B2 _08741_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07249_ _07249_/A _07249_/B vssd1 vssd1 vccd1 vccd1 _07300_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_6_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10208__A _10422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10260_ _06762_/B _09165_/X _10257_/Y _10258_/X vssd1 vssd1 vccd1 vccd1 _10260_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_103_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12423__A _12423_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10191_ _10192_/A _10192_/B _10192_/C vssd1 vssd1 vccd1 vccd1 _10193_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__08318__A2 _08741_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12901_ hold51/X hold242/X vssd1 vssd1 vccd1 vccd1 _12901_/X sky130_fd_sc_hd__and2b_1
XTAP_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12832_ _12832_/A _12856_/B vssd1 vssd1 vccd1 vccd1 _12832_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__13075__A1 _09716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12763_ reg1_val[28] _12782_/A vssd1 vssd1 vccd1 vccd1 _12773_/A sky130_fd_sc_hd__and2_1
XFILLER_0_29_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11714_ reg1_val[20] curr_PC[20] vssd1 vssd1 vccd1 vccd1 _11716_/A sky130_fd_sc_hd__or2_1
XFILLER_0_83_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_699 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12694_ _12695_/A _12695_/B _12695_/C vssd1 vssd1 vccd1 vccd1 _12701_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_71_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11645_ _11614_/X _11615_/Y _11618_/Y _11876_/A _11644_/X vssd1 vssd1 vccd1 vccd1
+ _11645_/X sky130_fd_sc_hd__a221o_1
XANTENNA__12050__A2 _07166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11576_ fanout29/X _11989_/A _12067_/A fanout27/X vssd1 vssd1 vccd1 vccd1 _11577_/B
+ sky130_fd_sc_hd__o22a_1
X_10527_ _10519_/Y _10520_/X _10526_/X vssd1 vssd1 vccd1 vccd1 _10527_/X sky130_fd_sc_hd__o21a_1
X_13315_ _13380_/CLK _13315_/D vssd1 vssd1 vccd1 vccd1 hold95/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13246_ hold53/X _06892_/B hold168/A _13246_/B2 vssd1 vssd1 vccd1 vccd1 _13246_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12338__B1 _11707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10458_ _10459_/A _10459_/B vssd1 vssd1 vccd1 vccd1 _10458_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_122_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13177_ hold263/X _12789_/B _13176_/X _12790_/A vssd1 vssd1 vccd1 vccd1 hold264/A
+ sky130_fd_sc_hd__a22o_1
X_10389_ _13290_/Q _10389_/B vssd1 vssd1 vccd1 vccd1 _10518_/B sky130_fd_sc_hd__or2_1
XANTENNA__07765__B1 _12818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12128_ _07169_/A _11343_/B _12254_/A1 _10113_/B _12127_/X vssd1 vssd1 vccd1 vccd1
+ _12128_/X sky130_fd_sc_hd__o221a_1
X_12059_ _12455_/S _12201_/C vssd1 vssd1 vccd1 vccd1 _12059_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__08309__A2 _08741_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06620_ _06621_/A _06621_/B vssd1 vssd1 vccd1 vccd1 _06647_/B sky130_fd_sc_hd__and2_1
XANTENNA__07162__A _09445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09270_ _11987_/A _09270_/B _09270_/C vssd1 vssd1 vccd1 vccd1 _09273_/C sky130_fd_sc_hd__and3_1
XFILLER_0_114_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08221_ _08745_/A _08221_/B vssd1 vssd1 vccd1 vccd1 _08225_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__13103__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08152_ _08722_/A _08152_/B vssd1 vssd1 vccd1 vccd1 _08159_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_125_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09993__B2 _09169_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07103_ _11269_/A _07103_/B vssd1 vssd1 vccd1 vccd1 _07636_/B sky130_fd_sc_hd__xnor2_1
X_08083_ _08081_/A _08081_/B _08082_/Y vssd1 vssd1 vccd1 vccd1 _08909_/B sky130_fd_sc_hd__a21boi_2
XFILLER_0_3_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08796__A2 fanout69/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07034_ _06774_/B _07050_/A _07050_/C _07223_/B vssd1 vssd1 vccd1 vccd1 _07036_/B
+ sky130_fd_sc_hd__a31o_4
XFILLER_0_70_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout115_A _08304_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11552__A1 _11142_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08985_ _08985_/A _08985_/B vssd1 vssd1 vccd1 vccd1 _09656_/C sky130_fd_sc_hd__nor2_1
X_07936_ _08727_/A2 _11558_/A _11751_/A _08727_/B1 vssd1 vssd1 vccd1 vccd1 _07937_/B
+ sky130_fd_sc_hd__o22a_2
X_07867_ _07878_/A _07878_/B vssd1 vssd1 vccd1 vccd1 _07867_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__06895__B _06896_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06818_ _10629_/A _06817_/Y _06740_/Y vssd1 vssd1 vccd1 vccd1 _06818_/X sky130_fd_sc_hd__o21a_1
XANTENNA__13057__A1 _07076_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09606_ _09606_/A _09606_/B vssd1 vssd1 vccd1 vccd1 _09607_/B sky130_fd_sc_hd__xor2_2
X_07798_ _06985_/A _06985_/B _10413_/A vssd1 vssd1 vccd1 vccd1 _07800_/B sky130_fd_sc_hd__a21oi_2
X_06749_ reg1_val[9] _07095_/A vssd1 vssd1 vccd1 vccd1 _06749_/Y sky130_fd_sc_hd__nand2_1
X_09537_ _09525_/Y _09526_/X _09534_/X _09536_/X vssd1 vssd1 vccd1 vccd1 _09537_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_78_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09468_ _09285_/A _09284_/B _09282_/Y vssd1 vssd1 vccd1 vccd1 _09478_/A sky130_fd_sc_hd__a21o_2
XANTENNA__07800__A _08724_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08419_ _08419_/A _08419_/B vssd1 vssd1 vccd1 vccd1 _08429_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_53_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09399_ _07033_/A _07033_/B _10664_/A vssd1 vssd1 vccd1 vccd1 _09401_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_46_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10830__A3 _12412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11430_ _11361_/Y _11649_/B _11429_/X vssd1 vssd1 vccd1 vccd1 _11430_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_104_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_363 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11361_ _11874_/A _11361_/B vssd1 vssd1 vccd1 vccd1 _11361_/Y sky130_fd_sc_hd__nand2_1
X_13100_ _13245_/A hold241/X vssd1 vssd1 vccd1 vccd1 _13349_/D sky130_fd_sc_hd__and2_1
X_10312_ _10312_/A _10312_/B vssd1 vssd1 vccd1 vccd1 _10314_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_104_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08631__A _09445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09736__A1 _10706_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11292_ _11292_/A _11292_/B _11292_/C vssd1 vssd1 vccd1 vccd1 _11293_/B sky130_fd_sc_hd__nor3_1
X_13031_ hold57/X _13236_/B _09594_/A _13077_/A2 _13030_/Y vssd1 vssd1 vccd1 vccd1
+ hold58/A sky130_fd_sc_hd__o221a_1
X_10243_ _06867_/B _10242_/X _11624_/A vssd1 vssd1 vccd1 vccd1 _10243_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__09736__B2 _10445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07747__B1 _11923_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11543__B2 _12254_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07247__A _09431_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07211__A2 _12830_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10174_ _10174_/A _10174_/B _10174_/C vssd1 vssd1 vccd1 vccd1 _10292_/B sky130_fd_sc_hd__and3_1
Xfanout192 _09083_/Y vssd1 vssd1 vccd1 vccd1 _09111_/S sky130_fd_sc_hd__buf_4
XANTENNA__06970__A1 _11343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout170 _07192_/Y vssd1 vssd1 vccd1 vccd1 _09568_/B sky130_fd_sc_hd__buf_8
Xfanout181 _12798_/A vssd1 vssd1 vccd1 vccd1 _07821_/A sky130_fd_sc_hd__buf_8
X_12815_ hold33/X _12818_/B _12814_/Y _13128_/A vssd1 vssd1 vccd1 vccd1 hold34/A sky130_fd_sc_hd__o211a_1
XFILLER_0_69_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08475__B2 _08739_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08475__A1 _07149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07710__A _11758_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12746_ _12746_/A _12746_/B _12746_/C _12746_/D vssd1 vssd1 vccd1 vccd1 _12746_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_29_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12677_ _12677_/A _12677_/B _12677_/C vssd1 vssd1 vccd1 vccd1 _12678_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_114_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11628_ _11532_/A _11532_/C _11532_/B vssd1 vssd1 vccd1 vccd1 _11629_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_107_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11559_ _11558_/A _12214_/B _11558_/C vssd1 vssd1 vccd1 vccd1 _11560_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_12_216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13229_ _13229_/A _13229_/B vssd1 vssd1 vccd1 vccd1 _13229_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__09356__B hold260/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12063__A _12261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09372__A _11142_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08770_ _08110_/A _08110_/B _08097_/Y vssd1 vssd1 vccd1 vccd1 _08774_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_18_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07721_ _08733_/A _07721_/B vssd1 vssd1 vccd1 vccd1 _07727_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__11837__A2 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08163__B1 _08216_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13039__A1 _10165_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07652_ _07656_/A _07656_/B vssd1 vssd1 vccd1 vccd1 _07652_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_125_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12247__C1 _12247_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06603_ reg1_val[27] _07144_/A vssd1 vssd1 vccd1 vccd1 _06606_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_88_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07583_ _07599_/A _07599_/B vssd1 vssd1 vccd1 vccd1 _07583_/X sky130_fd_sc_hd__and2b_1
X_09322_ _09108_/X _09110_/X _09336_/S vssd1 vssd1 vccd1 vccd1 _09322_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_47_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09253_ _09423_/B2 fanout9/A fanout5/X _12798_/A vssd1 vssd1 vccd1 vccd1 _09254_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_63_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07620__A _10448_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09184_ _09147_/X _09152_/Y _09183_/X _09151_/X vssd1 vssd1 vccd1 vccd1 _09184_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_90_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08218__B2 _12818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08204_ _08159_/A _08159_/B _08157_/X vssd1 vssd1 vccd1 vccd1 _08207_/B sky130_fd_sc_hd__o21ai_2
XFILLER_0_16_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08218__A1 fanout99/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10025__B2 _09433_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08135_ _08135_/A _08135_/B vssd1 vssd1 vccd1 vccd1 _08138_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_114_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08066_ _08809_/A _08809_/B vssd1 vssd1 vccd1 vccd1 _08848_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_101_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07017_ _07017_/A _12139_/A vssd1 vssd1 vccd1 vccd1 _07017_/X sky130_fd_sc_hd__or2_2
XFILLER_0_3_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09194__A2 fanout16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08968_ _08968_/A _08968_/B vssd1 vssd1 vccd1 vccd1 _08971_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_98_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08899_ _08899_/A _08899_/B vssd1 vssd1 vccd1 vccd1 _09049_/B sky130_fd_sc_hd__nor2_2
XANTENNA__11289__B1 fanout4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11828__A2 _12213_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07919_ _08742_/A _07919_/B vssd1 vssd1 vccd1 vccd1 _07923_/A sky130_fd_sc_hd__xnor2_2
X_10930_ _11171_/A _10930_/B vssd1 vssd1 vccd1 vccd1 _10931_/C sky130_fd_sc_hd__or2_1
XFILLER_0_85_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12600_ _12623_/A _12600_/B vssd1 vssd1 vccd1 vccd1 _12605_/D sky130_fd_sc_hd__xnor2_4
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10861_ _10739_/A _10861_/B _10861_/C _10861_/D vssd1 vssd1 vccd1 vccd1 _10862_/A
+ sky130_fd_sc_hd__and4b_1
XFILLER_0_14_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10792_ _10793_/A _10793_/B vssd1 vssd1 vccd1 vccd1 _10913_/B sky130_fd_sc_hd__nand2_1
XPHY_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12531_ _12537_/B _12531_/B vssd1 vssd1 vccd1 vccd1 new_PC[12] sky130_fd_sc_hd__and2_4
XFILLER_0_66_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12462_ reg1_val[3] curr_PC[3] _12622_/S vssd1 vssd1 vccd1 vccd1 _12464_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_81_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09406__B1 _10963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11413_ _11414_/A _11414_/B vssd1 vssd1 vccd1 vccd1 _11508_/B sky130_fd_sc_hd__nand2_1
XANTENNA__11987__A _11987_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12393_ reg1_val[30] _12429_/C vssd1 vssd1 vccd1 vccd1 _12393_/X sky130_fd_sc_hd__xor2_1
XANTENNA__12410__C1 _12455_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11344_ _06705_/X _11973_/B _11342_/Y _06707_/B _11343_/Y vssd1 vssd1 vccd1 vccd1
+ _11344_/X sky130_fd_sc_hd__a221o_2
XFILLER_0_120_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11275_ _11275_/A _11275_/B vssd1 vssd1 vccd1 vccd1 _11288_/A sky130_fd_sc_hd__xnor2_1
X_13014_ hold180/X _13016_/A2 _13016_/B1 hold195/X vssd1 vssd1 vccd1 vccd1 hold224/A
+ sky130_fd_sc_hd__a22o_1
X_10226_ _10227_/A _10227_/B vssd1 vssd1 vccd1 vccd1 _10226_/X sky130_fd_sc_hd__and2_1
Xhold4 hold4/A vssd1 vssd1 vccd1 vccd1 hold4/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10157_ _12076_/A _10157_/B vssd1 vssd1 vccd1 vccd1 _10159_/B sky130_fd_sc_hd__xnor2_1
X_10088_ _10088_/A _10088_/B vssd1 vssd1 vccd1 vccd1 _10090_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__07705__A _12210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09920__A _12138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09893__B1 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08536__A _08745_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09131__S _09142_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12729_ _12729_/A _12729_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[20] sky130_fd_sc_hd__nor2_8
XFILLER_0_127_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_758 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10558__A2 fanout30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07423__A2 _09238_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_396 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09940_ _09940_/A _09940_/B vssd1 vssd1 vccd1 vccd1 _09941_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_96_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09871_ _09871_/A _09871_/B vssd1 vssd1 vccd1 vccd1 _09932_/A sky130_fd_sc_hd__xor2_4
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06934__A1 _12341_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08822_ _08749_/A _08749_/B _08737_/X vssd1 vssd1 vccd1 vccd1 _08825_/A sky130_fd_sc_hd__a21oi_2
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08753_ _11758_/A _08753_/B vssd1 vssd1 vccd1 vccd1 _08755_/B sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout182_A _12798_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07704_ _12210_/A _07705_/B vssd1 vssd1 vccd1 vccd1 _07704_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__08136__B1 _09396_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08684_ _08685_/B vssd1 vssd1 vccd1 vccd1 _08684_/Y sky130_fd_sc_hd__inv_2
XTAP_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07635_ _07627_/A _08918_/A _07669_/B vssd1 vssd1 vccd1 vccd1 _07635_/X sky130_fd_sc_hd__o21ba_1
X_07566_ _07566_/A _07566_/B vssd1 vssd1 vccd1 vccd1 _07567_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_76_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09305_ _09706_/A _09649_/B _09071_/X _09304_/B _09304_/A vssd1 vssd1 vccd1 vccd1
+ _09307_/A sky130_fd_sc_hd__o32a_1
X_07497_ _07149_/A _12412_/A _09442_/A vssd1 vssd1 vccd1 vccd1 _07499_/B sky130_fd_sc_hd__a21oi_2
X_09236_ _09444_/A _12854_/A fanout7/X _09236_/B2 vssd1 vssd1 vccd1 vccd1 _09237_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_35_138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08165__B _09396_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09167_ _09168_/A _09170_/A vssd1 vssd1 vccd1 vccd1 _09167_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_44_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09098_ _09094_/X _09097_/X _09663_/S vssd1 vssd1 vccd1 vccd1 _09098_/X sky130_fd_sc_hd__mux2_1
X_08118_ _08119_/A _08119_/B vssd1 vssd1 vccd1 vccd1 _08118_/X sky130_fd_sc_hd__or2_1
XANTENNA__08181__A _08733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07509__B _12316_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08049_ _08844_/A _08049_/B vssd1 vssd1 vccd1 vccd1 _08069_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_102_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11060_ _11061_/A _11061_/B vssd1 vssd1 vccd1 vccd1 _11196_/B sky130_fd_sc_hd__and2_1
XANTENNA_fanout95_A _07076_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10011_ fanout59/X _10589_/A _08507_/B _10941_/B vssd1 vssd1 vccd1 vccd1 _10012_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_98_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12150__B _12261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08127__B1 _08727_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11962_ _11962_/A _11962_/B vssd1 vssd1 vccd1 vccd1 _11964_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09875__B1 fanout66/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11893_ hold225/A _11450_/B _11966_/B _11968_/B1 vssd1 vssd1 vccd1 vccd1 _11893_/X
+ sky130_fd_sc_hd__a31o_1
X_10913_ _10913_/A _10913_/B _10913_/C vssd1 vssd1 vccd1 vccd1 _10914_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_39_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10844_ _10844_/A _10844_/B _10842_/Y vssd1 vssd1 vccd1 vccd1 _10845_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_27_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10775_ _12254_/A1 _10762_/X _10774_/Y _10113_/A _10773_/X vssd1 vssd1 vccd1 vccd1
+ _10775_/Y sky130_fd_sc_hd__o221ai_1
X_12514_ _12523_/A _12514_/B vssd1 vssd1 vccd1 vccd1 _12516_/C sky130_fd_sc_hd__nand2_1
XANTENNA__07102__B2 _10571_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07102__A1 _10413_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07653__A2 _11989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12445_ _12626_/B _12446_/B vssd1 vssd1 vccd1 vccd1 _12453_/A sky130_fd_sc_hd__nand2_1
XANTENNA__11737__A1 _11142_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08602__A1 _08673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12376_ _12376_/A _12376_/B vssd1 vssd1 vccd1 vccd1 _12413_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_120_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08602__B2 _08671_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11327_ _11792_/A _11328_/B _11328_/C vssd1 vssd1 vccd1 vccd1 _11327_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_1_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09915__A _12808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11258_ _09614_/A _12150_/A _12067_/A _09613_/A vssd1 vssd1 vccd1 vccd1 _11259_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12341__A _12341_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11189_ _11188_/B _11188_/C _11188_/A vssd1 vssd1 vccd1 vccd1 _11190_/B sky130_fd_sc_hd__a21o_1
X_10209_ _10209_/A _10209_/B vssd1 vssd1 vccd1 vccd1 _10211_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__09126__S _09127_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07154__B _07154_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11122__C1 _09172_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07341__A1 _12846_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07341__B2 _09238_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07420_ _07420_/A _07420_/B vssd1 vssd1 vccd1 vccd1 fanout8/A sky130_fd_sc_hd__or2_1
XFILLER_0_15_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07351_ _10445_/A _12828_/A _12830_/A _10706_/B2 vssd1 vssd1 vccd1 vccd1 _07352_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_128_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11976__B2 _12254_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07282_ _12794_/A _07282_/B vssd1 vssd1 vccd1 vccd1 _07293_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_122_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09021_ _09021_/A _09021_/B vssd1 vssd1 vccd1 vccd1 _11221_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_31_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold201 hold201/A vssd1 vssd1 vccd1 vccd1 hold201/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13111__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold223 hold223/A vssd1 vssd1 vccd1 vccd1 hold223/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold212 hold212/A vssd1 vssd1 vccd1 vccd1 hold212/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold234 hold234/A vssd1 vssd1 vccd1 vccd1 hold234/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10400__A1 _12254_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold278 hold278/A vssd1 vssd1 vccd1 vccd1 hold278/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold267 hold267/A vssd1 vssd1 vccd1 vccd1 hold267/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold256 hold256/A vssd1 vssd1 vccd1 vccd1 hold256/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold245 hold245/A vssd1 vssd1 vccd1 vccd1 hold245/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10400__B2 _06924_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10036__A _10959_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold289 hold289/A vssd1 vssd1 vccd1 vccd1 hold289/X sky130_fd_sc_hd__dlygate4sd3_1
X_09923_ _09923_/A _09923_/B _09923_/C vssd1 vssd1 vccd1 vccd1 _10056_/B sky130_fd_sc_hd__and3_1
XFILLER_0_1_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09854_ _10748_/A _09854_/B vssd1 vssd1 vccd1 vccd1 _09958_/A sky130_fd_sc_hd__or2_1
XFILLER_0_0_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11900__A1 _12290_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08805_ _08805_/A _08805_/B vssd1 vssd1 vccd1 vccd1 _08806_/B sky130_fd_sc_hd__nor2_1
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09785_ _09786_/A _09786_/B vssd1 vssd1 vccd1 vccd1 _09785_/Y sky130_fd_sc_hd__nand2_1
X_06997_ reg1_val[18] reg1_val[19] _06997_/C vssd1 vssd1 vccd1 vccd1 _12726_/B sky130_fd_sc_hd__or3_4
XANTENNA__07064__B _07064_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08736_ _08736_/A _08736_/B vssd1 vssd1 vccd1 vccd1 _08738_/B sky130_fd_sc_hd__xnor2_1
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08667_ _08669_/B _08667_/B vssd1 vssd1 vccd1 vccd1 _08670_/A sky130_fd_sc_hd__and2b_1
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07618_ _11163_/A _07618_/B vssd1 vssd1 vccd1 vccd1 _07621_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__12208__A2 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07080__A _07080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08598_ _08598_/A _08598_/B vssd1 vssd1 vccd1 vccd1 _08627_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__08176__A _08731_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07549_ _07552_/B _07552_/A vssd1 vssd1 vccd1 vccd1 _07549_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_64_723 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10560_ _10561_/B _10560_/B vssd1 vssd1 vccd1 vccd1 _10562_/A sky130_fd_sc_hd__and2b_1
XANTENNA_fanout10_A fanout9/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09219_ _09220_/A _09220_/B vssd1 vssd1 vccd1 vccd1 _09415_/A sky130_fd_sc_hd__nor2_1
X_10491_ _10493_/B _10493_/A vssd1 vssd1 vccd1 vccd1 _10491_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_23_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12230_ _12414_/A _12230_/B vssd1 vssd1 vccd1 vccd1 _12286_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_16_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10942__A2 _07154_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12161_ _12017_/X _12092_/Y _12094_/B vssd1 vssd1 vccd1 vccd1 _12161_/Y sky130_fd_sc_hd__o21ai_1
X_11112_ _11111_/A _11111_/B _11111_/Y _09156_/Y vssd1 vssd1 vccd1 vccd1 _11137_/A
+ sky130_fd_sc_hd__o211a_1
XANTENNA__09735__A _10710_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12092_ _12094_/A vssd1 vssd1 vccd1 vccd1 _12092_/Y sky130_fd_sc_hd__inv_2
X_11043_ _10448_/A _06986_/B _12412_/A _11163_/A vssd1 vssd1 vccd1 vccd1 _11043_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_36_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12994_ hold174/X _13004_/A2 _13006_/B1 _13300_/Q vssd1 vssd1 vccd1 vccd1 hold175/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_98_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11945_ _11781_/A _11863_/A _11862_/A vssd1 vssd1 vccd1 vccd1 _11945_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_98_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11876_ _11876_/A _11876_/B vssd1 vssd1 vccd1 vccd1 _11876_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_27_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10827_ fanout74/X _09568_/A fanout13/X _10948_/B2 vssd1 vssd1 vccd1 vccd1 _10828_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_27_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10758_ _10632_/X _10636_/X _10754_/X _10756_/Y vssd1 vssd1 vccd1 vccd1 _10759_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12428_ _12428_/A _12428_/B _12428_/C vssd1 vssd1 vccd1 vccd1 _12428_/X sky130_fd_sc_hd__and3_1
X_10689_ _10689_/A _10689_/B vssd1 vssd1 vccd1 vccd1 _10693_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_23_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12359_ _06621_/A _09354_/B _12358_/Y _06619_/Y _11343_/B vssd1 vssd1 vccd1 vccd1
+ _12359_/X sky130_fd_sc_hd__o221a_1
XANTENNA__07149__B _09343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08051__A2 _08741_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11894__B _11973_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06920_ instruction[21] _06884_/Y _06919_/X _06694_/B vssd1 vssd1 vccd1 vccd1 reg2_idx[3]
+ sky130_fd_sc_hd__o211a_4
XANTENNA__12135__A1 _06881_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12071__A _12317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06851_ _08980_/B _06851_/B vssd1 vssd1 vccd1 vccd1 _06853_/C sky130_fd_sc_hd__nor2_1
XANTENNA__06770__C1 _12654_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06782_ reg1_val[4] _10252_/S vssd1 vssd1 vccd1 vccd1 _06782_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_89_130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09570_ _10165_/A _09570_/B _09570_/C vssd1 vssd1 vccd1 vccd1 _09573_/B sky130_fd_sc_hd__nand3_1
XANTENNA__12843__C1 _13214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08521_ _08521_/A _08521_/B vssd1 vssd1 vccd1 vccd1 _08538_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_77_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07314__A1 _10574_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08452_ _08487_/B _08487_/A vssd1 vssd1 vccd1 vccd1 _08452_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__07314__B2 _10575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12362__D_N _12361_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07403_ _07401_/A _07401_/B _07402_/Y vssd1 vssd1 vccd1 vccd1 _07598_/A sky130_fd_sc_hd__a21bo_2
XFILLER_0_58_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout145_A _09768_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08383_ _08383_/A _08383_/B vssd1 vssd1 vccd1 vccd1 _08384_/B sky130_fd_sc_hd__or2_1
XFILLER_0_18_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07334_ _07334_/A _07334_/B vssd1 vssd1 vccd1 vccd1 _07337_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_42_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07617__A2 _10818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08724__A _08724_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07265_ _12138_/A _07265_/B vssd1 vssd1 vccd1 vccd1 _07267_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_45_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09004_ _09004_/A _09004_/B vssd1 vssd1 vccd1 vccd1 _09004_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_5_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07196_ _10165_/A _07196_/B vssd1 vssd1 vccd1 vccd1 _07214_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_41_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07250__B1 _12834_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09555__A _11673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10924__A2 _10571_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12126__A1 _09354_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09906_ _09906_/A _09906_/B vssd1 vssd1 vccd1 vccd1 _09908_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_1_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09837_ _09837_/A _09837_/B _09837_/C vssd1 vssd1 vccd1 vccd1 _09837_/X sky130_fd_sc_hd__or3_2
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09768_ _09768_/A1 fanout9/A fanout5/X _07026_/X vssd1 vssd1 vccd1 vccd1 _09769_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08750__B1 _08216_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08719_ _08295_/Y _08719_/B vssd1 vssd1 vccd1 vccd1 _09036_/A sky130_fd_sc_hd__and2b_1
XANTENNA_fanout58_A fanout59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11730_ _10113_/A _10762_/X _10774_/Y _12254_/A1 _11729_/X vssd1 vssd1 vccd1 vccd1
+ _11730_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_95_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08502__B1 _08617_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09699_ _09699_/A _09699_/B _09699_/C _09699_/D vssd1 vssd1 vccd1 vccd1 _09699_/X
+ sky130_fd_sc_hd__or4_2
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11661_ _11661_/A _11661_/B vssd1 vssd1 vccd1 vccd1 _11663_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_64_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11592_ _11495_/A _11495_/B _11496_/Y vssd1 vssd1 vccd1 vccd1 _11594_/B sky130_fd_sc_hd__a21boi_1
X_10612_ _10612_/A _10612_/B vssd1 vssd1 vccd1 vccd1 _10615_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__12062__B1 fanout4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13331_ _13355_/CLK hold78/X vssd1 vssd1 vccd1 vccd1 _13331_/Q sky130_fd_sc_hd__dfxtp_1
X_10543_ _10543_/A _10543_/B vssd1 vssd1 vccd1 vccd1 _10546_/A sky130_fd_sc_hd__or2_2
XFILLER_0_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13262_ _13357_/CLK hold38/X vssd1 vssd1 vccd1 vccd1 hold37/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12365__A1 _10928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10474_ _10474_/A _10474_/B _10474_/C vssd1 vssd1 vccd1 vccd1 _10475_/B sky130_fd_sc_hd__and3_1
X_13193_ _13193_/A _13193_/B vssd1 vssd1 vccd1 vccd1 _13193_/Y sky130_fd_sc_hd__xnor2_1
X_12213_ _12213_/A _12214_/B vssd1 vssd1 vccd1 vccd1 _12213_/Y sky130_fd_sc_hd__nor2_1
X_12144_ _12145_/A _12145_/B _12145_/C vssd1 vssd1 vccd1 vccd1 _12146_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_20_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06595__A2 _06587_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06601__B _12686_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12075_ fanout29/X fanout12/X fanout8/X fanout27/X vssd1 vssd1 vccd1 vccd1 _12076_/B
+ sky130_fd_sc_hd__o22a_1
X_11026_ _12254_/A1 _11012_/B _11025_/X vssd1 vssd1 vccd1 vccd1 _11026_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_2_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08741__B1 _08617_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07135__D _07135_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12977_ _13013_/A hold221/X vssd1 vssd1 vccd1 vccd1 hold222/A sky130_fd_sc_hd__and2_1
X_11928_ _11926_/Y _11928_/B vssd1 vssd1 vccd1 vccd1 _11929_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_28_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11859_ _11859_/A _11859_/B vssd1 vssd1 vccd1 vccd1 _11861_/C sky130_fd_sc_hd__xor2_1
XANTENNA_29 reg2_val[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_18 reg1_val[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07050_ _07050_/A _07223_/B _07050_/C vssd1 vssd1 vccd1 vccd1 _08632_/B sky130_fd_sc_hd__or3_2
XFILLER_0_70_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09221__A1 _12842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09221__B2 _12844_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_166 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07952_ _08033_/A _08033_/B _07948_/Y vssd1 vssd1 vccd1 vccd1 _07962_/B sky130_fd_sc_hd__o21ba_1
X_06903_ instruction[18] _06921_/B vssd1 vssd1 vccd1 vccd1 _06903_/X sky130_fd_sc_hd__or2_1
XANTENNA__07535__A1 _07033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07883_ _08722_/A _07883_/B vssd1 vssd1 vccd1 vccd1 _07889_/A sky130_fd_sc_hd__xnor2_1
X_06834_ reg1_val[23] _07194_/A _06833_/Y vssd1 vssd1 vccd1 vccd1 _06834_/Y sky130_fd_sc_hd__a21oi_1
X_09622_ _09622_/A _09622_/B vssd1 vssd1 vccd1 vccd1 _09624_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__08732__B1 _08656_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09314__S _09351_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09553_ _09553_/A _09553_/B vssd1 vssd1 vccd1 vccd1 _09556_/A sky130_fd_sc_hd__nand2_1
XANTENNA__13084__A2 _06572_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06765_ _07036_/A reg1_val[6] vssd1 vssd1 vccd1 vccd1 _06765_/Y sky130_fd_sc_hd__nand2b_1
X_08504_ _08521_/A _08521_/B _08500_/X vssd1 vssd1 vccd1 vccd1 _08506_/B sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout262_A _12455_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12831__A2 _12818_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06696_ reg2_val[17] _06720_/B _06703_/B1 _06695_/Y vssd1 vssd1 vccd1 vccd1 _07130_/A
+ sky130_fd_sc_hd__o2bb2a_4
XFILLER_0_77_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09484_ _09484_/A _09484_/B vssd1 vssd1 vccd1 vccd1 _09953_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_77_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08435_ _08449_/A _08449_/B vssd1 vssd1 vccd1 vccd1 _08435_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_19_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08366_ _10949_/A _08414_/A vssd1 vssd1 vccd1 vccd1 _08366_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_46_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07317_ _07317_/A _07317_/B vssd1 vssd1 vccd1 vccd1 _07318_/B sky130_fd_sc_hd__nor2_1
XANTENNA__09269__B _10664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08263__A2 _08732_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08297_ _08297_/A _08297_/B vssd1 vssd1 vccd1 vccd1 _08300_/A sky130_fd_sc_hd__nand2_1
X_07248_ _07249_/A _07249_/B vssd1 vssd1 vccd1 vccd1 _07267_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_61_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07179_ _08741_/B2 _10948_/B2 _10963_/A fanout74/X vssd1 vssd1 vccd1 vccd1 _07180_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_103_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10190_ _10190_/A _10190_/B vssd1 vssd1 vccd1 vccd1 _10192_/C sky130_fd_sc_hd__xnor2_1
X_12900_ hold294/A hold55/X vssd1 vssd1 vccd1 vccd1 _13124_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__08723__B1 _08723_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12831_ hold47/X _12818_/B _12830_/Y _13235_/A vssd1 vssd1 vccd1 vccd1 hold48/A sky130_fd_sc_hd__o211a_1
XTAP_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12807__C1 _13128_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12762_ reg1_val[28] _12782_/A vssd1 vssd1 vccd1 vccd1 _12764_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_29_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11713_ _06676_/C _11711_/X _11712_/Y vssd1 vssd1 vccd1 vccd1 _11713_/X sky130_fd_sc_hd__a21o_1
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12693_ _12693_/A _12701_/A vssd1 vssd1 vccd1 vccd1 _12695_/C sky130_fd_sc_hd__nand2_1
X_11644_ _11644_/A _11644_/B _11624_/X vssd1 vssd1 vccd1 vccd1 _11644_/X sky130_fd_sc_hd__or3b_2
XANTENNA__12035__B1 _11624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11575_ _11575_/A _11575_/B vssd1 vssd1 vccd1 vccd1 _11579_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13314_ _13314_/CLK hold120/X vssd1 vssd1 vccd1 vccd1 hold118/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10526_ _06750_/A _10521_/Y _10523_/Y _10524_/X _10525_/Y vssd1 vssd1 vccd1 vccd1
+ _10526_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_24_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13245_ _13245_/A _13245_/B hold102/X vssd1 vssd1 vccd1 vccd1 hold103/A sky130_fd_sc_hd__and3_1
X_10457_ _10457_/A _10457_/B vssd1 vssd1 vccd1 vccd1 _10459_/B sky130_fd_sc_hd__or2_1
XFILLER_0_122_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06637__A_N _07140_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09195__A _09548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07708__A _11385_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13176_ hold277/A _13175_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13176_/X sky130_fd_sc_hd__mux2_1
X_10388_ _10384_/Y _10387_/Y _11886_/A vssd1 vssd1 vccd1 vccd1 _10388_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_58_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07765__B2 _08304_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07765__A1 fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12127_ _12307_/B1 _12126_/X _06633_/B vssd1 vssd1 vccd1 vccd1 _12127_/X sky130_fd_sc_hd__a21o_1
X_12058_ curr_PC[24] _12058_/B vssd1 vssd1 vccd1 vccd1 _12201_/C sky130_fd_sc_hd__and2_2
X_11009_ _11009_/A _11009_/B vssd1 vssd1 vccd1 vccd1 _11009_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_74_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09134__S _09142_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07443__A _09716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08220_ _07885_/B _08744_/A2 _08564_/B _08721_/B1 vssd1 vssd1 vccd1 vccd1 _08221_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_114_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08274__A _08742_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10309__A _10928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08151_ _10537_/A1 _07896_/A _08723_/B1 _08432_/B vssd1 vssd1 vccd1 vccd1 _08152_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_70_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07102_ _10413_/A _10570_/A _10567_/A _10571_/A vssd1 vssd1 vccd1 vccd1 _07103_/B
+ sky130_fd_sc_hd__o22a_1
X_08082_ _08900_/B _08900_/A vssd1 vssd1 vccd1 vccd1 _08082_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_31_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07033_ _07033_/A _07033_/B vssd1 vssd1 vccd1 vccd1 _07033_/X sky130_fd_sc_hd__and2_1
XFILLER_0_31_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07618__A _11163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout108_A _12073_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08984_ _08984_/A _08984_/B vssd1 vssd1 vccd1 vccd1 _08985_/B sky130_fd_sc_hd__and2_1
XFILLER_0_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07935_ _07938_/A _07938_/B vssd1 vssd1 vccd1 vccd1 _07935_/Y sky130_fd_sc_hd__nor2_1
X_09605_ _09606_/A _09606_/B vssd1 vssd1 vccd1 vccd1 _09605_/X sky130_fd_sc_hd__and2_1
X_07866_ _07912_/A _07865_/Y _07861_/Y vssd1 vssd1 vccd1 vccd1 _07878_/B sky130_fd_sc_hd__a21o_1
X_06817_ _10507_/A _06816_/X _06746_/X vssd1 vssd1 vccd1 vccd1 _06817_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__13057__A2 _13087_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07797_ _08740_/A _07797_/B vssd1 vssd1 vccd1 vccd1 _07805_/A sky130_fd_sc_hd__xnor2_1
X_09536_ _09520_/Y _09521_/X _09527_/X _09535_/X vssd1 vssd1 vccd1 vccd1 _09536_/X
+ sky130_fd_sc_hd__o211a_1
X_06748_ reg1_val[9] _07095_/A vssd1 vssd1 vccd1 vccd1 _06750_/B sky130_fd_sc_hd__and2_1
X_09467_ _09467_/A _09467_/B vssd1 vssd1 vccd1 vccd1 _09480_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_66_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06679_ reg2_val[19] _06720_/B _06596_/Y _06678_/Y vssd1 vssd1 vccd1 vccd1 _07210_/A
+ sky130_fd_sc_hd__o2bb2a_2
X_08418_ _08444_/A _08415_/B _08417_/X vssd1 vssd1 vccd1 vccd1 _08429_/A sky130_fd_sc_hd__o21ba_1
XFILLER_0_38_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07692__B1 _07819_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09398_ _09397_/B _09397_/C _09746_/A vssd1 vssd1 vccd1 vccd1 _09404_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__07800__B _07800_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08349_ _08349_/A _08349_/B vssd1 vssd1 vccd1 vccd1 _08376_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_117_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11360_ _11360_/A _11649_/A vssd1 vssd1 vccd1 vccd1 _11361_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_34_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10311_ _10312_/A _10312_/B vssd1 vssd1 vccd1 vccd1 _10471_/A sky130_fd_sc_hd__nor2_1
X_13030_ _06571_/Y _06572_/A rst vssd1 vssd1 vccd1 vccd1 _13030_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_14_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11291_ _11292_/A _11292_/B _11292_/C vssd1 vssd1 vccd1 vccd1 _11293_/A sky130_fd_sc_hd__o21a_1
X_10242_ _06814_/Y _10241_/Y _12388_/S vssd1 vssd1 vccd1 vccd1 _10242_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09736__A2 _10571_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07747__A1 _06574_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11543__A2 _11012_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07747__B2 _08436_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10173_ _10172_/B _10172_/C _10172_/A vssd1 vssd1 vccd1 vccd1 _10174_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout182 _12798_/A vssd1 vssd1 vccd1 vccd1 _08646_/B2 sky130_fd_sc_hd__clkbuf_4
Xfanout171 _09440_/B1 vssd1 vssd1 vccd1 vccd1 _08656_/B sky130_fd_sc_hd__buf_6
Xfanout160 _09653_/A vssd1 vssd1 vccd1 vccd1 _12170_/A sky130_fd_sc_hd__buf_4
XFILLER_0_88_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08359__A _08681_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout193 _09433_/A vssd1 vssd1 vccd1 vccd1 _08742_/A sky130_fd_sc_hd__buf_12
XANTENNA__07263__A _12076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13048__A2 _12788_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12814_ _12814_/A _12818_/B vssd1 vssd1 vccd1 vccd1 _12814_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_97_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12256__B1 _12255_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12745_ _12745_/A _12750_/A vssd1 vssd1 vccd1 vccd1 _12749_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_84_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08475__A2 _08436_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12676_ _12677_/A _12677_/C _12677_/B vssd1 vssd1 vccd1 vccd1 _12683_/B sky130_fd_sc_hd__a21o_1
XANTENNA__08094__A _08745_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11627_ _11627_/A _11627_/B vssd1 vssd1 vccd1 vccd1 _11629_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_37_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07435__B1 _10022_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09918__A _12804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11558_ _11558_/A _12214_/B _11558_/C vssd1 vssd1 vccd1 vccd1 _11682_/B sky130_fd_sc_hd__or3_1
XFILLER_0_123_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10509_ _10384_/A _10381_/Y _10383_/B vssd1 vssd1 vccd1 vccd1 _10513_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_80_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09129__S _09669_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11489_ _11489_/A _11489_/B vssd1 vssd1 vccd1 vccd1 _11503_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_122_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13228_ _13235_/A _13228_/B vssd1 vssd1 vccd1 vccd1 _13376_/D sky130_fd_sc_hd__and2_1
XFILLER_0_0_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13159_ _12885_/X _13159_/B vssd1 vssd1 vccd1 vccd1 _13160_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_85_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07720_ _08732_/A2 _11751_/A _11766_/A _08656_/B vssd1 vssd1 vccd1 vccd1 _07721_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10799__A _10959_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08163__A1 _08798_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
X_07651_ _08731_/A _07651_/B vssd1 vssd1 vccd1 vccd1 _07656_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__08163__B2 _07821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06602_ reg2_val[27] _06771_/A _06596_/Y _06601_/Y vssd1 vssd1 vccd1 vccd1 _07144_/A
+ sky130_fd_sc_hd__o2bb2a_4
XFILLER_0_94_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07582_ _07582_/A _07582_/B vssd1 vssd1 vccd1 vccd1 _07599_/B sky130_fd_sc_hd__xnor2_2
X_09321_ _09104_/X _09107_/X _09330_/S vssd1 vssd1 vccd1 vccd1 _09321_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_88_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12519__A _12680_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09252_ _07500_/A _07500_/B _07498_/X vssd1 vssd1 vccd1 vccd1 _09256_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_7_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09183_ _09108_/S _12430_/A _09171_/X _09161_/Y vssd1 vssd1 vccd1 vccd1 _09183_/X
+ sky130_fd_sc_hd__a211o_1
X_08203_ _08150_/A _08149_/B _08147_/Y vssd1 vssd1 vccd1 vccd1 _08207_/A sky130_fd_sc_hd__a21o_1
XANTENNA__08218__A2 _08732_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10025__A2 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout225_A _12794_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08134_ _08135_/A _08135_/B vssd1 vssd1 vccd1 vccd1 _08134_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_71_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08065_ _08724_/A _08065_/B vssd1 vssd1 vccd1 vccd1 _08809_/B sky130_fd_sc_hd__xnor2_1
X_07016_ _10248_/S _07016_/B vssd1 vssd1 vccd1 vccd1 _07016_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_101_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08967_ _08960_/A _08960_/B _08961_/X vssd1 vssd1 vccd1 vccd1 _08971_/A sky130_fd_sc_hd__a21o_2
X_08898_ _08898_/A _08898_/B _08898_/C vssd1 vssd1 vccd1 vccd1 _08899_/B sky130_fd_sc_hd__and3_1
XANTENNA__11289__A1 _09745_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11289__B2 _10418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07918_ _08732_/A1 _08741_/A2 _08617_/B _10927_/A1 vssd1 vssd1 vccd1 vccd1 _07919_/B
+ sky130_fd_sc_hd__o22a_1
X_07849_ _07824_/B _07824_/C _07824_/A vssd1 vssd1 vccd1 vccd1 _07849_/Y sky130_fd_sc_hd__a21oi_1
X_10860_ _11102_/A _11102_/B vssd1 vssd1 vccd1 vccd1 _10861_/B sky130_fd_sc_hd__nor2_1
X_09519_ hold248/A hold290/A vssd1 vssd1 vccd1 vccd1 _09519_/X sky130_fd_sc_hd__or2_1
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10791_ _11269_/A _10791_/B vssd1 vssd1 vccd1 vccd1 _10793_/B sky130_fd_sc_hd__xnor2_1
XPHY_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12530_ _12530_/A _12530_/B _12530_/C vssd1 vssd1 vccd1 vccd1 _12531_/B sky130_fd_sc_hd__nand3_1
X_12461_ _12467_/B _12461_/B vssd1 vssd1 vccd1 vccd1 new_PC[2] sky130_fd_sc_hd__and2_4
XANTENNA__09406__A1 _11065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09406__B2 _11653_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11412_ _11412_/A _11412_/B vssd1 vssd1 vccd1 vccd1 _11414_/B sky130_fd_sc_hd__xor2_2
XANTENNA__08642__A _09897_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12392_ _12392_/A _12392_/B vssd1 vssd1 vccd1 vccd1 _12392_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_62_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11987__B _11987_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11343_ _11343_/A _11343_/B vssd1 vssd1 vccd1 vccd1 _11343_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_120_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11274_ _11392_/A _11274_/B vssd1 vssd1 vccd1 vccd1 _11275_/B sky130_fd_sc_hd__nor2_1
X_13013_ _13013_/A hold181/X vssd1 vssd1 vccd1 vccd1 hold182/A sky130_fd_sc_hd__and2_1
X_10225_ _10225_/A _10225_/B vssd1 vssd1 vccd1 vccd1 _10227_/B sky130_fd_sc_hd__xor2_4
XANTENNA__09590__B1 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10156_ fanout29/X _10818_/A _10963_/A _07688_/B vssd1 vssd1 vccd1 vccd1 _10157_/B
+ sky130_fd_sc_hd__o22a_1
Xhold5 hold5/A vssd1 vssd1 vccd1 vccd1 hold5/X sky130_fd_sc_hd__dlygate4sd3_1
X_10087_ _09940_/A _09940_/B _09938_/Y vssd1 vssd1 vccd1 vccd1 _10088_/B sky130_fd_sc_hd__a21oi_4
XANTENNA__08089__A _08745_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09893__A1 _09567_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09893__B2 _07192_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07721__A _08733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10989_ _10735_/X _10857_/Y _10858_/X vssd1 vssd1 vccd1 vccd1 _10989_/Y sky130_fd_sc_hd__a21oi_1
X_12728_ _12746_/A _12728_/B _12728_/C vssd1 vssd1 vccd1 vccd1 _12729_/B sky130_fd_sc_hd__and3_2
XFILLER_0_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12659_ reg1_val[7] _12659_/B vssd1 vssd1 vccd1 vccd1 _12660_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_127_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09870_ _09870_/A _09870_/B vssd1 vssd1 vccd1 vccd1 _09871_/B sky130_fd_sc_hd__nand2_2
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12802__A _12802_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09383__A _09716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09581__B1 _11558_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08821_ _11758_/A _08763_/B _08766_/A vssd1 vssd1 vccd1 vccd1 _08826_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_29_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08752_ _08752_/A _08752_/B vssd1 vssd1 vccd1 vccd1 _08753_/B sky130_fd_sc_hd__nor2_1
XANTENNA__08136__A1 _08752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08683_ _08683_/A _08683_/B vssd1 vssd1 vccd1 vccd1 _08685_/B sky130_fd_sc_hd__xor2_1
X_07703_ _07703_/A _07703_/B vssd1 vssd1 vccd1 vccd1 _07705_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__08136__B2 _08798_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07634_ _08919_/A _08919_/B _07630_/X vssd1 vssd1 vccd1 vccd1 _07669_/B sky130_fd_sc_hd__a21oi_1
XTAP_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07895__B1 _07955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07565_ _07566_/A _07566_/B vssd1 vssd1 vccd1 vccd1 _07565_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_75_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07496_ _09897_/A _07496_/B vssd1 vssd1 vccd1 vccd1 _07499_/A sky130_fd_sc_hd__xnor2_2
X_09304_ _09304_/A _09304_/B vssd1 vssd1 vccd1 vccd1 _09304_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_63_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11153__A _12317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09235_ _09235_/A _09235_/B vssd1 vssd1 vccd1 vccd1 _09247_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_35_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_564 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09166_ _12428_/A _11973_/B _08680_/A vssd1 vssd1 vccd1 vccd1 _09166_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_121_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09097_ _09095_/X _09096_/X _09330_/S vssd1 vssd1 vccd1 vccd1 _09097_/X sky130_fd_sc_hd__mux2_1
X_08117_ _08724_/A _08117_/B vssd1 vssd1 vccd1 vccd1 _08119_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_101_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07078__A _11470_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08048_ _08752_/A _09614_/A _11908_/A vssd1 vssd1 vccd1 vccd1 _08049_/B sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout88_A _07204_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10010_ _10010_/A vssd1 vssd1 vccd1 vccd1 _10019_/A sky130_fd_sc_hd__inv_2
XANTENNA__10706__B1 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09999_ _10780_/A _09995_/X _09996_/X _09998_/Y vssd1 vssd1 vccd1 vccd1 dest_val[5]
+ sky130_fd_sc_hd__a22o_4
X_11961_ reg1_val[23] curr_PC[23] vssd1 vssd1 vccd1 vccd1 _11962_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08127__A1 _08732_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08127__B2 _10927_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09875__A1 _11294_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09875__B2 _10418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10912_ _10913_/A _10913_/B _10913_/C vssd1 vssd1 vccd1 vccd1 _11081_/A sky130_fd_sc_hd__a21o_1
X_11892_ _11450_/B _11966_/B hold225/A vssd1 vssd1 vccd1 vccd1 _11892_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_79_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10843_ _10844_/A _10844_/B _10842_/Y vssd1 vssd1 vccd1 vccd1 _10843_/X sky130_fd_sc_hd__o21ba_1
X_10774_ _10252_/S _09827_/X _09181_/X vssd1 vssd1 vccd1 vccd1 _10774_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_94_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07638__B1 _07688_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12513_ _12673_/B _12513_/B vssd1 vssd1 vccd1 vccd1 _12514_/B sky130_fd_sc_hd__or2_1
XFILLER_0_81_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07102__A2 _10570_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11998__A _12261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12444_ _12626_/A curr_PC[0] _12448_/S vssd1 vssd1 vccd1 vccd1 _12446_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_124_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08602__A2 _08741_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12375_ _12373_/A _12373_/B _12373_/C vssd1 vssd1 vccd1 vccd1 _12376_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_34_172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11002__S _12174_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11326_ _11707_/A _11326_/B _11326_/C vssd1 vssd1 vccd1 vccd1 _11326_/X sky130_fd_sc_hd__and3_1
XFILLER_0_50_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11257_ _11178_/B _11181_/B _11176_/Y vssd1 vssd1 vccd1 vccd1 _11266_/A sky130_fd_sc_hd__a21o_1
XANTENNA__09915__B _10797_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11188_ _11188_/A _11188_/B _11188_/C vssd1 vssd1 vccd1 vccd1 _11188_/X sky130_fd_sc_hd__and3_1
X_10208_ _10422_/A _10208_/B vssd1 vssd1 vccd1 vccd1 _10209_/B sky130_fd_sc_hd__xor2_1
X_10139_ curr_PC[6] _10138_/B _11142_/S vssd1 vssd1 vccd1 vccd1 _10139_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_89_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09142__S _09142_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07341__A2 _09440_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07350_ _07350_/A _07350_/B vssd1 vssd1 vccd1 vccd1 _07362_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_58_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09020_ _09014_/Y _09018_/Y _08491_/B _09021_/A vssd1 vssd1 vccd1 vccd1 _09020_/X
+ sky130_fd_sc_hd__a211o_1
X_07281_ _07281_/A _07281_/B vssd1 vssd1 vccd1 vccd1 _07294_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_5_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold202 hold202/A vssd1 vssd1 vccd1 vccd1 hold202/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11728__A2 _09527_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold224 hold224/A vssd1 vssd1 vccd1 vccd1 hold224/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold213 hold213/A vssd1 vssd1 vccd1 vccd1 hold213/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold235 hold235/A vssd1 vssd1 vccd1 vccd1 hold235/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07801__B1 _08724_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10936__B1 _10574_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold257 hold257/A vssd1 vssd1 vccd1 vccd1 hold257/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold246 hold246/A vssd1 vssd1 vccd1 vccd1 hold246/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold268 hold268/A vssd1 vssd1 vccd1 vccd1 hold268/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold279 hold279/A vssd1 vssd1 vccd1 vccd1 hold279/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10751__S _12174_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09922_ _09922_/A _09922_/B vssd1 vssd1 vccd1 vccd1 _09923_/C sky130_fd_sc_hd__xnor2_1
X_09853_ _09853_/A _09853_/B _09853_/C vssd1 vssd1 vccd1 vccd1 _09854_/B sky130_fd_sc_hd__nor3_1
XANTENNA__09554__B1 _10413_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09784_ _09598_/A _12264_/B _09604_/B _09602_/X vssd1 vssd1 vccd1 vccd1 _09786_/B
+ sky130_fd_sc_hd__a31o_1
X_08804_ _08805_/A _08805_/B vssd1 vssd1 vccd1 vccd1 _08853_/B sky130_fd_sc_hd__and2_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10052__A _11564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06996_ reg1_val[16] reg1_val[17] vssd1 vssd1 vccd1 vccd1 _06997_/C sky130_fd_sc_hd__or2_1
X_08735_ _08735_/A _08735_/B vssd1 vssd1 vccd1 vccd1 _08736_/B sky130_fd_sc_hd__xor2_2
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07064__C _07100_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08666_ _08666_/A _08666_/B vssd1 vssd1 vccd1 vccd1 _08669_/B sky130_fd_sc_hd__xor2_1
XANTENNA__07868__B1 _11558_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08597_ _07752_/B _08727_/A2 _08673_/B _12802_/A vssd1 vssd1 vccd1 vccd1 _08598_/B
+ sky130_fd_sc_hd__o22a_1
X_07617_ fanout74/X _10818_/A _10963_/A _10948_/B2 vssd1 vssd1 vccd1 vccd1 _07618_/B
+ sky130_fd_sc_hd__o22a_1
X_07548_ _09548_/A _07548_/B vssd1 vssd1 vccd1 vccd1 _07552_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_72_91 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07479_ _12840_/A _10167_/A1 _10022_/B1 _12842_/A vssd1 vssd1 vccd1 vccd1 _07480_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_64_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09218_ _10165_/A _09218_/B vssd1 vssd1 vccd1 vccd1 _09220_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_63_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10490_ _10490_/A _10490_/B vssd1 vssd1 vccd1 vccd1 _10493_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_16_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08192__A _08740_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09149_ _12626_/A curr_PC[0] vssd1 vssd1 vccd1 vccd1 _09149_/X sky130_fd_sc_hd__or2_1
XFILLER_0_44_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12160_ _12160_/A _12160_/B vssd1 vssd1 vccd1 vccd1 _12280_/A sky130_fd_sc_hd__or2_2
XANTENNA__10927__B1 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11111_ _11111_/A _11111_/B vssd1 vssd1 vccd1 vccd1 _11111_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_102_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12091_ _12093_/A _12093_/B _12093_/C vssd1 vssd1 vccd1 vccd1 _12094_/A sky130_fd_sc_hd__a21o_1
X_11042_ _11470_/A _11042_/B vssd1 vssd1 vccd1 vccd1 _11046_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__11058__A _11261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12993_ _13013_/A hold184/X vssd1 vssd1 vccd1 vccd1 _13299_/D sky130_fd_sc_hd__and2_1
XFILLER_0_98_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08367__A _10949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07859__B1 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11944_ _11944_/A _11944_/B vssd1 vssd1 vccd1 vccd1 _12165_/B sky130_fd_sc_hd__or2_2
X_11875_ _11875_/A _11875_/B vssd1 vssd1 vccd1 vccd1 _11876_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_39_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10826_ _10665_/A _10665_/B _10681_/A vssd1 vssd1 vccd1 vccd1 _10838_/A sky130_fd_sc_hd__o21bai_1
XFILLER_0_109_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10757_ _10754_/X _10756_/Y _10632_/X _10636_/X vssd1 vssd1 vccd1 vccd1 _10757_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_54_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13212__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10688_ _10689_/A _10689_/B vssd1 vssd1 vccd1 vccd1 _10835_/A sky130_fd_sc_hd__and2_1
XFILLER_0_14_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12427_ _12426_/A _12426_/B _12426_/C vssd1 vssd1 vccd1 vccd1 _12428_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_2_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08036__B1 _08656_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12358_ _06621_/A _09158_/Y _09154_/Y vssd1 vssd1 vccd1 vccd1 _12358_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_77_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09645__B _09647_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12289_ _12287_/A _12287_/B _12383_/A _12170_/A vssd1 vssd1 vccd1 vccd1 _12290_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_10_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11309_ _11310_/A _11310_/B vssd1 vssd1 vccd1 vccd1 _11417_/A sky130_fd_sc_hd__nand2_1
X_06850_ reg1_val[30] _07345_/A _06849_/X vssd1 vssd1 vccd1 vccd1 _06851_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_93_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06781_ reg1_val[4] _11233_/S vssd1 vssd1 vccd1 vccd1 _06781_/X sky130_fd_sc_hd__and2_1
XFILLER_0_89_142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08520_ _08540_/A _08540_/B vssd1 vssd1 vccd1 vccd1 _08543_/B sky130_fd_sc_hd__or2_1
XANTENNA__08277__A _08745_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07314__A2 _12808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08451_ _08451_/A _08451_/B vssd1 vssd1 vccd1 vccd1 _08487_/B sky130_fd_sc_hd__xnor2_1
X_07402_ _07600_/B _07600_/A vssd1 vssd1 vccd1 vccd1 _07402_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_85_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08382_ _08382_/A _08382_/B _08382_/C vssd1 vssd1 vccd1 vccd1 _08382_/Y sky130_fd_sc_hd__nor3_1
XFILLER_0_42_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12527__A _12686_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07333_ _07333_/A _07333_/B vssd1 vssd1 vccd1 vccd1 _07334_/B sky130_fd_sc_hd__and2_1
XFILLER_0_45_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout138_A _12812_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07264_ _12794_/A fanout16/X _07282_/B _08671_/B2 vssd1 vssd1 vccd1 vccd1 _07265_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_116_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12359__C1 _11343_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09003_ _10625_/B _10625_/C vssd1 vssd1 vccd1 vccd1 _10748_/B sky130_fd_sc_hd__and2_1
XANTENNA__13020__B1 _13213_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07195_ _09567_/B _12838_/A _09568_/B _12840_/A vssd1 vssd1 vccd1 vccd1 _07196_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout305_A _07149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08740__A _08740_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07250__B2 _10022_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07250__A1 _12832_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire3 wire3/A vssd1 vssd1 vccd1 vccd1 wire3/X sky130_fd_sc_hd__buf_1
XANTENNA__10137__A1 _11876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09905_ fanout75/X _11847_/A _11923_/A _08304_/B vssd1 vssd1 vccd1 vccd1 _09906_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_67_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09836_ _09835_/B _10124_/C hold291/A vssd1 vssd1 vccd1 vccd1 _09837_/C sky130_fd_sc_hd__a21oi_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08750__A1 _07752_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13087__B1 _07504_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09767_ _09594_/A _09594_/B _09592_/X vssd1 vssd1 vccd1 vccd1 _09771_/A sky130_fd_sc_hd__o21a_1
X_06979_ reg1_val[15] _06979_/B vssd1 vssd1 vccd1 vccd1 _09906_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__08750__B2 _07955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09698_ _09152_/Y _09672_/X _12299_/B _09111_/S _09697_/X vssd1 vssd1 vccd1 vccd1
+ _09699_/D sky130_fd_sc_hd__a221o_1
X_08718_ _08341_/Y _08719_/B _08295_/Y vssd1 vssd1 vccd1 vccd1 _08718_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08502__A1 _09423_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08649_ _08652_/A _08643_/B _08643_/C vssd1 vssd1 vccd1 vccd1 _08650_/C sky130_fd_sc_hd__a21o_1
XANTENNA__08502__B2 _12802_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11660_ _11751_/A _12261_/A vssd1 vssd1 vccd1 vccd1 _11661_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_64_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11591_ _11591_/A _11591_/B vssd1 vssd1 vccd1 vccd1 _11594_/A sky130_fd_sc_hd__xnor2_1
X_10611_ _10611_/A _10611_/B vssd1 vssd1 vccd1 vccd1 _10612_/B sky130_fd_sc_hd__xor2_2
XANTENNA__12062__B2 _12150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12062__A1 _12213_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13330_ _13340_/CLK _13330_/D vssd1 vssd1 vccd1 vccd1 hold76/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10542_ _10542_/A _10542_/B vssd1 vssd1 vccd1 vccd1 _10543_/B sky130_fd_sc_hd__and2_1
X_13261_ _13357_/CLK hold34/X vssd1 vssd1 vccd1 vccd1 hold33/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12365__A2 _07508_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12212_ _12212_/A _12212_/B vssd1 vssd1 vccd1 vccd1 _12219_/A sky130_fd_sc_hd__xnor2_1
X_10473_ _10474_/A _10474_/B _10474_/C vssd1 vssd1 vccd1 vccd1 _10603_/B sky130_fd_sc_hd__a21oi_2
X_13192_ _13214_/A hold253/X vssd1 vssd1 vccd1 vccd1 _13368_/D sky130_fd_sc_hd__and2_1
XFILLER_0_32_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11573__B1 _12213_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12172__A _12290_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12143_ _12217_/A _12143_/B vssd1 vssd1 vccd1 vccd1 _12145_/C sky130_fd_sc_hd__or2_1
XFILLER_0_20_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12074_ _12145_/A _12074_/B vssd1 vssd1 vccd1 vccd1 _12078_/A sky130_fd_sc_hd__nor2_1
X_11025_ _11015_/Y _11016_/X _11024_/Y _10113_/A _11023_/X vssd1 vssd1 vccd1 vccd1
+ _11025_/X sky130_fd_sc_hd__o221a_1
XANTENNA__08741__A1 _12820_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06752__B1 _06751_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08741__B2 _08741_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12976_ _13290_/Q _13016_/A2 _13006_/B1 hold220/X vssd1 vssd1 vccd1 vccd1 hold221/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11927_ _11927_/A _11927_/B vssd1 vssd1 vccd1 vccd1 _11928_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_74_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11858_ _11859_/B _11859_/A vssd1 vssd1 vccd1 vccd1 _11943_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_27_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_19 reg1_val[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11789_ _12098_/A _11789_/B vssd1 vssd1 vccd1 vccd1 _11822_/B sky130_fd_sc_hd__xnor2_2
X_10809_ _10810_/A _10810_/B vssd1 vssd1 vccd1 vccd1 _10809_/X sky130_fd_sc_hd__and2_1
XFILLER_0_27_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10064__B1 _10963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11013__C1 _09172_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09221__A2 _10167_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07176__A _10448_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07951_ _08724_/A _07951_/B vssd1 vssd1 vccd1 vccd1 _08033_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_120_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06902_ instruction[15] _06902_/B vssd1 vssd1 vccd1 vccd1 dest_idx[4] sky130_fd_sc_hd__and2_4
XFILLER_0_10_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12810__A _12810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07882_ _08432_/B fanout99/X _08436_/A _10537_/A1 vssd1 vssd1 vccd1 vccd1 _07883_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_128_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06833_ _06828_/Y _06832_/X _11959_/A vssd1 vssd1 vccd1 vccd1 _06833_/Y sky130_fd_sc_hd__a21oi_1
X_09621_ _10422_/A _09621_/B vssd1 vssd1 vccd1 vccd1 _09622_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__07535__A2 _07033_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08732__B2 _10927_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08732__A1 _08732_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06764_ _06805_/A _06702_/A _12659_/B _06763_/X vssd1 vssd1 vccd1 vccd1 _07036_/A
+ sky130_fd_sc_hd__a31o_4
X_09552_ _09552_/A _09552_/B vssd1 vssd1 vccd1 vccd1 _09553_/B sky130_fd_sc_hd__nand2_1
XANTENNA__10330__A _11180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08503_ _09433_/A _08503_/B vssd1 vssd1 vccd1 vccd1 _08521_/B sky130_fd_sc_hd__xnor2_1
X_06695_ _06695_/A _12634_/B vssd1 vssd1 vccd1 vccd1 _06695_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__08496__B1 _08656_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09483_ _09484_/A _09484_/B vssd1 vssd1 vccd1 vccd1 _09483_/X sky130_fd_sc_hd__and2_1
X_08434_ _08434_/A _08434_/B vssd1 vssd1 vccd1 vccd1 _08449_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_19_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08365_ _08363_/Y _08416_/B _08360_/Y vssd1 vssd1 vccd1 vccd1 _08387_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_46_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07316_ _07317_/A _07317_/B vssd1 vssd1 vccd1 vccd1 _07573_/A sky130_fd_sc_hd__and2_1
XFILLER_0_34_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08296_ _08296_/A _08296_/B vssd1 vssd1 vccd1 vccd1 _08297_/B sky130_fd_sc_hd__or2_1
XFILLER_0_104_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07247_ _09431_/A _07247_/B vssd1 vssd1 vccd1 vccd1 _07249_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_61_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07178_ _11020_/A _07178_/B vssd1 vssd1 vccd1 vccd1 _07178_/Y sky130_fd_sc_hd__xnor2_4
XANTENNA__09748__B1 _11766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06702__B _12629_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout70_A _07819_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09819_ _06870_/C _09817_/X _09818_/Y vssd1 vssd1 vccd1 vccd1 _09819_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__09505__S _09505_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08723__B2 _08304_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08723__A1 fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12830_ _12830_/A _12830_/B vssd1 vssd1 vccd1 vccd1 _12830_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__10530__A1 _06924_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12761_ _12761_/A _12766_/C vssd1 vssd1 vccd1 vccd1 loadstore_address[27] sky130_fd_sc_hd__xnor2_4
XTAP_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11712_ _06676_/C _11711_/X _09156_/Y vssd1 vssd1 vccd1 vccd1 _11712_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__08645__A _08645_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12692_ reg1_val[13] _12692_/B vssd1 vssd1 vccd1 vccd1 _12701_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_127_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11643_ _11968_/B1 _11633_/X _11634_/Y _11642_/X vssd1 vssd1 vccd1 vccd1 _11644_/A
+ sky130_fd_sc_hd__o31ai_1
XFILLER_0_84_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11574_ _12073_/A _11574_/B vssd1 vssd1 vccd1 vccd1 _11575_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_24_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13313_ _13314_/CLK hold217/X vssd1 vssd1 vccd1 vccd1 hold215/A sky130_fd_sc_hd__dfxtp_1
X_10525_ _07095_/A _12404_/A _11973_/B _06750_/B _06881_/X vssd1 vssd1 vccd1 vccd1
+ _10525_/Y sky130_fd_sc_hd__a221oi_1
XFILLER_0_91_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13244_ hold299/A hold297/A hold63/X hold101/X vssd1 vssd1 vccd1 vccd1 hold102/A
+ sky130_fd_sc_hd__a31o_1
X_10456_ _10455_/B _10455_/C _10455_/A vssd1 vssd1 vccd1 vccd1 _10457_/B sky130_fd_sc_hd__a21oi_1
X_13175_ _13175_/A _13175_/B vssd1 vssd1 vccd1 vccd1 _13175_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_122_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10387_ _10252_/S _10245_/X _10386_/X vssd1 vssd1 vccd1 vccd1 _10387_/Y sky130_fd_sc_hd__a21oi_2
X_12126_ _12402_/A0 _09354_/B _12126_/S vssd1 vssd1 vccd1 vccd1 _12126_/X sky130_fd_sc_hd__mux2_1
XANTENNA__06612__B _06612_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07765__A2 fanout99/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12057_ curr_PC[24] _12058_/B vssd1 vssd1 vccd1 vccd1 _12057_/X sky130_fd_sc_hd__or2_1
X_11008_ reg1_val[12] curr_PC[12] _10888_/B vssd1 vssd1 vccd1 vccd1 _11009_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_74_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12959_ _13233_/B _12959_/B vssd1 vssd1 vccd1 vccd1 fanout2/A sky130_fd_sc_hd__or2_2
XFILLER_0_90_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08150_ _08150_/A _08150_/B vssd1 vssd1 vccd1 vccd1 _08161_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__10037__B1 _10818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07101_ _11385_/A _11470_/B vssd1 vssd1 vccd1 vccd1 _09745_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_28_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08081_ _08081_/A _08081_/B vssd1 vssd1 vccd1 vccd1 _08900_/B sky130_fd_sc_hd__xnor2_1
X_07032_ _10422_/A _07037_/B _07524_/A vssd1 vssd1 vccd1 vccd1 _07033_/B sky130_fd_sc_hd__or3b_4
XFILLER_0_3_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06803__A _09343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08983_ _08983_/A _08983_/B vssd1 vssd1 vccd1 vccd1 _08984_/B sky130_fd_sc_hd__or2_1
XANTENNA__12540__A _12698_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07934_ _08733_/A _07934_/B vssd1 vssd1 vccd1 vccd1 _07938_/B sky130_fd_sc_hd__xnor2_4
X_07865_ _07912_/B vssd1 vssd1 vccd1 vccd1 _07865_/Y sky130_fd_sc_hd__inv_2
X_09604_ _09604_/A _09604_/B vssd1 vssd1 vccd1 vccd1 _09606_/B sky130_fd_sc_hd__xnor2_2
X_06816_ _10378_/A _06815_/X _06753_/X vssd1 vssd1 vccd1 vccd1 _06816_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_97_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07796_ _12820_/A fanout87/X fanout82/X _08741_/B2 vssd1 vssd1 vccd1 vccd1 _07797_/B
+ sky130_fd_sc_hd__o22a_1
X_06747_ reg1_val[9] _07095_/A vssd1 vssd1 vccd1 vccd1 _06750_/A sky130_fd_sc_hd__nor2_1
X_09535_ _09684_/B _12403_/A1 _09354_/B _06798_/B _09531_/X vssd1 vssd1 vccd1 vccd1
+ _09535_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_93_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06678_ _06695_/A _12644_/B vssd1 vssd1 vccd1 vccd1 _06678_/Y sky130_fd_sc_hd__nor2_1
X_09466_ _09466_/A _09466_/B vssd1 vssd1 vccd1 vccd1 _09467_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_66_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08417_ _08456_/A _08456_/B vssd1 vssd1 vccd1 vccd1 _08417_/X sky130_fd_sc_hd__and2b_1
XANTENNA__07692__A1 _08671_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_532 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07692__B2 _07821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09397_ _09746_/A _09397_/B _09397_/C vssd1 vssd1 vccd1 vccd1 _09404_/A sky130_fd_sc_hd__and3_1
XFILLER_0_34_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11225__C1 _09156_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08348_ _08379_/A _08379_/B vssd1 vssd1 vccd1 vccd1 _08382_/A sky130_fd_sc_hd__nor2_1
XANTENNA__08641__B1 _09440_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08279_ _08275_/A _08275_/B _08278_/Y vssd1 vssd1 vccd1 vccd1 _08301_/A sky130_fd_sc_hd__o21ai_2
X_10310_ _12810_/A _12316_/B vssd1 vssd1 vccd1 vccd1 _10312_/B sky130_fd_sc_hd__or2_1
X_11290_ _12261_/A _11290_/B vssd1 vssd1 vccd1 vccd1 _11292_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_22_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10241_ _06767_/X _10107_/Y _06769_/B vssd1 vssd1 vccd1 vccd1 _10241_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__11528__B1 _11624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07747__A2 _11989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10172_ _10172_/A _10172_/B _10172_/C vssd1 vssd1 vccd1 vccd1 _10174_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_28_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12450__A _12629_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout183 _07016_/Y vssd1 vssd1 vccd1 vccd1 _12798_/A sky130_fd_sc_hd__clkbuf_8
Xfanout172 _07167_/Y vssd1 vssd1 vccd1 vccd1 _09440_/B1 sky130_fd_sc_hd__buf_8
Xfanout161 _08979_/X vssd1 vssd1 vccd1 vccd1 _09653_/A sky130_fd_sc_hd__buf_4
Xfanout150 _09906_/A vssd1 vssd1 vccd1 vccd1 _08724_/A sky130_fd_sc_hd__buf_12
Xfanout194 _09433_/A vssd1 vssd1 vccd1 vccd1 _10165_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_0_69_410 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07380__B1 _10571_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07263__B _07263_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12813_ hold7/X _12856_/B _12812_/Y _13128_/A vssd1 vssd1 vccd1 vccd1 hold8/A sky130_fd_sc_hd__o211a_1
XANTENNA__12256__A1 _06924_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12744_ reg1_val[24] _12782_/A vssd1 vssd1 vccd1 vccd1 _12750_/A sky130_fd_sc_hd__nand2_1
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06604__A_N _07144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12675_ _12671_/A _12675_/B vssd1 vssd1 vccd1 vccd1 _12677_/C sky130_fd_sc_hd__nand2b_1
X_11626_ reg1_val[19] curr_PC[19] vssd1 vssd1 vccd1 vccd1 _11627_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_65_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07435__B2 _12840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07435__A1 _12838_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09918__B _12316_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11557_ _11557_/A _11557_/B vssd1 vssd1 vccd1 vccd1 _11558_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10508_ _10507_/A _10507_/B _10507_/Y _11624_/A vssd1 vssd1 vccd1 vccd1 _10508_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_80_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12625__A _12626_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11488_ _11488_/A _11488_/B vssd1 vssd1 vccd1 vccd1 _11489_/B sky130_fd_sc_hd__xor2_1
X_13227_ hold268/X _12789_/B _13226_/X _12790_/A vssd1 vssd1 vccd1 vccd1 _13228_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10439_ _10439_/A _10439_/B vssd1 vssd1 vccd1 vccd1 _10440_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_20_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10145__A _10959_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13158_ _13242_/A hold280/X vssd1 vssd1 vccd1 vccd1 _13361_/D sky130_fd_sc_hd__and2_1
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13089_ hold59/X fanout1/X hold70/X vssd1 vssd1 vccd1 vccd1 _13089_/X sky130_fd_sc_hd__a21o_1
X_12109_ _06854_/X _12108_/X _12174_/S vssd1 vssd1 vccd1 vccd1 _12110_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_85_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08163__A2 fanout69/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07650_ _07149_/A _12214_/A _08436_/B _12067_/A vssd1 vssd1 vccd1 vccd1 _07651_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_18_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06601_ _06635_/A _12686_/B vssd1 vssd1 vccd1 vccd1 _06601_/Y sky130_fd_sc_hd__nor2_1
X_07581_ _07581_/A _07581_/B vssd1 vssd1 vccd1 vccd1 _07599_/A sky130_fd_sc_hd__xnor2_4
X_09320_ _09318_/X _09319_/X _09663_/S vssd1 vssd1 vccd1 vccd1 _09320_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_88_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09251_ _09251_/A _12264_/B vssd1 vssd1 vccd1 vccd1 _09257_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_75_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08202_ _11564_/A _08162_/Y _08167_/A vssd1 vssd1 vccd1 vccd1 _08208_/A sky130_fd_sc_hd__o21ai_2
X_09182_ _09182_/A _09182_/B vssd1 vssd1 vccd1 vccd1 _12430_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_8_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout120_A _12828_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08133_ _11385_/A _08133_/B vssd1 vssd1 vccd1 vccd1 _08135_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_16_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08064_ fanout75/X _08723_/B1 _07885_/B _08304_/B vssd1 vssd1 vccd1 vccd1 _08065_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_114_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07015_ _09666_/S _09351_/B _12341_/A _07064_/B vssd1 vssd1 vccd1 vccd1 _07016_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_101_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08966_ _09072_/B vssd1 vssd1 vccd1 vccd1 _09485_/B sky130_fd_sc_hd__inv_2
X_08897_ _08898_/A _08898_/B _08898_/C vssd1 vssd1 vccd1 vccd1 _08897_/X sky130_fd_sc_hd__a21o_1
X_07917_ _07916_/B _07916_/C _07916_/A vssd1 vssd1 vccd1 vccd1 _07964_/A sky130_fd_sc_hd__o21ba_1
XANTENNA__11289__A2 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07848_ _07807_/A _07806_/C _07806_/B vssd1 vssd1 vccd1 vccd1 _07848_/X sky130_fd_sc_hd__a21o_1
X_09518_ _11886_/A _09518_/B vssd1 vssd1 vccd1 vccd1 _09518_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_79_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07779_ _07811_/A _07811_/B vssd1 vssd1 vccd1 vccd1 _07781_/C sky130_fd_sc_hd__nand2_1
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12429__B _12429_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07114__B1 _11171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout33_A _12261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10790_ _10571_/A _12150_/A _12067_/A _10570_/A vssd1 vssd1 vccd1 vccd1 _10791_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11997__B1 fanout4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09449_ _10418_/A fanout69/X _08216_/B _09745_/B vssd1 vssd1 vccd1 vccd1 _09450_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_93_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12460_ _12460_/A _12460_/B _12460_/C vssd1 vssd1 vccd1 vccd1 _12461_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_47_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12391_ _09077_/A _09077_/B _12426_/A vssd1 vssd1 vccd1 vccd1 _12392_/B sky130_fd_sc_hd__a21o_1
XANTENNA__12410__A1 _06612_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11411_ _11412_/A _11412_/B vssd1 vssd1 vccd1 vccd1 _11508_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_105_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11342_ _06705_/X _09527_/B _12307_/B1 vssd1 vssd1 vccd1 vccd1 _11342_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__12445__A _12626_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10421__B1 _10930_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11987__C fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11273_ _11272_/B _11272_/C _11272_/A vssd1 vssd1 vccd1 vccd1 _11274_/B sky130_fd_sc_hd__o21a_1
X_13012_ hold207/A _13016_/A2 _13016_/B1 hold180/X vssd1 vssd1 vccd1 vccd1 hold181/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09754__A _11470_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10224_ _10224_/A _10224_/B vssd1 vssd1 vccd1 vccd1 _10225_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_30_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09590__A1 _09238_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10155_ _10155_/A _10155_/B vssd1 vssd1 vccd1 vccd1 _10159_/A sky130_fd_sc_hd__xor2_1
XANTENNA__11921__B1 fanout4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07274__A _07485_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold6 hold6/A vssd1 vssd1 vccd1 vccd1 hold6/X sky130_fd_sc_hd__dlygate4sd3_1
X_10086_ _10086_/A _10086_/B vssd1 vssd1 vccd1 vccd1 _10088_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__07353__B1 _07178_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09893__A2 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11524__A _12174_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10988_ _10988_/A _10988_/B vssd1 vssd1 vccd1 vccd1 _11100_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_29_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12727_ _12728_/B _12728_/C _12746_/A vssd1 vssd1 vccd1 vccd1 _12729_/A sky130_fd_sc_hd__a21oi_4
XFILLER_0_127_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12658_ reg1_val[7] _12659_/B vssd1 vssd1 vccd1 vccd1 _12658_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_115_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11609_ _11609_/A vssd1 vssd1 vccd1 vccd1 _11609_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_111_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12589_ _12595_/B _12589_/B vssd1 vssd1 vccd1 vccd1 new_PC[21] sky130_fd_sc_hd__xnor2_4
XFILLER_0_53_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12802__B _12818_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09581__A1 _10941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08820_ _08762_/B _08767_/B _08760_/Y vssd1 vssd1 vccd1 vccd1 _08831_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_0_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09581__B2 fanout94/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08751_ _11385_/A _08751_/B vssd1 vssd1 vccd1 vccd1 _08754_/B sky130_fd_sc_hd__xnor2_1
X_08682_ _08983_/A _08983_/B vssd1 vssd1 vccd1 vccd1 _08984_/A sky130_fd_sc_hd__nand2_1
X_07702_ _07794_/A _07794_/B vssd1 vssd1 vccd1 vccd1 _07808_/A sky130_fd_sc_hd__or2_2
XANTENNA__08136__A2 _09609_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07344__B1 _07220_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07633_ _07633_/A _07633_/B vssd1 vssd1 vccd1 vccd1 _08919_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_45_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07895__A1 _07099_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07564_ _07564_/A _07564_/B vssd1 vssd1 vccd1 vccd1 _07566_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_48_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07495_ _12848_/A _09238_/B _09440_/B1 _10941_/B vssd1 vssd1 vccd1 vccd1 _07496_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_75_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09303_ _08971_/A _08971_/B _07685_/A _07685_/B vssd1 vssd1 vccd1 vccd1 _09304_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_48_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09234_ _09906_/A _09234_/B vssd1 vssd1 vccd1 vccd1 _09235_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_35_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09165_ _09165_/A instruction[6] instruction[5] vssd1 vssd1 vccd1 vccd1 _09165_/X
+ sky130_fd_sc_hd__or3b_2
XFILLER_0_8_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08116_ _08304_/B _07896_/A _07955_/A fanout75/X vssd1 vssd1 vccd1 vccd1 _08117_/B
+ sky130_fd_sc_hd__o22a_1
X_09096_ reg1_val[4] reg1_val[27] _09108_/S vssd1 vssd1 vccd1 vccd1 _09096_/X sky130_fd_sc_hd__mux2_1
XANTENNA__07359__A _11163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08047_ _08046_/A _08811_/A _08752_/A _09614_/A vssd1 vssd1 vccd1 vccd1 _08844_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_101_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10706__A1 _10445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10706__B2 _10706_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09998_ _10780_/A _10138_/B vssd1 vssd1 vccd1 vccd1 _09998_/Y sky130_fd_sc_hd__nor2_1
X_08949_ _08950_/A _08950_/B vssd1 vssd1 vccd1 vccd1 _08949_/X sky130_fd_sc_hd__and2_1
X_11960_ reg1_val[23] curr_PC[23] vssd1 vssd1 vccd1 vccd1 _11962_/A sky130_fd_sc_hd__or2_1
XANTENNA__08127__A2 _08727_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11131__A1 _12307_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07335__B1 _12836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09875__A2 _07087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07822__A _11908_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10911_ _10813_/A _10813_/B _10809_/X vssd1 vssd1 vccd1 vccd1 _10916_/A sky130_fd_sc_hd__a21oi_1
X_11891_ hold236/A _11891_/B vssd1 vssd1 vccd1 vccd1 _11966_/B sky130_fd_sc_hd__or2_1
XFILLER_0_128_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10842_ _10701_/A _10701_/B _10699_/X vssd1 vssd1 vccd1 vccd1 _10842_/Y sky130_fd_sc_hd__a21oi_1
X_10773_ _10765_/Y _10766_/X _10768_/X _10772_/X vssd1 vssd1 vccd1 vccd1 _10773_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_109_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07638__A1 _12794_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07638__B2 _08671_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10259__A2_N _12404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12512_ _12673_/B _12513_/B vssd1 vssd1 vccd1 vccd1 _12523_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_66_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09749__A _11163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12443_ _07064_/B _06939_/Y _12421_/X _12442_/Y _12455_/S vssd1 vssd1 vccd1 vccd1
+ dest_val[31] sky130_fd_sc_hd__o221a_4
XFILLER_0_50_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12374_ _12374_/A vssd1 vssd1 vccd1 vccd1 _12376_/A sky130_fd_sc_hd__inv_2
XFILLER_0_1_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11325_ _11792_/A _11360_/A _11649_/A vssd1 vssd1 vccd1 vccd1 _11326_/C sky130_fd_sc_hd__or3_1
X_11256_ _11034_/B _11650_/B _11650_/C vssd1 vssd1 vccd1 vccd1 _11360_/A sky130_fd_sc_hd__and3b_1
XFILLER_0_50_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_49 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11187_ _11187_/A _11187_/B vssd1 vssd1 vccd1 vccd1 _11188_/C sky130_fd_sc_hd__or2_1
X_10207_ _07087_/X _11472_/A _10574_/B fanout66/X vssd1 vssd1 vccd1 vccd1 _10208_/B
+ sky130_fd_sc_hd__o22a_1
X_10138_ curr_PC[6] _10138_/B vssd1 vssd1 vccd1 vccd1 _10403_/C sky130_fd_sc_hd__and2_1
X_10069_ _10069_/A _10069_/B vssd1 vssd1 vccd1 vccd1 _10070_/B sky130_fd_sc_hd__nor2_1
XANTENNA__11122__A1 _11886_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07732__A _08740_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07280_ _09746_/A _07280_/B vssd1 vssd1 vccd1 vccd1 _07281_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_122_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08563__A _08742_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10397__C1 _10396_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold225 hold225/A vssd1 vssd1 vccd1 vccd1 hold225/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold203 hold203/A vssd1 vssd1 vccd1 vccd1 hold203/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold214 hold214/A vssd1 vssd1 vccd1 vccd1 hold214/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07801__A1 _07800_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10936__B2 fanout27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10936__A1 fanout30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold236 hold236/A vssd1 vssd1 vccd1 vccd1 hold236/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold247 hold247/A vssd1 vssd1 vccd1 vccd1 hold247/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold269 hold269/A vssd1 vssd1 vccd1 vccd1 hold269/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold258 hold258/A vssd1 vssd1 vccd1 vccd1 hold258/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09921_ _09922_/A _09922_/B vssd1 vssd1 vccd1 vccd1 _10056_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_1_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09554__A1 fanout30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09554__B2 _07688_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09852_ _11142_/S _09850_/Y _09851_/X _09849_/Y vssd1 vssd1 vccd1 vccd1 dest_val[4]
+ sky130_fd_sc_hd__a31o_4
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09783_ _09912_/A _09783_/B vssd1 vssd1 vccd1 vccd1 _09786_/A sky130_fd_sc_hd__and2_1
X_08803_ _11564_/A _08803_/B vssd1 vssd1 vccd1 vccd1 _08805_/B sky130_fd_sc_hd__xnor2_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout285_A _06587_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06995_ reg1_val[20] reg1_val[21] reg1_val[22] vssd1 vssd1 vccd1 vccd1 _06998_/B
+ sky130_fd_sc_hd__or3_1
X_08734_ _08735_/A _08735_/B vssd1 vssd1 vccd1 vccd1 _08734_/Y sky130_fd_sc_hd__nor2_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08665_ _08683_/A _08683_/B vssd1 vssd1 vccd1 vccd1 _08667_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_49_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07868__A1 _08732_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07868__B2 _08656_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08596_ _08645_/A _08596_/B vssd1 vssd1 vccd1 vccd1 _08627_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__10872__B1 _11707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07616_ _10710_/A _07616_/B vssd1 vssd1 vccd1 vccd1 _07621_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__11164__A _11164_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07547_ _12798_/A fanout16/X _07282_/B _09423_/B2 vssd1 vssd1 vccd1 vccd1 _07548_/B
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_118_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07478_ _07478_/A _07478_/B vssd1 vssd1 vccd1 vccd1 _07481_/A sky130_fd_sc_hd__nor2_1
XANTENNA__09490__B1 _11707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08473__A _10444_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09217_ _12846_/A _09567_/B _09568_/B _12848_/A vssd1 vssd1 vccd1 vccd1 _09218_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_63_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07089__A _07089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09148_ _12626_/A curr_PC[0] vssd1 vssd1 vccd1 vccd1 _09345_/A sky130_fd_sc_hd__nand2_1
X_09079_ _09542_/A _09079_/B vssd1 vssd1 vccd1 vccd1 _09079_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_16_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10927__B2 _11367_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10927__A1 _10927_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11110_ _06821_/X _11109_/X _12174_/S vssd1 vssd1 vccd1 vccd1 _11111_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_32_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12090_ _12159_/B _12090_/B vssd1 vssd1 vccd1 vccd1 _12093_/C sky130_fd_sc_hd__nand2_1
XANTENNA__11352__A1 _09156_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07536__B _10567_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11041_ _10941_/A _12316_/A fanout12/X fanout94/X vssd1 vssd1 vccd1 vccd1 _11042_/B
+ sky130_fd_sc_hd__o22a_1
X_12992_ hold183/X _13004_/A2 _13006_/B1 hold174/X vssd1 vssd1 vccd1 vccd1 hold184/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08648__A _08655_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07859__A1 _12818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07859__B2 _12820_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11943_ _11943_/A _11943_/B _11943_/C vssd1 vssd1 vccd1 vccd1 _11944_/B sky130_fd_sc_hd__and3_1
XFILLER_0_52_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11874_ _11874_/A _11874_/B vssd1 vssd1 vccd1 vccd1 _11875_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_67_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10825_ _10825_/A _10825_/B vssd1 vssd1 vccd1 vccd1 _10839_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_55_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10756_ reg1_val[11] curr_PC[11] vssd1 vssd1 vccd1 vccd1 _10756_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_82_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12109__S _12174_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06834__A2 _07194_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10687_ _11180_/A _10687_/B vssd1 vssd1 vccd1 vccd1 _10689_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__10418__A _10418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06615__B _12698_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12426_ _12426_/A _12426_/B _12426_/C vssd1 vssd1 vccd1 vccd1 _12428_/B sky130_fd_sc_hd__or3_1
XANTENNA__09233__B1 _12832_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08036__A1 _10927_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08036__B2 _11367_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10379__C1 _11624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09784__A1 _09598_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12357_ _13312_/Q _12434_/B1 _12399_/B _12401_/B1 vssd1 vssd1 vccd1 vccd1 _12357_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_23_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12288_ _12170_/A _12287_/X _12383_/A vssd1 vssd1 vccd1 vccd1 _12290_/B sky130_fd_sc_hd__a21oi_1
X_11308_ _11308_/A _11308_/B vssd1 vssd1 vccd1 vccd1 _11310_/B sky130_fd_sc_hd__xnor2_1
X_11239_ _08980_/Y _11237_/Y _11238_/X _09169_/Y vssd1 vssd1 vccd1 vccd1 _11249_/A
+ sky130_fd_sc_hd__o211a_1
XANTENNA__10153__A _11172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07547__B1 _07282_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06780_ _06805_/A _06686_/A _12649_/B _06778_/X vssd1 vssd1 vccd1 vccd1 _07050_/A
+ sky130_fd_sc_hd__a31oi_4
XFILLER_0_89_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08450_ _08457_/A _08457_/B _08435_/Y vssd1 vssd1 vccd1 vccd1 _08487_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07401_ _07401_/A _07401_/B vssd1 vssd1 vccd1 vccd1 _07600_/B sky130_fd_sc_hd__xnor2_2
X_08381_ _08381_/A _08381_/B vssd1 vssd1 vccd1 vccd1 _08382_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__12808__A _12808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07332_ _07333_/A _07333_/B vssd1 vssd1 vccd1 vccd1 _07334_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_73_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07263_ _12076_/A _07263_/B vssd1 vssd1 vccd1 vccd1 _07263_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_0_45_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07194_ _07194_/A _07194_/B vssd1 vssd1 vccd1 vccd1 _07194_/X sky130_fd_sc_hd__xor2_1
X_09002_ _09002_/A _09002_/B vssd1 vssd1 vccd1 vccd1 _10625_/C sky130_fd_sc_hd__xor2_2
XFILLER_0_14_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_493 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09328__S _09669_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07250__A2 _10167_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09904_ _10710_/A _09904_/B vssd1 vssd1 vccd1 vccd1 _09908_/A sky130_fd_sc_hd__xnor2_1
X_09835_ hold291/A _09835_/B _10124_/C vssd1 vssd1 vccd1 vccd1 _09837_/B sky130_fd_sc_hd__and3_1
XANTENNA__07538__B1 _11987_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13087__B2 _13087_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09766_ _09766_/A _12316_/B vssd1 vssd1 vccd1 vccd1 _09772_/A sky130_fd_sc_hd__or2_1
X_06978_ reg1_val[15] _06979_/B vssd1 vssd1 vccd1 vccd1 _11164_/A sky130_fd_sc_hd__xor2_4
XANTENNA__08750__A2 fanout69/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09697_ _09156_/Y _09686_/Y _09687_/Y _09696_/Y vssd1 vssd1 vccd1 vccd1 _09697_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_68_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08717_ _08295_/B _08295_/C _08295_/A vssd1 vssd1 vccd1 vccd1 _08719_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_95_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08648_ _08655_/A _08655_/B vssd1 vssd1 vccd1 vccd1 _08650_/B sky130_fd_sc_hd__nor2_1
XANTENNA__08502__A2 _08741_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_327 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11325__C _11649_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08579_ _12802_/A _08661_/A2 _08673_/B _12804_/A vssd1 vssd1 vccd1 vccd1 _08580_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_76_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11590_ _11591_/A _11591_/B vssd1 vssd1 vccd1 vccd1 _11687_/B sky130_fd_sc_hd__nand2_1
X_10610_ _10611_/A _10611_/B vssd1 vssd1 vccd1 vccd1 _10610_/X sky130_fd_sc_hd__or2_1
XANTENNA__12062__A2 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11270__B1 _11470_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10541_ _10542_/A _10542_/B vssd1 vssd1 vccd1 vccd1 _10543_/A sky130_fd_sc_hd__nor2_1
X_13260_ _13357_/CLK hold8/X vssd1 vssd1 vccd1 vccd1 hold7/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09215__B1 _08507_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12211_ _12212_/A _12212_/B vssd1 vssd1 vccd1 vccd1 _12211_/X sky130_fd_sc_hd__and2b_1
X_10472_ _10603_/A _10472_/B vssd1 vssd1 vccd1 vccd1 _10474_/C sky130_fd_sc_hd__or2_1
X_13191_ hold252/X _13213_/A2 _13190_/X _13213_/B2 vssd1 vssd1 vccd1 vccd1 hold253/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07777__B1 _09396_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12365__A3 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11573__A1 fanout24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12142_ _12142_/A _12142_/B vssd1 vssd1 vccd1 vccd1 _12143_/B sky130_fd_sc_hd__and2_1
XANTENNA__11573__B2 _07819_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12073_ _12073_/A _12073_/B vssd1 vssd1 vccd1 vccd1 _12074_/B sky130_fd_sc_hd__and2_1
XFILLER_0_20_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11024_ _10119_/S _09510_/X _09181_/X vssd1 vssd1 vccd1 vccd1 _11024_/Y sky130_fd_sc_hd__o21ai_2
XANTENNA__08741__A2 _08741_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12975_ _13009_/A hold158/X vssd1 vssd1 vccd1 vccd1 hold159/A sky130_fd_sc_hd__and2_1
XFILLER_0_99_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07282__A _12794_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_2_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13378_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_87_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11926_ _11927_/A _11927_/B vssd1 vssd1 vccd1 vccd1 _11926_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_86_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11857_ _11943_/A _11857_/B vssd1 vssd1 vccd1 vccd1 _11859_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_103_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09454__B1 _10575_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11788_ _11427_/B _11787_/Y _12099_/A vssd1 vssd1 vccd1 vccd1 _11789_/B sky130_fd_sc_hd__a21oi_1
X_10808_ _12210_/A _10808_/B vssd1 vssd1 vccd1 vccd1 _10810_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10739_ _10739_/A _11102_/A vssd1 vssd1 vccd1 vccd1 _10992_/A sky130_fd_sc_hd__or2_1
XANTENNA__10064__A1 _11065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10064__B2 fanout24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10148__A _10148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13389_ instruction[15] vssd1 vssd1 vccd1 vccd1 loadstore_dest[4] sky130_fd_sc_hd__buf_12
XFILLER_0_88_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12409_ _12389_/Y _12390_/X _12408_/X vssd1 vssd1 vccd1 vccd1 _12409_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_11_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07950_ fanout75/X _07885_/B _08721_/B1 _08304_/B vssd1 vssd1 vccd1 vccd1 _07951_/B
+ sky130_fd_sc_hd__o22a_1
X_06901_ instruction[14] _06902_/B vssd1 vssd1 vccd1 vccd1 dest_idx[3] sky130_fd_sc_hd__and2_4
XFILLER_0_128_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08193__B1 _07752_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07881_ _07881_/A _07881_/B vssd1 vssd1 vccd1 vccd1 _07902_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_128_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13069__A1 _07037_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06832_ _06829_/Y _06831_/X _11880_/A vssd1 vssd1 vccd1 vccd1 _06832_/X sky130_fd_sc_hd__a21o_1
X_09620_ _11065_/A _11653_/A _08752_/B _11146_/A vssd1 vssd1 vccd1 vccd1 _09621_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11707__A _11707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08732__A2 _08732_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06763_ reg2_val[6] _06799_/B vssd1 vssd1 vccd1 vccd1 _06763_/X sky130_fd_sc_hd__and2_1
X_09551_ _09552_/A _09552_/B vssd1 vssd1 vccd1 vccd1 _09553_/A sky130_fd_sc_hd__or2_1
X_08502_ _09423_/B2 _08741_/A2 _08617_/B _12802_/A vssd1 vssd1 vccd1 vccd1 _08503_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_77_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10827__B1 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06694_ instruction[27] _06694_/B vssd1 vssd1 vccd1 vccd1 _12634_/B sky130_fd_sc_hd__and2_4
XANTENNA__08496__A1 _07896_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08496__B2 _08723_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09482_ _09484_/A _09484_/B vssd1 vssd1 vccd1 vccd1 _09482_/X sky130_fd_sc_hd__or2_2
XFILLER_0_93_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08433_ _08469_/A _08722_/A _08469_/B vssd1 vssd1 vccd1 vccd1 _08449_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_58_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout150_A _09906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08364_ _08364_/A _08364_/B vssd1 vssd1 vccd1 vccd1 _08416_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_46_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07315_ _11987_/A _07315_/B vssd1 vssd1 vccd1 vccd1 _07317_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_18_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08295_ _08295_/A _08295_/B _08295_/C vssd1 vssd1 vccd1 vccd1 _08295_/Y sky130_fd_sc_hd__nor3_1
XFILLER_0_6_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07246_ _12828_/A _10589_/A _12830_/A _08507_/B vssd1 vssd1 vccd1 vccd1 _07247_/B
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_5_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08751__A _11385_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07177_ _07074_/A _07074_/C _07074_/B vssd1 vssd1 vccd1 vccd1 _07178_/B sky130_fd_sc_hd__o21a_1
XANTENNA__09748__A1 _10948_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09748__B2 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07367__A _12794_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout310 instruction[7] vssd1 vssd1 vccd1 vccd1 _12341_/A sky130_fd_sc_hd__buf_8
XANTENNA__09582__A _11384_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09818_ _06870_/C _09817_/X _11624_/A vssd1 vssd1 vccd1 vccd1 _09818_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__08723__A2 _07896_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12807__A1 _07035_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09749_ _11163_/A _09749_/B vssd1 vssd1 vccd1 vccd1 _09751_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__07931__B1 _11766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12760_ reg1_val[27] _12782_/A vssd1 vssd1 vccd1 vccd1 _12766_/C sky130_fd_sc_hd__xnor2_4
XTAP_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11711_ _06827_/Y _11710_/Y _12174_/S vssd1 vssd1 vccd1 vccd1 _11711_/X sky130_fd_sc_hd__mux2_1
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12691_ reg1_val[13] _12692_/B vssd1 vssd1 vccd1 vccd1 _12693_/A sky130_fd_sc_hd__or2_1
XFILLER_0_37_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11642_ _12247_/C1 _11636_/X _11637_/Y _11641_/X vssd1 vssd1 vccd1 vccd1 _11642_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_83_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09436__B1 _10022_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13312_ _13314_/CLK hold171/X vssd1 vssd1 vccd1 vccd1 _13312_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11573_ fanout24/X _12150_/A _12213_/A _07819_/B vssd1 vssd1 vccd1 vccd1 _11574_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_9_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10524_ hold288/A _11452_/B1 _10646_/B _09837_/A vssd1 vssd1 vccd1 vccd1 _10524_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_107_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09757__A _10165_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13243_ hold101/X _06892_/B _12786_/Y _06572_/A vssd1 vssd1 vccd1 vccd1 _13245_/B
+ sky130_fd_sc_hd__a22o_1
X_10455_ _10455_/A _10455_/B _10455_/C vssd1 vssd1 vccd1 vccd1 _10457_/A sky130_fd_sc_hd__and3_1
X_13174_ _13174_/A _13174_/B vssd1 vssd1 vccd1 vccd1 _13175_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_60_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12125_ hold207/A _12434_/B1 _12191_/B _12401_/B1 vssd1 vssd1 vccd1 vccd1 _12125_/X
+ sky130_fd_sc_hd__a31o_1
X_10386_ _11231_/S _09114_/X _10385_/X _11233_/S vssd1 vssd1 vccd1 vccd1 _10386_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_102_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12056_ _11707_/A _12029_/X _12030_/Y _12055_/X vssd1 vssd1 vccd1 vccd1 _12056_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__08175__B1 _08732_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11007_ _11007_/A _11007_/B vssd1 vssd1 vccd1 vccd1 _11009_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12958_ hold86/X _12958_/B vssd1 vssd1 vccd1 vccd1 _12959_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_90_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12889_ hold43/X hold287/A vssd1 vssd1 vccd1 vccd1 _12889_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_87_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11482__B1 fanout4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11909_ fanout24/X fanout12/X fanout8/X _07819_/B vssd1 vssd1 vccd1 vccd1 _11910_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_23_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10037__B2 fanout27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10037__A1 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07100_ _07100_/A _07100_/B vssd1 vssd1 vccd1 vccd1 _12814_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_15_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08080_ _08078_/A _08078_/B _08079_/Y vssd1 vssd1 vccd1 vccd1 _08900_/A sky130_fd_sc_hd__o21ai_1
X_07031_ _07524_/A _10422_/A _07037_/B vssd1 vssd1 vccd1 vccd1 _07033_/A sky130_fd_sc_hd__nand3b_4
XFILLER_0_24_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06803__B _09666_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07187__A _09433_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08982_ _08982_/A _08982_/B vssd1 vssd1 vccd1 vccd1 _09656_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_48_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07933_ _11367_/A _08732_/A2 _08656_/B _11472_/A vssd1 vssd1 vccd1 vccd1 _07934_/B
+ sky130_fd_sc_hd__o22a_2
X_07864_ _08745_/A _07864_/B vssd1 vssd1 vccd1 vccd1 _07912_/B sky130_fd_sc_hd__xnor2_1
X_06815_ _06867_/B _06814_/Y _06759_/X vssd1 vssd1 vccd1 vccd1 _06815_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_98_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09603_ _09603_/A _09603_/B vssd1 vssd1 vccd1 vccd1 _09604_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_97_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07795_ _07808_/A _07808_/B vssd1 vssd1 vccd1 vccd1 _07809_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_3_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06746_ _07095_/A reg1_val[9] vssd1 vssd1 vccd1 vccd1 _06746_/X sky130_fd_sc_hd__and2b_1
X_09534_ _12394_/A _09512_/Y _09518_/Y _06924_/X vssd1 vssd1 vccd1 vccd1 _09534_/X
+ sky130_fd_sc_hd__a211o_1
X_06677_ instruction[29] _06694_/B vssd1 vssd1 vccd1 vccd1 _12644_/B sky130_fd_sc_hd__and2_4
XFILLER_0_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09465_ _09465_/A _09465_/B vssd1 vssd1 vccd1 vccd1 _09466_/B sky130_fd_sc_hd__nor2_1
X_08416_ _08416_/A _08416_/B vssd1 vssd1 vccd1 vccd1 _08456_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__11172__A _11172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07692__A2 fanout24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09396_ _11294_/A _09396_/B vssd1 vssd1 vccd1 vccd1 _09397_/C sky130_fd_sc_hd__or2_1
XFILLER_0_19_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08347_ _08347_/A _08347_/B vssd1 vssd1 vccd1 vccd1 _08379_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_117_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08641__B2 _08671_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08641__A1 _08673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09577__A _10449_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08278_ _08332_/B _08332_/A vssd1 vssd1 vccd1 vccd1 _08278_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_6_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07229_ _07230_/B _07230_/A vssd1 vssd1 vccd1 vccd1 _07376_/B sky130_fd_sc_hd__and2b_1
X_10240_ _09653_/A _08994_/A _08994_/B _09163_/X _10239_/Y vssd1 vssd1 vccd1 vccd1
+ _10270_/B sky130_fd_sc_hd__a311oi_1
XANTENNA__07097__A _11384_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10171_ _10172_/A _10172_/B _10172_/C vssd1 vssd1 vccd1 vccd1 _10292_/A sky130_fd_sc_hd__and3_1
Xfanout140 _07089_/Y vssd1 vssd1 vccd1 vccd1 _12810_/A sky130_fd_sc_hd__buf_8
Xfanout162 _11633_/B vssd1 vssd1 vccd1 vccd1 _11450_/B sky130_fd_sc_hd__buf_4
Xfanout173 _09236_/B2 vssd1 vssd1 vccd1 vccd1 _08727_/B1 sky130_fd_sc_hd__clkbuf_8
Xfanout195 _07183_/X vssd1 vssd1 vccd1 vccd1 _09433_/A sky130_fd_sc_hd__buf_8
Xfanout184 _08671_/B2 vssd1 vssd1 vccd1 vccd1 _08798_/B2 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07380__A1 _10664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07380__B2 _10818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12812_ _12812_/A _12856_/B vssd1 vssd1 vccd1 vccd1 _12812_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__08656__A _08673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12743_ reg1_val[24] _12782_/A vssd1 vssd1 vccd1 vccd1 _12745_/A sky130_fd_sc_hd__or2_1
XFILLER_0_84_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12674_ _12674_/A _12683_/A vssd1 vssd1 vccd1 vccd1 _12677_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_37_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11625_ reg1_val[19] curr_PC[19] vssd1 vssd1 vccd1 vccd1 _11627_/A sky130_fd_sc_hd__or2_1
XFILLER_0_71_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12964__B1 _13213_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07435__A2 _10167_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08391__A _12626_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11556_ _11557_/A _11557_/B vssd1 vssd1 vccd1 vccd1 _11682_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_4_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10507_ _10507_/A _10507_/B vssd1 vssd1 vccd1 vccd1 _10507_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_80_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12625__B _12626_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13226_ hold266/X _13225_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13226_/X sky130_fd_sc_hd__mux2_1
XANTENNA__06623__B _12692_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11487_ _11488_/A _11488_/B vssd1 vssd1 vccd1 vccd1 _11487_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_0_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10438_ _10439_/A _10439_/B vssd1 vssd1 vccd1 vccd1 _10438_/Y sky130_fd_sc_hd__nand2_1
X_13157_ hold279/X _06892_/B _13156_/X _13246_/B2 vssd1 vssd1 vccd1 vccd1 hold280/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10369_ _08977_/A _08977_/B _09706_/X _10368_/X vssd1 vssd1 vccd1 vccd1 _10369_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13088_ hold70/X hold59/X fanout1/X vssd1 vssd1 vccd1 vccd1 hold302/A sky130_fd_sc_hd__nand3_1
X_12108_ _06648_/D _12033_/Y _12049_/S vssd1 vssd1 vccd1 vccd1 _12108_/X sky130_fd_sc_hd__o21a_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12039_ reg1_val[24] curr_PC[24] vssd1 vssd1 vccd1 vccd1 _12040_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_18_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10161__A _10941_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06600_ instruction[37] _06634_/B vssd1 vssd1 vccd1 vccd1 _12686_/B sky130_fd_sc_hd__and2_4
X_07580_ _07580_/A _07580_/B vssd1 vssd1 vccd1 vccd1 _07581_/B sky130_fd_sc_hd__nor2_2
XANTENNA__11455__B1 _11454_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09250_ _09379_/A _09249_/C _09249_/A vssd1 vssd1 vccd1 vccd1 _09258_/B sky130_fd_sc_hd__a21o_1
XANTENNA__08320__B1 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08201_ _08214_/A _08214_/B _08190_/Y vssd1 vssd1 vccd1 vccd1 _08210_/A sky130_fd_sc_hd__a21o_1
XANTENNA__12816__A _12816_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09181_ _11233_/S _09181_/B vssd1 vssd1 vccd1 vccd1 _09181_/X sky130_fd_sc_hd__or2_4
XFILLER_0_62_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08132_ _07821_/A fanout69/X _08216_/B _07752_/B vssd1 vssd1 vccd1 vccd1 _08133_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_16_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08063_ _08722_/A _08063_/B vssd1 vssd1 vccd1 vccd1 _08809_/A sky130_fd_sc_hd__xnor2_2
XANTENNA_fanout113_A _08732_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07014_ _12076_/A _12139_/A _07012_/X vssd1 vssd1 vccd1 vccd1 _07014_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__10336__A _11172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10946__B1_N _10448_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08965_ _08965_/A _08965_/B vssd1 vssd1 vccd1 vccd1 _09072_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_11_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07916_ _07916_/A _07916_/B _07916_/C vssd1 vssd1 vccd1 vccd1 _08073_/A sky130_fd_sc_hd__or3_1
X_08896_ _08898_/A _08898_/B _08898_/C vssd1 vssd1 vccd1 vccd1 _08899_/A sky130_fd_sc_hd__a21oi_1
X_07847_ _07847_/A _07847_/B vssd1 vssd1 vccd1 vccd1 _07908_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__08476__A _08681_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07778_ _07833_/A _07778_/B vssd1 vssd1 vccd1 vccd1 _07811_/B sky130_fd_sc_hd__xnor2_1
X_06729_ reg1_val[12] _07074_/A vssd1 vssd1 vccd1 vccd1 _10897_/S sky130_fd_sc_hd__and2_1
XANTENNA__11446__B1 _12455_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09517_ _09517_/A _09517_/B vssd1 vssd1 vccd1 vccd1 _09518_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_39_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07114__B2 _12804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07114__A1 fanout23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11997__A1 _12150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11997__B2 _12067_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09448_ _10707_/A _09448_/B vssd1 vssd1 vccd1 vccd1 _09452_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09379_ _09379_/A _09379_/B vssd1 vssd1 vccd1 vccd1 _09393_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_53_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11630__A _12244_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12390_ _12389_/A _12389_/B _09156_/Y vssd1 vssd1 vccd1 vccd1 _12390_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_74_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11410_ _11410_/A _11410_/B vssd1 vssd1 vccd1 vccd1 _11412_/B sky130_fd_sc_hd__xnor2_2
X_11341_ hold292/A _11341_/B _11536_/C vssd1 vssd1 vccd1 vccd1 _11341_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_105_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12410__A2 _06939_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10421__A1 _07087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10421__B2 fanout66/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11272_ _11272_/A _11272_/B _11272_/C vssd1 vssd1 vccd1 vccd1 _11392_/A sky130_fd_sc_hd__nor3_2
X_13011_ _13013_/A hold208/X vssd1 vssd1 vccd1 vccd1 hold209/A sky130_fd_sc_hd__and2_1
XFILLER_0_120_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10223_ _10224_/A _10224_/B vssd1 vssd1 vccd1 vccd1 _10223_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_30_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09590__A2 _12854_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10154_ _10155_/A _10155_/B vssd1 vssd1 vccd1 vccd1 _10154_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__11921__B2 _11989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11921__A1 _12067_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold7 hold7/A vssd1 vssd1 vccd1 vccd1 hold7/X sky130_fd_sc_hd__dlygate4sd3_1
X_10085_ _10085_/A _10085_/B vssd1 vssd1 vccd1 vccd1 _10086_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_89_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07353__A1 _12822_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08550__B1 _09440_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07353__B2 fanout69/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06618__B _06838_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08302__B1 _07821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10987_ _10987_/A _10987_/B _10987_/C vssd1 vssd1 vccd1 vccd1 _10988_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_29_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11988__B2 _11172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12726_ _12741_/B _12726_/B vssd1 vssd1 vccd1 vccd1 _12728_/C sky130_fd_sc_hd__nand2_1
X_12657_ _12656_/A _12655_/A _12655_/B vssd1 vssd1 vccd1 vccd1 _12661_/A sky130_fd_sc_hd__o21ba_2
XFILLER_0_37_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11608_ _11608_/A _11787_/A vssd1 vssd1 vccd1 vccd1 _11609_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_123_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06616__B1 _06771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12588_ _12595_/A _12584_/Y _12580_/A vssd1 vssd1 vccd1 vccd1 _12589_/B sky130_fd_sc_hd__o21ai_2
XFILLER_0_80_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11539_ _11539_/A _11539_/B vssd1 vssd1 vccd1 vccd1 _11539_/X sky130_fd_sc_hd__or2_2
XFILLER_0_40_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13209_ hold261/X _13213_/A2 _13208_/X _13213_/B2 vssd1 vssd1 vccd1 vccd1 hold262/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_111_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09581__A2 _09745_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08750_ _07752_/B fanout69/X _08216_/B _07955_/A vssd1 vssd1 vccd1 vccd1 _08751_/B
+ sky130_fd_sc_hd__o22a_1
X_08681_ _08681_/A _08985_/A vssd1 vssd1 vccd1 vccd1 _08983_/B sky130_fd_sc_hd__nor2_1
X_07701_ _08728_/A _07701_/B vssd1 vssd1 vccd1 vccd1 _07794_/B sky130_fd_sc_hd__xnor2_1
X_07632_ _07292_/A _07292_/B _07293_/B vssd1 vssd1 vccd1 vccd1 _07633_/B sky130_fd_sc_hd__o21bai_1
XFILLER_0_76_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07895__A2 _07099_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11979__A1 _09156_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07563_ _07563_/A _07563_/B vssd1 vssd1 vccd1 vccd1 _07566_/A sky130_fd_sc_hd__xnor2_4
X_09302_ _09302_/A _09302_/B vssd1 vssd1 vccd1 vccd1 _09953_/A sky130_fd_sc_hd__xnor2_4
X_07494_ _09594_/A _07494_/B vssd1 vssd1 vccd1 vccd1 _07500_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_75_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout230_A _09505_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09233_ fanout74/X _12830_/A _12832_/A _10948_/B2 vssd1 vssd1 vccd1 vccd1 _09234_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_0_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13141__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_15_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13384_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_90_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09164_ instruction[4] instruction[6] instruction[5] instruction[3] vssd1 vssd1 vccd1
+ vccd1 _11973_/B sky130_fd_sc_hd__and4bb_4
XFILLER_0_44_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08115_ _08740_/A _08115_/B vssd1 vssd1 vccd1 vccd1 _08119_/A sky130_fd_sc_hd__xnor2_1
X_09095_ reg1_val[5] reg1_val[26] _09108_/S vssd1 vssd1 vccd1 vccd1 _09095_/X sky130_fd_sc_hd__mux2_1
X_08046_ _08046_/A _08046_/B _08046_/C vssd1 vssd1 vccd1 vccd1 _08811_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_102_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11903__A1 _11142_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10706__A2 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10167__B1 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09997_ curr_PC[4] curr_PC[5] _09997_/C vssd1 vssd1 vccd1 vccd1 _10138_/B sky130_fd_sc_hd__and3_1
X_08948_ _08948_/A _08948_/B vssd1 vssd1 vccd1 vccd1 _08950_/B sky130_fd_sc_hd__xnor2_2
X_08879_ _08880_/A _08880_/B vssd1 vssd1 vccd1 vccd1 _08898_/A sky130_fd_sc_hd__nand2_1
XANTENNA__11667__B1 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07335__A1 _12838_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07335__B2 _10167_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09875__A3 _07087_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10910_ _10848_/A _10848_/B _10849_/Y vssd1 vssd1 vccd1 vccd1 _10985_/A sky130_fd_sc_hd__o21ai_1
X_11890_ hold246/A _11636_/B _11970_/B _11889_/Y _12247_/C1 vssd1 vssd1 vccd1 vccd1
+ _11890_/X sky130_fd_sc_hd__a311o_1
XFILLER_0_86_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10841_ _10714_/A _10714_/B _10715_/Y vssd1 vssd1 vccd1 vccd1 _10846_/A sky130_fd_sc_hd__a21bo_1
X_10772_ _06963_/A _12404_/A _10770_/Y _10771_/X vssd1 vssd1 vccd1 vccd1 _10772_/X
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__07638__A2 fanout30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12511_ reg1_val[10] curr_PC[10] _12586_/S vssd1 vssd1 vccd1 vccd1 _12513_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_54_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12456__A _12634_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12442_ _12424_/Y _12425_/X _12441_/X vssd1 vssd1 vccd1 vccd1 _12442_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_0_66_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12395__A1 _12394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08599__B1 _09440_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12373_ _12373_/A _12373_/B _12373_/C vssd1 vssd1 vccd1 vccd1 _12374_/A sky130_fd_sc_hd__or3_1
XFILLER_0_35_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11324_ _11792_/A _11360_/A _11649_/A vssd1 vssd1 vccd1 vccd1 _11326_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_50_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11255_ _12448_/S _11251_/X _11252_/X _11254_/Y vssd1 vssd1 vccd1 vccd1 dest_val[15]
+ sky130_fd_sc_hd__a22o_4
X_10206_ _10206_/A _10206_/B vssd1 vssd1 vccd1 vccd1 _10209_/A sky130_fd_sc_hd__nor2_1
XANTENNA__11519__B _11649_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11186_ _11187_/A _11187_/B vssd1 vssd1 vccd1 vccd1 _11188_/B sky130_fd_sc_hd__nand2_1
X_10137_ _11876_/A _10106_/Y _10136_/X _10104_/Y vssd1 vssd1 vccd1 vccd1 _10137_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_89_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10068_ _10069_/A _10069_/B vssd1 vssd1 vccd1 vccd1 _10070_/A sky130_fd_sc_hd__and2_1
XANTENNA__13226__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12709_ _12709_/A _12709_/B vssd1 vssd1 vccd1 vccd1 _12712_/A sky130_fd_sc_hd__or2_2
XFILLER_0_127_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12366__A fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold215 hold215/A vssd1 vssd1 vccd1 vccd1 hold215/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold226 hold226/A vssd1 vssd1 vccd1 vccd1 hold226/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold204 hold204/A vssd1 vssd1 vccd1 vccd1 hold204/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10936__A2 _09745_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold237 hold237/A vssd1 vssd1 vccd1 vccd1 hold237/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold248 hold248/A vssd1 vssd1 vccd1 vccd1 hold248/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold259 hold259/A vssd1 vssd1 vccd1 vccd1 hold259/X sky130_fd_sc_hd__dlygate4sd3_1
X_09920_ _12138_/A _09920_/B vssd1 vssd1 vccd1 vccd1 _09922_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_1_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10614__A _10615_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09554__A2 _07089_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09851_ curr_PC[4] _09997_/C vssd1 vssd1 vccd1 vccd1 _09851_/X sky130_fd_sc_hd__or2_1
XFILLER_0_0_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09782_ _09782_/A _09782_/B vssd1 vssd1 vccd1 vccd1 _09783_/B sky130_fd_sc_hd__or2_1
X_06994_ reg1_val[13] reg1_val[14] reg1_val[15] _06994_/D vssd1 vssd1 vccd1 vccd1
+ _07254_/B sky130_fd_sc_hd__or4_4
X_08802_ _07821_/A _09609_/B _09396_/B _07752_/B vssd1 vssd1 vccd1 vccd1 _08803_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08733_ _08733_/A _08733_/B vssd1 vssd1 vccd1 vccd1 _08735_/B sky130_fd_sc_hd__xnor2_2
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13136__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout278_A _13246_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08664_ _08731_/A _08664_/B vssd1 vssd1 vccd1 vccd1 _08683_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07868__A2 _11472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08595_ _08730_/A1 _08723_/B1 _08038_/A _12804_/A vssd1 vssd1 vccd1 vccd1 _08596_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_49_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07615_ _11294_/A _10589_/A _08507_/B _10418_/A vssd1 vssd1 vccd1 vccd1 _07616_/B
+ sky130_fd_sc_hd__o22a_1
X_07546_ _07350_/A _07350_/B _07348_/Y vssd1 vssd1 vccd1 vccd1 _07552_/A sky130_fd_sc_hd__a21o_2
XFILLER_0_119_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09216_ _09431_/A _09216_/B vssd1 vssd1 vccd1 vccd1 _09220_/A sky130_fd_sc_hd__xnor2_1
X_07477_ _07477_/A _07477_/B vssd1 vssd1 vccd1 vccd1 _07478_/B sky130_fd_sc_hd__and2_1
XFILLER_0_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11180__A _11180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09147_ _09115_/X _09146_/X _09147_/S vssd1 vssd1 vccd1 vccd1 _09147_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_32_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09078_ _09653_/A _10658_/A vssd1 vssd1 vccd1 vccd1 _09079_/B sky130_fd_sc_hd__nand2_1
XANTENNA__12129__A1 _09111_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08029_ _08029_/A _08029_/B vssd1 vssd1 vccd1 vccd1 _08031_/B sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout93_A _07833_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11040_ _11040_/A _11040_/B vssd1 vssd1 vccd1 vccd1 _11048_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__09524__S _12388_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07833__A _07833_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12991_ _13013_/A hold206/X vssd1 vssd1 vccd1 vccd1 _13298_/D sky130_fd_sc_hd__and2_1
XFILLER_0_98_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07859__A2 fanout87/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11942_ _11942_/A vssd1 vssd1 vccd1 vccd1 _11944_/A sky130_fd_sc_hd__inv_2
X_11873_ _11874_/A _11872_/B _11872_/C vssd1 vssd1 vccd1 vccd1 _11873_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_39_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10824_ _10971_/B _10822_/B _10822_/C vssd1 vssd1 vccd1 vccd1 _10825_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_109_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08664__A _08731_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10755_ reg1_val[11] curr_PC[11] vssd1 vssd1 vccd1 vccd1 _10755_/X sky130_fd_sc_hd__and2_1
XFILLER_0_82_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10686_ _10574_/A _10575_/B _10930_/B _10575_/A vssd1 vssd1 vccd1 vccd1 _10687_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10418__B _11171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12425_ _08980_/B _12422_/X _12423_/Y _09157_/X vssd1 vssd1 vccd1 vccd1 _12425_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__09233__A1 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08036__A2 _08732_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12356_ _12434_/B1 _12399_/B _13312_/Q vssd1 vssd1 vccd1 vccd1 _12356_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__07244__B1 _12836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09784__A2 _12264_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09233__B2 _10948_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12633__B _12634_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11307_ _11308_/A _11308_/B vssd1 vssd1 vccd1 vccd1 _11307_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_23_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12287_ _12287_/A _12287_/B vssd1 vssd1 vccd1 vccd1 _12287_/X sky130_fd_sc_hd__or2_1
XFILLER_0_10_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11238_ _11450_/B _11346_/B hold183/A vssd1 vssd1 vccd1 vccd1 _11238_/X sky130_fd_sc_hd__a21o_1
XANTENNA__07547__A1 _12798_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07547__B2 _09423_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08744__B1 _08564_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11169_ _11292_/B _11169_/B vssd1 vssd1 vccd1 vccd1 _11187_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_93_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07400_ _08958_/A _08958_/B _07397_/Y vssd1 vssd1 vccd1 vccd1 _07600_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_58_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08380_ _08424_/A _08424_/B vssd1 vssd1 vccd1 vccd1 _08382_/B sky130_fd_sc_hd__and2_1
XFILLER_0_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07331_ _09433_/A _07331_/B vssd1 vssd1 vccd1 vccd1 _07333_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_58_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07262_ _07262_/A _07262_/B vssd1 vssd1 vccd1 vccd1 _07262_/X sky130_fd_sc_hd__or2_1
XFILLER_0_5_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07193_ _07191_/A _07220_/C _07134_/Y _07074_/B vssd1 vssd1 vccd1 vccd1 _07194_/B
+ sky130_fd_sc_hd__o31a_1
X_09001_ _10503_/B _10503_/C vssd1 vssd1 vccd1 vccd1 _10625_/B sky130_fd_sc_hd__and2_1
XANTENNA__12824__A _12824_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07235__B1 _12840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10909__A2 _10782_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10790__B1 _12067_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09903_ _12214_/A _10589_/A _08507_/B fanout59/X vssd1 vssd1 vccd1 vccd1 _09904_/B
+ sky130_fd_sc_hd__o22a_1
X_09834_ hold284/A hold240/A hold244/A hold260/A vssd1 vssd1 vccd1 vccd1 _10124_/C
+ sky130_fd_sc_hd__or4_2
XFILLER_0_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09765_ _09765_/A _09765_/B vssd1 vssd1 vccd1 vccd1 _09774_/A sky130_fd_sc_hd__xor2_1
X_06977_ reg1_val[13] reg1_val[14] _06994_/D _07364_/B1 vssd1 vssd1 vccd1 vccd1 _06979_/B
+ sky130_fd_sc_hd__o31a_4
XANTENNA__11175__A _11261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09696_ _09689_/Y _09690_/X _09695_/X vssd1 vssd1 vccd1 vccd1 _09696_/Y sky130_fd_sc_hd__o21ai_1
X_08716_ _08427_/Y _08711_/A _08711_/B _08714_/X _08713_/Y vssd1 vssd1 vccd1 vccd1
+ _09028_/B sky130_fd_sc_hd__a41o_1
XFILLER_0_96_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08647_ _08728_/A _08647_/B vssd1 vssd1 vccd1 vccd1 _08655_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_68_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08578_ _08584_/A _08584_/B vssd1 vssd1 vccd1 vccd1 _08578_/X sky130_fd_sc_hd__and2b_1
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07529_ _09716_/A _07529_/B vssd1 vssd1 vccd1 vccd1 _07577_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_64_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07474__B1 _09568_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11270__A1 _11164_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10540_ _11384_/A _10540_/B vssd1 vssd1 vccd1 vccd1 _10542_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__09215__A1 _12838_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10471_ _10471_/A _10471_/B _10471_/C vssd1 vssd1 vccd1 vccd1 _10472_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_121_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11022__A1 _12307_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09215__B2 _12840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12210_ _12210_/A _12210_/B vssd1 vssd1 vccd1 vccd1 _12212_/B sky130_fd_sc_hd__xnor2_1
X_13190_ hold275/A _13189_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13190_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_121_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07777__B2 _07885_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07777__A1 _08723_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11573__A2 _12150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12141_ _12142_/A _12142_/B vssd1 vssd1 vccd1 vccd1 _12217_/A sky130_fd_sc_hd__nor2_1
X_12072_ _12073_/A _12073_/B vssd1 vssd1 vccd1 vccd1 _12145_/A sky130_fd_sc_hd__nor2_1
X_11023_ _11018_/Y _11019_/X _11020_/Y _11022_/X vssd1 vssd1 vccd1 vccd1 _11023_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_99_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12825__A2 _12818_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12974_ hold157/X _13016_/A2 _13016_/B1 _13290_/Q vssd1 vssd1 vccd1 vccd1 hold158/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_63_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07282__B _07282_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11925_ _12317_/A _11925_/B vssd1 vssd1 vccd1 vccd1 _11927_/B sky130_fd_sc_hd__xnor2_1
XANTENNA_clkbuf_4_0_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12628__B _12629_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11856_ _11856_/A _11856_/B vssd1 vssd1 vccd1 vccd1 _11857_/B sky130_fd_sc_hd__or2_1
XANTENNA__06626__B _07343_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09454__A1 fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11787_ _11787_/A _11787_/B vssd1 vssd1 vccd1 vccd1 _11787_/Y sky130_fd_sc_hd__nor2_1
X_10807_ _10418_/A fanout29/X fanout27/X _09745_/B vssd1 vssd1 vccd1 vccd1 _10808_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_125_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10738_ _10491_/Y _10613_/X _10614_/X vssd1 vssd1 vccd1 vccd1 _10738_/X sky130_fd_sc_hd__a21o_1
XANTENNA__10064__A2 _11171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10148__B _12316_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11013__A1 _11886_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12408_ _11876_/A _12392_/X _12395_/X _12407_/Y vssd1 vssd1 vccd1 vccd1 _12408_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__11549__C1 _11548_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10669_ _10669_/A _10669_/B _10669_/C vssd1 vssd1 vccd1 vccd1 _10681_/A sky130_fd_sc_hd__and3_1
X_13388_ instruction[14] vssd1 vssd1 vccd1 vccd1 loadstore_dest[3] sky130_fd_sc_hd__buf_12
X_12339_ _12383_/B _12337_/X _12338_/Y vssd1 vssd1 vccd1 vccd1 _12339_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_11_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10164__A _10710_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06900_ instruction[13] _06902_/B vssd1 vssd1 vccd1 vccd1 dest_idx[2] sky130_fd_sc_hd__and2_4
XANTENNA__07473__A _10710_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07880_ _07850_/X _07969_/A _07905_/B vssd1 vssd1 vccd1 vccd1 _07880_/X sky130_fd_sc_hd__o21ba_1
XANTENNA__08193__A1 fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08193__B2 _08304_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06831_ _11797_/A _06831_/B vssd1 vssd1 vccd1 vccd1 _06831_/X sky130_fd_sc_hd__or2_1
XFILLER_0_37_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06762_ _06760_/Y _06762_/B vssd1 vssd1 vccd1 vccd1 _06867_/B sky130_fd_sc_hd__nand2b_2
X_09550_ _09716_/A _09550_/B vssd1 vssd1 vccd1 vccd1 _09552_/B sky130_fd_sc_hd__xor2_1
X_08501_ _08501_/A _08501_/B vssd1 vssd1 vccd1 vccd1 _08521_/A sky130_fd_sc_hd__xnor2_1
X_09481_ _09481_/A _09481_/B vssd1 vssd1 vccd1 vccd1 _09484_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__10827__A1 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10827__B2 _10948_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06693_ _11540_/A _06693_/B vssd1 vssd1 vccd1 vccd1 _06693_/X sky130_fd_sc_hd__or2_1
XANTENNA__07153__C1 _06838_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08496__A2 _09238_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08432_ _08673_/A _08432_/B vssd1 vssd1 vccd1 vccd1 _08469_/B sky130_fd_sc_hd__or2_1
XFILLER_0_77_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08363_ _08416_/A vssd1 vssd1 vccd1 vccd1 _08363_/Y sky130_fd_sc_hd__inv_2
XANTENNA_fanout143_A _12802_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07314_ _10574_/A _12808_/A _12810_/A _10575_/A vssd1 vssd1 vccd1 vccd1 _07315_/B
+ sky130_fd_sc_hd__o22a_1
X_08294_ _08340_/B _08340_/A vssd1 vssd1 vccd1 vccd1 _08295_/C sky130_fd_sc_hd__and2b_1
XFILLER_0_6_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07245_ _10165_/A _07245_/B vssd1 vssd1 vccd1 vccd1 _07249_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_46_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09748__A2 _11847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07176_ _10448_/A _07176_/B vssd1 vssd1 vccd1 vccd1 _07603_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13088__C fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07367__B fanout9/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout300 _13242_/A vssd1 vssd1 vccd1 vccd1 _13109_/A sky130_fd_sc_hd__buf_4
X_09817_ _06811_/X _09816_/X _12388_/S vssd1 vssd1 vccd1 vccd1 _09817_/X sky130_fd_sc_hd__mux2_1
XANTENNA__07383__A _10422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09748_ _10948_/B2 _11847_/A _11766_/A fanout74/X vssd1 vssd1 vccd1 vccd1 _09749_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12268__B1 _12138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07931__A1 _08730_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07931__B2 _08038_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12807__A2 _13087_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout56_A _10941_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11710_ _11623_/A _11621_/B _11638_/A vssd1 vssd1 vccd1 vccd1 _11710_/Y sky130_fd_sc_hd__o21bai_1
X_09679_ _12244_/S _09672_/X _09677_/Y _09678_/X _09172_/B vssd1 vssd1 vccd1 vccd1
+ _09699_/C sky130_fd_sc_hd__o221a_1
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12690_ _12695_/B _12690_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[12] sky130_fd_sc_hd__and2_4
XFILLER_0_127_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11641_ _10113_/A _10883_/A _10901_/Y _12254_/A1 _11640_/X vssd1 vssd1 vccd1 vccd1
+ _11641_/X sky130_fd_sc_hd__o221a_1
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09436__A1 _12844_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07447__B1 _09768_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09436__B2 _12846_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11572_ _12317_/A _11572_/B vssd1 vssd1 vccd1 vccd1 _11575_/A sky130_fd_sc_hd__xnor2_1
X_13311_ _13311_/CLK _13311_/D vssd1 vssd1 vccd1 vccd1 hold169/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_119_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10523_ _09835_/B _10646_/B hold288/A vssd1 vssd1 vccd1 vccd1 _10523_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_25_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12464__A _12639_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13242_ _13242_/A hold300/X hold173/X vssd1 vssd1 vccd1 vccd1 _13381_/D sky130_fd_sc_hd__and3_1
X_10454_ _10454_/A _10454_/B _10454_/C vssd1 vssd1 vccd1 vccd1 _10455_/C sky130_fd_sc_hd__or3_1
X_13173_ _13245_/A hold278/X vssd1 vssd1 vccd1 vccd1 _13364_/D sky130_fd_sc_hd__and2_1
XFILLER_0_110_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10385_ _11118_/A _10385_/B vssd1 vssd1 vccd1 vccd1 _10385_/X sky130_fd_sc_hd__or2_1
XFILLER_0_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12124_ _12434_/B1 _12191_/B hold207/A vssd1 vssd1 vccd1 vccd1 _12124_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_32_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08389__A _09897_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12055_ _11876_/A _12031_/X _12032_/Y _12054_/X vssd1 vssd1 vccd1 vccd1 _12055_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__08175__A1 _08730_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11006_ reg1_val[13] curr_PC[13] vssd1 vssd1 vccd1 vccd1 _11007_/B sky130_fd_sc_hd__nand2_1
XANTENNA__07293__A _12138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08175__B2 _08038_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12957_ hold86/X _12958_/B hold250/X vssd1 vssd1 vccd1 vccd1 _13233_/B sky130_fd_sc_hd__a21boi_1
XFILLER_0_99_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12888_ hold282/A hold23/X vssd1 vssd1 vccd1 vccd1 _13154_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_114_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07686__B1 _07955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11482__A1 _11751_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11482__B2 _11558_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11908_ _11908_/A _11908_/B vssd1 vssd1 vccd1 vccd1 _11912_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_68_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11839_ _11839_/A _11839_/B vssd1 vssd1 vccd1 vccd1 _11840_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_128_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09948__A _09949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10037__A2 _10664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_36 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_718 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07030_ reg1_val[22] _07030_/B vssd1 vssd1 vccd1 vccd1 _07037_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_70_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_423 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08981_ _09445_/A _08685_/A _08677_/X _08984_/A vssd1 vssd1 vccd1 vccd1 _08982_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_11_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07932_ _08731_/A _07932_/B vssd1 vssd1 vccd1 vccd1 _07938_/A sky130_fd_sc_hd__xnor2_4
X_07863_ _08741_/B2 _08744_/A2 _08564_/B _08732_/A1 vssd1 vssd1 vccd1 vccd1 _07864_/B
+ sky130_fd_sc_hd__o22a_1
X_06814_ _10109_/A _06813_/Y _06765_/Y vssd1 vssd1 vccd1 vccd1 _06814_/Y sky130_fd_sc_hd__o21ai_1
X_09602_ _09603_/A _09603_/B vssd1 vssd1 vccd1 vccd1 _09602_/X sky130_fd_sc_hd__and2b_1
XANTENNA__11170__B1 fanout48/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09533_ _12423_/A _09497_/Y _09532_/Y _09152_/B vssd1 vssd1 vccd1 vccd1 _09533_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_64_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07794_ _07794_/A _07794_/B vssd1 vssd1 vccd1 vccd1 _07808_/B sky130_fd_sc_hd__nand2_1
X_06745_ _06805_/A _06702_/A _12673_/B _06744_/X vssd1 vssd1 vccd1 vccd1 _07095_/A
+ sky130_fd_sc_hd__a31o_4
XFILLER_0_64_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06676_ _11959_/A _11880_/A _06676_/C _11797_/A vssd1 vssd1 vccd1 vccd1 _06874_/B
+ sky130_fd_sc_hd__or4_1
X_09464_ _09465_/A _09465_/B vssd1 vssd1 vccd1 vccd1 _09466_/A sky130_fd_sc_hd__and2_1
XFILLER_0_109_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08415_ _08444_/A _08415_/B vssd1 vssd1 vccd1 vccd1 _08456_/A sky130_fd_sc_hd__xnor2_1
X_09395_ _07099_/A _07099_/B _11146_/A vssd1 vssd1 vccd1 vccd1 _09397_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_19_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08346_ _08346_/A _08346_/B vssd1 vssd1 vccd1 vccd1 _08379_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_117_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12422__B1 _12423_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08641__A2 _09238_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08277_ _08745_/A _08277_/B vssd1 vssd1 vccd1 vccd1 _08332_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07228_ _08584_/A _07228_/B vssd1 vssd1 vccd1 vccd1 _07230_/B sky130_fd_sc_hd__xnor2_1
X_07159_ reg1_val[5] _07159_/B vssd1 vssd1 vccd1 vccd1 _09898_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_30_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09593__A _09593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10170_ _10169_/A _10169_/B _10169_/C vssd1 vssd1 vccd1 vccd1 _10172_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_100_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout130 _07218_/X vssd1 vssd1 vccd1 vccd1 _10167_/A1 sky130_fd_sc_hd__buf_8
Xfanout163 _08979_/X vssd1 vssd1 vccd1 vccd1 _11633_/B sky130_fd_sc_hd__clkbuf_4
Xfanout141 _12808_/A vssd1 vssd1 vccd1 vccd1 _07885_/B sky130_fd_sc_hd__buf_6
Xfanout174 _09236_/B2 vssd1 vssd1 vccd1 vccd1 _08673_/B sky130_fd_sc_hd__clkbuf_4
Xfanout152 _10707_/A vssd1 vssd1 vccd1 vccd1 _10448_/A sky130_fd_sc_hd__buf_6
Xfanout196 _07220_/B vssd1 vssd1 vccd1 vccd1 _07074_/B sky130_fd_sc_hd__buf_4
Xfanout185 _07006_/Y vssd1 vssd1 vccd1 vccd1 _08671_/B2 sky130_fd_sc_hd__buf_8
XANTENNA__11161__B1 _12316_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07380__A2 _10570_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12811_ hold55/X _12856_/B _12810_/Y _13128_/A vssd1 vssd1 vccd1 vccd1 hold56/A sky130_fd_sc_hd__o211a_1
XFILLER_0_97_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08656__B _08656_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12742_ _12742_/A _12746_/D vssd1 vssd1 vccd1 vccd1 loadstore_address[23] sky130_fd_sc_hd__xnor2_4
XFILLER_0_96_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09409__A1 _09251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12673_ reg1_val[10] _12673_/B vssd1 vssd1 vccd1 vccd1 _12683_/A sky130_fd_sc_hd__nand2_1
X_11624_ _11624_/A _11624_/B _11624_/C vssd1 vssd1 vccd1 vccd1 _11624_/X sky130_fd_sc_hd__or3_1
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08672__A _08681_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08093__B1 _08564_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11555_ _12261_/A _11555_/B vssd1 vssd1 vccd1 vccd1 _11557_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__10707__A _10707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10506_ _06816_/X _10505_/X _12388_/S vssd1 vssd1 vccd1 vccd1 _10507_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_40_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11486_ _11486_/A _11486_/B vssd1 vssd1 vccd1 vccd1 _11488_/B sky130_fd_sc_hd__xor2_1
X_13225_ _13225_/A _13225_/B vssd1 vssd1 vccd1 vccd1 _13225_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__12177__C1 _11624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10437_ _12076_/A _10437_/B vssd1 vssd1 vccd1 vccd1 _10439_/B sky130_fd_sc_hd__xnor2_1
X_13156_ hold282/A _13155_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13156_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_103_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10368_ _10368_/A _10496_/A _10617_/A _10741_/A vssd1 vssd1 vccd1 vccd1 _10368_/X
+ sky130_fd_sc_hd__or4_2
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13087_ hold70/X _13236_/B _07504_/Y _13087_/B2 _13086_/Y vssd1 vssd1 vccd1 vccd1
+ hold71/A sky130_fd_sc_hd__o221a_1
X_12107_ _12106_/A _12106_/B _12106_/Y _09163_/X vssd1 vssd1 vccd1 vccd1 _12107_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10299_ _10413_/C _10413_/D vssd1 vssd1 vccd1 vccd1 _10302_/A sky130_fd_sc_hd__xnor2_1
X_12038_ reg1_val[24] curr_PC[24] vssd1 vssd1 vccd1 vccd1 _12038_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__11152__B1 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10161__B _10589_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07659__B1 _11751_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08320__B2 _07955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08320__A1 _07752_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08200_ _08200_/A _08200_/B vssd1 vssd1 vccd1 vccd1 _08214_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__12816__B _12818_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09180_ _11233_/S _09181_/B vssd1 vssd1 vccd1 vccd1 _09182_/B sky130_fd_sc_hd__nor2_1
XANTENNA__08582__A _08681_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08131_ _08129_/Y _08140_/B _08126_/Y vssd1 vssd1 vccd1 vccd1 _08135_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_71_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08062_ _10537_/A1 _08721_/B1 _08739_/A1 _08432_/B vssd1 vssd1 vccd1 vccd1 _08063_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_70_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07013_ _11172_/A _07013_/B vssd1 vssd1 vccd1 vccd1 _12139_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_12_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12832__A _12832_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout106_A _11987_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_776 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08964_ _08965_/A _08965_/B vssd1 vssd1 vccd1 vccd1 _08964_/X sky130_fd_sc_hd__and2_1
XANTENNA__13132__B2 _12790_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07915_ _07915_/A _07915_/B vssd1 vssd1 vccd1 vccd1 _07916_/C sky130_fd_sc_hd__xor2_1
XFILLER_0_75_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08895_ _08895_/A _08895_/B vssd1 vssd1 vccd1 vccd1 _08898_/C sky130_fd_sc_hd__xor2_1
XFILLER_0_75_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07846_ _07846_/A _07846_/B vssd1 vssd1 vccd1 vccd1 _07847_/B sky130_fd_sc_hd__xor2_1
XANTENNA__07898__B1 _11564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07777_ _08723_/B1 _09609_/B _09396_/B _07885_/B vssd1 vssd1 vccd1 vccd1 _07778_/B
+ sky130_fd_sc_hd__o22a_1
X_06728_ _07074_/A reg1_val[12] vssd1 vssd1 vccd1 vccd1 _06728_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__11446__A1 _07130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09516_ _09514_/Y _09516_/B vssd1 vssd1 vccd1 vccd1 _09517_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_79_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09447_ _10706_/B2 fanout48/X _10930_/B _10445_/A vssd1 vssd1 vccd1 vccd1 _09448_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07114__A2 _12802_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11997__A2 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06659_ _06657_/Y _06703_/B1 _06771_/A reg2_val[22] vssd1 vssd1 vccd1 vccd1 _07191_/A
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_38_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09378_ _09294_/A _09294_/B _09295_/Y vssd1 vssd1 vccd1 vccd1 _09481_/A sky130_fd_sc_hd__o21ai_4
XFILLER_0_47_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08329_ _08329_/A _08329_/B vssd1 vssd1 vccd1 vccd1 _08331_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_19_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11340_ _11341_/B _11536_/C hold292/A vssd1 vssd1 vccd1 vccd1 _11340_/X sky130_fd_sc_hd__a21o_1
XANTENNA__06724__B _11020_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10421__A2 _07087_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13010_ hold218/A _13016_/A2 _13016_/B1 hold207/X vssd1 vssd1 vccd1 vccd1 hold208/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__06673__A_N _07135_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11271_ _11271_/A fanout8/X vssd1 vssd1 vccd1 vccd1 _11272_/C sky130_fd_sc_hd__nor2_1
X_10222_ _10086_/A _10086_/B _10084_/Y vssd1 vssd1 vccd1 vccd1 _10224_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_100_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10153_ _11172_/A _10153_/B vssd1 vssd1 vccd1 vccd1 _10155_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__11382__B1 _12316_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11921__A2 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold8 hold8/A vssd1 vssd1 vccd1 vccd1 hold8/X sky130_fd_sc_hd__dlygate4sd3_1
X_10084_ _10085_/A _10085_/B vssd1 vssd1 vccd1 vccd1 _10084_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__08550__B2 _07955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08550__A1 _09423_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07353__A2 fanout94/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08302__B2 _08432_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08302__A1 _10537_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10986_ _10987_/A _10987_/B _10987_/C vssd1 vssd1 vccd1 vccd1 _10988_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_127_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12725_ _12725_/A _12725_/B _12725_/C _12725_/D vssd1 vssd1 vccd1 vccd1 _12728_/B
+ sky130_fd_sc_hd__or4_2
XFILLER_0_72_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12656_ _12656_/A _12656_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[6] sky130_fd_sc_hd__xor2_4
X_12587_ _12611_/A _12587_/B vssd1 vssd1 vccd1 vccd1 _12595_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__11540__B _11973_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11607_ _11420_/Y _11787_/A _11605_/Y vssd1 vssd1 vccd1 vccd1 _11607_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_25_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10437__A _12076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10948__B1 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11538_ hold263/A _11341_/B _11635_/B _09837_/A vssd1 vssd1 vccd1 vccd1 _11539_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_111_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11469_ _11469_/A _11469_/B vssd1 vssd1 vccd1 vccd1 _11478_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_0_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13208_ hold254/X _13207_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13208_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_110_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13139_ _12893_/X _13139_/B vssd1 vssd1 vccd1 vccd1 _13140_/B sky130_fd_sc_hd__nand2b_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11125__B1 _12247_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07700_ _08727_/A2 _11847_/A _11923_/A _08727_/B1 vssd1 vssd1 vccd1 vccd1 _07701_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08680_ _08680_/A _09364_/A vssd1 vssd1 vccd1 vccd1 _08985_/A sky130_fd_sc_hd__or2_2
X_07631_ _07631_/A _07631_/B vssd1 vssd1 vccd1 vccd1 _08919_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_45_74 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07562_ _07562_/A _07562_/B vssd1 vssd1 vccd1 vccd1 _07567_/A sky130_fd_sc_hd__and2_2
XFILLER_0_76_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09301_ _09302_/A _09302_/B vssd1 vssd1 vccd1 vccd1 _09301_/X sky130_fd_sc_hd__and2_1
XFILLER_0_48_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07493_ _09444_/A _12852_/A _12854_/A _09236_/B2 vssd1 vssd1 vccd1 vccd1 _07494_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_76_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09232_ _09232_/A _09232_/B vssd1 vssd1 vccd1 vccd1 _09235_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_35_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09163_ _09163_/A _09170_/A vssd1 vssd1 vccd1 vccd1 _09163_/X sky130_fd_sc_hd__or2_4
XFILLER_0_8_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout223_A _06890_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08114_ _08721_/B1 fanout87/X fanout82/X _08739_/A1 vssd1 vssd1 vccd1 vccd1 _08115_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_16_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09094_ _09092_/X _09093_/X _09330_/S vssd1 vssd1 vccd1 vccd1 _09094_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_71_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08045_ _08042_/B _08042_/C _08042_/A vssd1 vssd1 vccd1 vccd1 _08046_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_3_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10167__A1 _10167_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10167__B2 _07222_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09309__B1 _12290_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09996_ curr_PC[3] curr_PC[4] _09701_/B curr_PC[5] vssd1 vssd1 vccd1 vccd1 _09996_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__12313__C1 _06881_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08947_ _08948_/B _08948_/A vssd1 vssd1 vccd1 vccd1 _08947_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_98_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11667__B2 _07819_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11667__A1 fanout24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11906__A _12210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08878_ _08878_/A _08878_/B vssd1 vssd1 vccd1 vccd1 _08880_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__07335__A2 _10022_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07829_ _11758_/A _07829_/B vssd1 vssd1 vccd1 vccd1 _07831_/B sky130_fd_sc_hd__xnor2_1
X_10840_ _10704_/B _10717_/B _10704_/A vssd1 vssd1 vccd1 vccd1 _10850_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_94_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10771_ hold285/A _11341_/B _10893_/B _09837_/A vssd1 vssd1 vccd1 vccd1 _10771_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_67_746 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_5_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12510_ _12516_/B _12510_/B vssd1 vssd1 vccd1 vccd1 new_PC[9] sky130_fd_sc_hd__and2_4
XFILLER_0_124_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12441_ _06923_/Y _12430_/X _12440_/X _12428_/X vssd1 vssd1 vccd1 vccd1 _12441_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__11360__B _11649_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08048__B1 _11908_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08599__A1 _08646_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08599__B2 _09423_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12372_ _12372_/A _12372_/B vssd1 vssd1 vccd1 vccd1 _12373_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_34_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11323_ _11421_/B _11323_/B vssd1 vssd1 vccd1 vccd1 _11649_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11254_ _12448_/S _11357_/C vssd1 vssd1 vccd1 vccd1 _11254_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_120_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11355__B1 _11142_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10205_ _10205_/A _10205_/B vssd1 vssd1 vccd1 vccd1 _10206_/B sky130_fd_sc_hd__nor2_1
XANTENNA__08220__B1 _08564_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11185_ _11185_/A vssd1 vssd1 vccd1 vccd1 _11187_/B sky130_fd_sc_hd__inv_2
X_10136_ _10109_/Y _10110_/X _10135_/X vssd1 vssd1 vccd1 vccd1 _10136_/X sky130_fd_sc_hd__a21o_1
X_10067_ _11261_/A _10067_/B vssd1 vssd1 vccd1 vccd1 _10069_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__09720__B1 _10567_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06629__B _12673_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10945__B1_N _10448_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10969_ _10969_/A _10969_/B vssd1 vssd1 vccd1 vccd1 _10983_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_128_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12708_ reg1_val[16] _12741_/B vssd1 vssd1 vccd1 vccd1 _12709_/B sky130_fd_sc_hd__and2_1
XFILLER_0_115_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08039__B1 _07149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13032__B1 _06892_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12639_ reg1_val[3] _12639_/B vssd1 vssd1 vccd1 vccd1 _12640_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_25_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold216 hold216/A vssd1 vssd1 vccd1 vccd1 hold216/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold205 hold228/X vssd1 vssd1 vccd1 vccd1 hold205/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold227 hold227/A vssd1 vssd1 vccd1 vccd1 hold227/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold249 hold249/A vssd1 vssd1 vccd1 vccd1 hold249/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold238 hold238/A vssd1 vssd1 vccd1 vccd1 hold238/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07014__A1 _12076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11897__B2 _12254_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09850_ curr_PC[4] _09997_/C vssd1 vssd1 vccd1 vccd1 _09850_/Y sky130_fd_sc_hd__nand2_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06773__B1 _12429_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06993_ _07374_/A _06993_/B vssd1 vssd1 vccd1 vccd1 _07057_/A sky130_fd_sc_hd__and2_1
X_09781_ _09782_/A _09782_/B vssd1 vssd1 vccd1 vccd1 _09912_/A sky130_fd_sc_hd__nand2_1
X_08801_ _08801_/A _08801_/B vssd1 vssd1 vccd1 vccd1 _08805_/A sky130_fd_sc_hd__xor2_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08732_ _08732_/A1 _08732_/A2 _08656_/B _10927_/A1 vssd1 vssd1 vccd1 vccd1 _08733_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08663_ _08730_/A1 _07752_/B _08436_/B _07821_/A vssd1 vssd1 vccd1 vccd1 _08664_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout173_A _09236_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08100__A _08728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08594_ _08594_/A _08594_/B vssd1 vssd1 vccd1 vccd1 _08611_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__10872__A2 _10871_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07614_ _07624_/B _07993_/A _07624_/A vssd1 vssd1 vccd1 vccd1 _07627_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_119_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07545_ _07545_/A _07545_/B vssd1 vssd1 vccd1 vccd1 _07555_/A sky130_fd_sc_hd__xnor2_2
X_07476_ _07477_/A _07477_/B vssd1 vssd1 vccd1 vccd1 _07478_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_76_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11821__A1 _11142_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11461__A _12073_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09215_ _12838_/A _10589_/A _08507_/B _12840_/A vssd1 vssd1 vccd1 vccd1 _09216_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_91_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09146_ _10385_/B _09145_/X _11231_/S vssd1 vssd1 vccd1 vccd1 _09146_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09866__A _11172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09077_ _09077_/A _09077_/B _12392_/A _12426_/C vssd1 vssd1 vccd1 vccd1 _10658_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_71_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08028_ _08028_/A _08028_/B vssd1 vssd1 vccd1 vccd1 _08078_/A sky130_fd_sc_hd__xnor2_1
X_09979_ hold187/A _10120_/C _10391_/A2 vssd1 vssd1 vccd1 vccd1 _09980_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__06764__B1 _06763_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10540__A _11384_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12990_ hold205/X _13004_/A2 _13006_/B1 hold183/X vssd1 vssd1 vccd1 vccd1 hold206/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_98_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11941_ _11943_/A _11943_/B _11943_/C vssd1 vssd1 vccd1 vccd1 _11942_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_98_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11872_ _11874_/A _11872_/B _11872_/C vssd1 vssd1 vccd1 vccd1 _11872_/X sky130_fd_sc_hd__and3_1
XFILLER_0_67_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10823_ _10823_/A vssd1 vssd1 vccd1 vccd1 _10825_/A sky130_fd_sc_hd__inv_2
XFILLER_0_109_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11812__A1 _12307_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10754_ reg1_val[11] curr_PC[11] vssd1 vssd1 vccd1 vccd1 _10754_/X sky130_fd_sc_hd__or2_1
XFILLER_0_82_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10685_ _12076_/A _10685_/B vssd1 vssd1 vccd1 vccd1 _10689_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__11025__C1 _11023_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12424_ _12422_/X _12423_/Y _08980_/B vssd1 vssd1 vccd1 vccd1 _12424_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__09233__A2 _12830_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12355_ hold169/A _12355_/B vssd1 vssd1 vccd1 vccd1 _12399_/B sky130_fd_sc_hd__or2_1
XANTENNA__07244__B2 _09567_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07244__A1 _12838_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11576__B1 _12067_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07296__A _10165_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11306_ _11306_/A _11306_/B vssd1 vssd1 vccd1 vccd1 _11308_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12286_ _12170_/B _12286_/B vssd1 vssd1 vccd1 vccd1 _12287_/B sky130_fd_sc_hd__nand2b_2
X_11237_ hold183/A _11346_/B vssd1 vssd1 vccd1 vccd1 _11237_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__07547__A2 fanout16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08744__A1 fanout99/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08744__B2 _12818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11168_ _11168_/A _11168_/B vssd1 vssd1 vccd1 vccd1 _11169_/B sky130_fd_sc_hd__nor2_1
X_10119_ _10116_/X _10118_/X _10119_/S vssd1 vssd1 vccd1 vccd1 _10119_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_93_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11099_ _10857_/Y _10988_/A _10988_/B vssd1 vssd1 vccd1 vccd1 _11319_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_26_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12056__A1 _11707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07330_ _12842_/A _09568_/B _12840_/A _09567_/B vssd1 vssd1 vccd1 vccd1 _07331_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_46_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09000_ _09000_/A _09000_/B vssd1 vssd1 vccd1 vccd1 _10503_/C sky130_fd_sc_hd__or2_1
X_07261_ _12076_/A _07263_/B _10928_/A vssd1 vssd1 vccd1 vccd1 _07262_/B sky130_fd_sc_hd__a21boi_1
XFILLER_0_115_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12359__A2 _09354_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07192_ _07187_/B _10024_/A vssd1 vssd1 vccd1 vccd1 _07192_/Y sky130_fd_sc_hd__nand2b_2
XFILLER_0_26_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12824__B _12830_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07235__B2 _09238_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07235__A1 _12842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10909__A3 _10871_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06734__A_N _06963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10790__A1 _10571_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10790__B2 _10570_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12840__A _12840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09902_ _10448_/A _09902_/B vssd1 vssd1 vccd1 vccd1 _09910_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_1_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09833_ hold187/A _10391_/A2 _10120_/C _11968_/B1 vssd1 vssd1 vccd1 vccd1 _09833_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07934__A _08733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout290_A _06799_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06976_ reg1_val[13] _06994_/D _07200_/A vssd1 vssd1 vccd1 vccd1 _06982_/B sky130_fd_sc_hd__o21a_1
X_09764_ _09764_/A _09764_/B vssd1 vssd1 vccd1 vccd1 _09765_/B sky130_fd_sc_hd__xor2_2
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09695_ _06789_/Y _12403_/A1 _12402_/A0 _09686_/B _09694_/X vssd1 vssd1 vccd1 vccd1
+ _09695_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_96_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08715_ _08382_/Y _08715_/B vssd1 vssd1 vccd1 vccd1 _09026_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__09160__A1 _11624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08646_ _08671_/B2 _08661_/A2 _08673_/B _08646_/B2 vssd1 vssd1 vccd1 vccd1 _08647_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_68_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08577_ _08577_/A _08577_/B vssd1 vssd1 vccd1 vccd1 _08584_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_76_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07528_ _09768_/A1 fanout23/X _11171_/A _12808_/A vssd1 vssd1 vccd1 vccd1 _07529_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_64_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07474__A1 _12844_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07474__B2 _12846_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07459_ _07459_/A _07459_/B vssd1 vssd1 vccd1 vccd1 _07560_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__08671__B1 _08436_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11270__A2 _07076_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10470_ _10471_/A _10471_/B _10471_/C vssd1 vssd1 vccd1 vccd1 _10603_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_17_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09129_ _09125_/X _09128_/X _09669_/S vssd1 vssd1 vccd1 vccd1 _09129_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09215__A2 _10589_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06732__B _06799_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07777__A2 _09609_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12140_ _07012_/X _12412_/A _12139_/Y _12076_/A vssd1 vssd1 vccd1 vccd1 _12142_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12071_ _12317_/A _12071_/B vssd1 vssd1 vccd1 vccd1 _12073_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_4_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11022_ _12307_/B1 _11021_/X _06725_/B vssd1 vssd1 vccd1 vccd1 _11022_/X sky130_fd_sc_hd__a21o_1
XANTENNA__11366__A _12317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12973_ _13009_/A hold186/X vssd1 vssd1 vccd1 vccd1 _13289_/D sky130_fd_sc_hd__and2_1
XANTENNA__06752__A3 _12669_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09151__A1 _12429_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10297__B1 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11924_ _12150_/A fanout15/X fanout36/X _12213_/A vssd1 vssd1 vccd1 vccd1 _11925_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_86_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08675__A _08728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06907__B _06921_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10049__B1 _10930_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11855_ _11856_/A _11856_/B vssd1 vssd1 vccd1 vccd1 _11943_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_28_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09454__A2 _10574_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11786_ _11605_/Y _11787_/B _11784_/Y vssd1 vssd1 vccd1 vccd1 _12099_/A sky130_fd_sc_hd__o21ai_1
X_10806_ _11180_/A _10806_/B vssd1 vssd1 vccd1 vccd1 _10810_/A sky130_fd_sc_hd__xnor2_1
X_10737_ _10737_/A _10737_/B vssd1 vssd1 vccd1 vccd1 _11102_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_27_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12407_ _12397_/Y _12398_/X _12406_/X vssd1 vssd1 vccd1 vccd1 _12407_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_113_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10668_ _10959_/A _10668_/B vssd1 vssd1 vccd1 vccd1 _10669_/C sky130_fd_sc_hd__or2_1
XANTENNA__12644__B _12644_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13387_ instruction[13] vssd1 vssd1 vccd1 vccd1 loadstore_dest[2] sky130_fd_sc_hd__buf_12
X_10599_ _10441_/A _10441_/B _10429_/X vssd1 vssd1 vccd1 vccd1 _10601_/A sky130_fd_sc_hd__a21o_1
XANTENNA__10445__A _10445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06976__B1 _07200_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12338_ _12383_/B _12337_/X _11707_/A vssd1 vssd1 vccd1 vccd1 _12338_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_23_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12269_ _12210_/A _12317_/A _07263_/B _12412_/A _12268_/X vssd1 vssd1 vccd1 vccd1
+ _12321_/B sky130_fd_sc_hd__a41o_1
XANTENNA__09914__B1 _07036_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08193__A2 _07821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06830_ reg1_val[20] _07223_/A vssd1 vssd1 vccd1 vccd1 _06831_/B sky130_fd_sc_hd__nand2_1
X_06761_ reg1_val[7] _07080_/A vssd1 vssd1 vccd1 vccd1 _06762_/B sky130_fd_sc_hd__nand2_1
X_06692_ _11540_/A _06693_/B vssd1 vssd1 vccd1 vccd1 _06866_/B sky130_fd_sc_hd__nor2_1
X_08500_ _08501_/A _08501_/B vssd1 vssd1 vccd1 vccd1 _08500_/X sky130_fd_sc_hd__or2_1
X_09480_ _09480_/A _09480_/B vssd1 vssd1 vccd1 vccd1 _09481_/B sky130_fd_sc_hd__xor2_4
XANTENNA__10827__A2 _09568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08431_ _08740_/A _08431_/B vssd1 vssd1 vccd1 vccd1 _08469_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08362_ _09445_/A _08362_/B vssd1 vssd1 vccd1 vccd1 _08416_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_85_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07313_ _07522_/A _07313_/B vssd1 vssd1 vccd1 vccd1 _07317_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_46_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08293_ _08293_/A _08293_/B vssd1 vssd1 vccd1 vccd1 _08340_/B sky130_fd_sc_hd__xnor2_1
X_07244_ _12838_/A _09568_/B _12836_/A _09567_/B vssd1 vssd1 vccd1 vccd1 _07245_/B
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_73_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout136_A _12814_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07929__A _11908_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07175_ _11294_/A _10706_/B2 _08732_/A1 _10445_/A vssd1 vssd1 vccd1 vccd1 _07176_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_42_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10763__A1 _12244_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout301 _13242_/A vssd1 vssd1 vccd1 vccd1 _13245_/A sky130_fd_sc_hd__buf_4
XANTENNA__09905__B1 _11923_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11712__B1 _09156_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09816_ _06789_/Y _09684_/B _09684_/C _06791_/B vssd1 vssd1 vccd1 vccd1 _09816_/X
+ sky130_fd_sc_hd__o31a_1
X_06959_ _11231_/S _10248_/S _09666_/S _09351_/B vssd1 vssd1 vccd1 vccd1 _06964_/A
+ sky130_fd_sc_hd__or4_4
X_09747_ _09746_/B _09746_/C _09746_/A vssd1 vssd1 vccd1 vccd1 _09751_/B sky130_fd_sc_hd__a21o_1
XANTENNA__12268__A1 fanout16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07931__A2 _11847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10279__B1 _10570_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09678_ _09673_/X _09675_/X _09676_/Y _11886_/A vssd1 vssd1 vccd1 vccd1 _09678_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08629_ _08637_/B _08637_/A vssd1 vssd1 vccd1 vccd1 _08629_/X sky130_fd_sc_hd__and2b_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11640_ _07210_/A _11343_/B _11639_/X _06683_/B vssd1 vssd1 vccd1 vccd1 _11640_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_83_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09436__A2 _10167_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12440__A1 _09169_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07447__A1 fanout30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07447__B2 _07688_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11571_ _11847_/A fanout15/X fanout36/X _11923_/A vssd1 vssd1 vccd1 vccd1 _11572_/B
+ sky130_fd_sc_hd__o22a_1
X_13310_ _13314_/CLK _13310_/D vssd1 vssd1 vccd1 vccd1 hold195/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10522_ hold273/A hold294/A _10522_/C vssd1 vssd1 vccd1 vccd1 _10646_/B sky130_fd_sc_hd__or3_2
XFILLER_0_91_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13241_ hold172/X hold63/X hold166/X vssd1 vssd1 vccd1 vccd1 hold173/A sky130_fd_sc_hd__a21o_1
X_10453_ _10454_/A _10454_/B _10454_/C vssd1 vssd1 vccd1 vccd1 _10455_/B sky130_fd_sc_hd__o21ai_1
X_13172_ hold277/X _06890_/Y _13171_/X _13246_/B2 vssd1 vssd1 vccd1 vccd1 hold278/A
+ sky130_fd_sc_hd__a22o_1
X_10384_ _10384_/A _10384_/B vssd1 vssd1 vccd1 vccd1 _10384_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_60_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12123_ hold218/A _12123_/B vssd1 vssd1 vccd1 vccd1 _12191_/B sky130_fd_sc_hd__or2_1
X_12054_ _09172_/B _12042_/X _12053_/Y _12036_/X vssd1 vssd1 vccd1 vccd1 _12054_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__08175__A2 _10927_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11005_ reg1_val[13] curr_PC[13] vssd1 vssd1 vccd1 vccd1 _11007_/A sky130_fd_sc_hd__or2_1
XANTENNA__12259__A1 _11673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12956_ _12860_/B _13229_/B _12860_/A vssd1 vssd1 vccd1 vccd1 _12958_/B sky130_fd_sc_hd__o21ba_1
XFILLER_0_87_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12639__B _12639_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12887_ hold23/X hold282/A vssd1 vssd1 vccd1 vccd1 _12887_/X sky130_fd_sc_hd__and2b_1
XANTENNA__07686__A1 _09613_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07686__B2 _09614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11482__A2 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11907_ _11908_/A _11908_/B vssd1 vssd1 vccd1 vccd1 _11992_/A sky130_fd_sc_hd__and2b_1
XTAP_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10690__B1 _10574_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11838_ _11839_/A _11839_/B vssd1 vssd1 vccd1 vccd1 _11915_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09948__B _09949_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11769_ _11767_/X _11769_/B vssd1 vssd1 vccd1 vccd1 _11770_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_126_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08980_ _12423_/A _08980_/B vssd1 vssd1 vccd1 vccd1 _08980_/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07931_ _08730_/A1 _11847_/A _11766_/A _08038_/A vssd1 vssd1 vccd1 vccd1 _07932_/B
+ sky130_fd_sc_hd__o22a_2
XANTENNA__09363__A1 _09442_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07862_ _07862_/A _07862_/B vssd1 vssd1 vccd1 vccd1 _07912_/A sky130_fd_sc_hd__xor2_1
X_06813_ _09964_/A _06812_/X _06774_/X vssd1 vssd1 vccd1 vccd1 _06813_/Y sky130_fd_sc_hd__a21oi_1
X_09601_ _12264_/B _09601_/B vssd1 vssd1 vccd1 vccd1 _09603_/B sky130_fd_sc_hd__xnor2_2
X_09532_ _12423_/A _09532_/B vssd1 vssd1 vccd1 vccd1 _09532_/Y sky130_fd_sc_hd__nor2_1
X_07793_ _07881_/A _07881_/B _07789_/X vssd1 vssd1 vccd1 vccd1 _07810_/A sky130_fd_sc_hd__o21ai_2
X_06744_ reg2_val[9] _06799_/B vssd1 vssd1 vccd1 vccd1 _06744_/X sky130_fd_sc_hd__and2_1
X_06675_ _11811_/S _06675_/B vssd1 vssd1 vccd1 vccd1 _11797_/A sky130_fd_sc_hd__nor2_2
X_09463_ _09463_/A _09463_/B vssd1 vssd1 vccd1 vccd1 _09465_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_66_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09394_ _09203_/A _09203_/B _09200_/A vssd1 vssd1 vccd1 vccd1 _09413_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_59_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08414_ _08414_/A _08414_/B vssd1 vssd1 vccd1 vccd1 _08415_/B sky130_fd_sc_hd__or2_1
X_08345_ _08345_/A _08345_/B vssd1 vssd1 vccd1 vccd1 _08346_/B sky130_fd_sc_hd__or2_1
XFILLER_0_19_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08276_ _08723_/B1 _08744_/A2 _08564_/B _07885_/B vssd1 vssd1 vccd1 vccd1 _08277_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_6_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07227_ _10167_/A1 _12834_/A _10022_/B1 _12836_/A vssd1 vssd1 vccd1 vccd1 _07228_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_14_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07158_ reg1_val[5] _07159_/B vssd1 vssd1 vccd1 vccd1 _09897_/A sky130_fd_sc_hd__xor2_4
XANTENNA__09874__A _11470_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09085__S _09108_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07089_ _07089_/A _07089_/B vssd1 vssd1 vccd1 vccd1 _07089_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_0_2_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout131 _09567_/B vssd1 vssd1 vccd1 vccd1 _08741_/A2 sky130_fd_sc_hd__buf_8
Xfanout120 _12828_/A vssd1 vssd1 vccd1 vccd1 _11367_/A sky130_fd_sc_hd__buf_6
Xfanout164 _10391_/A2 vssd1 vssd1 vccd1 vccd1 _12434_/B1 sky130_fd_sc_hd__buf_4
Xfanout142 _10148_/A vssd1 vssd1 vccd1 vccd1 _12808_/A sky130_fd_sc_hd__buf_8
Xfanout153 _08722_/A vssd1 vssd1 vccd1 vccd1 _10707_/A sky130_fd_sc_hd__buf_8
Xfanout197 _12791_/Y vssd1 vssd1 vccd1 vccd1 _13087_/B2 sky130_fd_sc_hd__buf_4
Xfanout186 _08740_/A vssd1 vssd1 vccd1 vccd1 _10710_/A sky130_fd_sc_hd__buf_12
Xfanout175 _07139_/Y vssd1 vssd1 vccd1 vccd1 _09236_/B2 sky130_fd_sc_hd__buf_4
XANTENNA__11161__A1 _09609_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11161__B2 _09396_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12810_ _12810_/A _12856_/B vssd1 vssd1 vccd1 vccd1 _12810_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_97_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12741_ reg1_val[23] _12741_/B vssd1 vssd1 vccd1 vccd1 _12746_/D sky130_fd_sc_hd__xnor2_4
XFILLER_0_84_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12672_ reg1_val[10] _12673_/B vssd1 vssd1 vccd1 vccd1 _12674_/A sky130_fd_sc_hd__or2_1
X_11623_ _11623_/A _11623_/B _11623_/C vssd1 vssd1 vccd1 vccd1 _11624_/C sky130_fd_sc_hd__and3_1
XANTENNA__09409__A2 _12264_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08093__A1 _08436_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11554_ _11766_/A fanout9/X fanout4/X _11751_/A vssd1 vssd1 vccd1 vccd1 _11555_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08093__B2 fanout99/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10505_ _06754_/Y _10376_/X _06756_/B vssd1 vssd1 vccd1 vccd1 _10505_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_80_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11485_ _12210_/A _11485_/B vssd1 vssd1 vccd1 vccd1 _11486_/B sky130_fd_sc_hd__xnor2_1
X_13224_ _12861_/X _13224_/B vssd1 vssd1 vccd1 vccd1 _13225_/B sky130_fd_sc_hd__nand2b_1
X_10436_ _11065_/A fanout30/X _07688_/B _11146_/A vssd1 vssd1 vccd1 vccd1 _10437_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11924__B1 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13155_ _13155_/A _13155_/B vssd1 vssd1 vccd1 vccd1 _13155_/Y sky130_fd_sc_hd__xnor2_1
X_10367_ _10100_/A _10366_/Y _10365_/Y vssd1 vssd1 vccd1 vccd1 _10864_/A sky130_fd_sc_hd__a21oi_2
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13086_ _06566_/Y _06572_/A rst vssd1 vssd1 vccd1 vccd1 _13086_/Y sky130_fd_sc_hd__a21oi_1
X_12106_ _12106_/A _12106_/B vssd1 vssd1 vccd1 vccd1 _12106_/Y sky130_fd_sc_hd__nor2_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10298_ _11163_/A _10298_/B vssd1 vssd1 vccd1 vccd1 _10413_/D sky130_fd_sc_hd__xnor2_1
X_12037_ _11964_/A _11964_/B _11962_/B vssd1 vssd1 vccd1 vccd1 _12041_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_18_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11152__B2 _11558_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11152__A1 _11472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07108__B1 _07688_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12939_ _12877_/X _12939_/B vssd1 vssd1 vccd1 vccd1 _13184_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_88_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07659__A1 _09567_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07659__B2 _09568_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08320__A2 fanout87/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08130_ _08130_/A _08130_/B vssd1 vssd1 vccd1 vccd1 _08140_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_28_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08061_ _08067_/A _08067_/B vssd1 vssd1 vccd1 vccd1 _08061_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_114_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07012_ _12076_/A _11172_/A _07013_/B vssd1 vssd1 vccd1 vccd1 _07012_/X sky130_fd_sc_hd__and3b_1
XFILLER_0_3_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06830__B _07223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08963_ _08965_/A _08965_/B vssd1 vssd1 vccd1 vccd1 _08963_/X sky130_fd_sc_hd__or2_1
XANTENNA__13132__A2 _12789_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07914_ _07913_/A _07913_/B _07913_/C vssd1 vssd1 vccd1 vccd1 _07916_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_75_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08894_ _08895_/B _08895_/A vssd1 vssd1 vccd1 vccd1 _08901_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_79_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07845_ _07846_/A _07846_/B vssd1 vssd1 vccd1 vccd1 _07845_/Y sky130_fd_sc_hd__nand2_1
X_07776_ _07776_/A _07776_/B vssd1 vssd1 vccd1 vccd1 _07811_/A sky130_fd_sc_hd__xor2_1
XANTENNA__11446__A2 _11343_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09515_ reg1_val[2] curr_PC[2] vssd1 vssd1 vccd1 vccd1 _09516_/B sky130_fd_sc_hd__nand2_1
X_06727_ _06805_/A _06702_/A _12692_/B _06726_/X vssd1 vssd1 vccd1 vccd1 _07074_/A
+ sky130_fd_sc_hd__a31o_4
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09446_ _09446_/A _09446_/B vssd1 vssd1 vccd1 vccd1 _09459_/A sky130_fd_sc_hd__xnor2_2
XPHY_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06658_ reg2_val[22] _06771_/A _06703_/B1 _06657_/Y vssd1 vssd1 vccd1 vccd1 _07135_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_66_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06589_ instruction[1] instruction[2] instruction[0] pred_val vssd1 vssd1 vccd1 vccd1
+ _06589_/X sky130_fd_sc_hd__or4bb_4
X_09377_ _09299_/A _09299_/B _09297_/X vssd1 vssd1 vccd1 vccd1 _09484_/A sky130_fd_sc_hd__a21oi_4
XFILLER_0_62_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10808__A _12210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08328_ _08349_/A _08349_/B _08317_/Y vssd1 vssd1 vccd1 vccd1 _08335_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_105_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08259_ _08724_/A _08259_/B vssd1 vssd1 vccd1 vccd1 _08330_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__10421__A3 _10575_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11270_ _11164_/A _07076_/B fanout6/X _11470_/A vssd1 vssd1 vccd1 vccd1 _11272_/B
+ sky130_fd_sc_hd__o31a_1
X_10221_ _10221_/A _10221_/B vssd1 vssd1 vccd1 vccd1 _10224_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__11382__A1 _11653_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11382__B2 _08752_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10152_ _11065_/A fanout23/X _11171_/A _11146_/A vssd1 vssd1 vccd1 vccd1 _10153_/B
+ sky130_fd_sc_hd__o22a_1
X_10083_ _09929_/A _09928_/B _09928_/A vssd1 vssd1 vccd1 vccd1 _10085_/B sky130_fd_sc_hd__o21ba_1
Xhold9 hold9/A vssd1 vssd1 vccd1 vccd1 hold9/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08550__A2 _09238_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08302__A2 _08671_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10985_ _10985_/A _10985_/B vssd1 vssd1 vccd1 vccd1 _10987_/C sky130_fd_sc_hd__xor2_1
X_12724_ reg1_val[20] _12741_/B vssd1 vssd1 vccd1 vccd1 _12746_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_127_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06915__B _06921_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12655_ _12655_/A _12655_/B vssd1 vssd1 vccd1 vccd1 _12656_/B sky130_fd_sc_hd__or2_2
X_12586_ reg1_val[21] curr_PC[21] _12586_/S vssd1 vssd1 vccd1 vccd1 _12587_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_38_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11606_ _11606_/A _11700_/A vssd1 vssd1 vccd1 vccd1 _11787_/A sky130_fd_sc_hd__or2_2
X_11537_ _11341_/B _11635_/B hold263/A vssd1 vssd1 vccd1 vccd1 _11539_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_53_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10948__B2 _10948_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10948__A1 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11468_ _11908_/A _11468_/B vssd1 vssd1 vccd1 vccd1 _11469_/B sky130_fd_sc_hd__xnor2_1
X_13207_ _13207_/A _13207_/B vssd1 vssd1 vccd1 vccd1 _13207_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_110_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11399_ _11288_/A _11288_/B _11296_/X vssd1 vssd1 vccd1 vccd1 _11410_/A sky130_fd_sc_hd__o21ba_1
X_10419_ _11172_/A _10419_/B _10419_/C vssd1 vssd1 vccd1 vccd1 _10424_/A sky130_fd_sc_hd__nand3_1
X_13138_ _13235_/A hold270/X vssd1 vssd1 vccd1 vccd1 _13357_/D sky130_fd_sc_hd__and2_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13069_ _07037_/B _13077_/A2 hold127/X vssd1 vssd1 vccd1 vccd1 _13337_/D sky130_fd_sc_hd__o21a_1
XANTENNA__07762__A _08722_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07630_ _07631_/A _07631_/B vssd1 vssd1 vccd1 vccd1 _07630_/X sky130_fd_sc_hd__and2b_1
XANTENNA__11284__A _12210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07561_ _07561_/A _07561_/B vssd1 vssd1 vccd1 vccd1 _07562_/B sky130_fd_sc_hd__or2_1
XFILLER_0_45_86 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09300_ _09302_/A _09302_/B vssd1 vssd1 vccd1 vccd1 _09300_/X sky130_fd_sc_hd__or2_1
XFILLER_0_48_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07492_ _09209_/B _07492_/B vssd1 vssd1 vccd1 vccd1 _07501_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_8_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09231_ _09231_/A _09231_/B vssd1 vssd1 vccd1 vccd1 _09232_/B sky130_fd_sc_hd__or2_1
XANTENNA__11223__S _12174_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09162_ _09163_/A _09170_/A vssd1 vssd1 vccd1 vccd1 _12428_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_16_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08113_ _08722_/A _08113_/B vssd1 vssd1 vccd1 vccd1 _08120_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_16_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09093_ reg1_val[6] reg1_val[25] _09108_/S vssd1 vssd1 vccd1 vccd1 _09093_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_43_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08044_ _08598_/A _08044_/B vssd1 vssd1 vccd1 vccd1 _08046_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07937__A _08598_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10363__A _10364_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10167__A2 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09995_ _09958_/X _09959_/Y _09961_/Y _11876_/A _09994_/X vssd1 vssd1 vccd1 vccd1
+ _09995_/X sky130_fd_sc_hd__a221o_1
X_08946_ _08946_/A _08946_/B vssd1 vssd1 vccd1 vccd1 _08948_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__11667__A2 _12213_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08877_ _08878_/A _08878_/B vssd1 vssd1 vccd1 vccd1 _08877_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__10875__B1 _11876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07828_ _07752_/B _07087_/A _07087_/B _08752_/B _07955_/A vssd1 vssd1 vccd1 vccd1
+ _07829_/B sky130_fd_sc_hd__o32a_1
XFILLER_0_79_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07759_ _07759_/A _07759_/B _07759_/C vssd1 vssd1 vccd1 vccd1 _07814_/A sky130_fd_sc_hd__and3_1
XANTENNA__11922__A _12261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10770_ _11452_/B1 _10893_/B hold285/A vssd1 vssd1 vccd1 vccd1 _10770_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__09493__B1 _09163_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout31_A _12412_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09429_ _09429_/A _09429_/B vssd1 vssd1 vccd1 vccd1 _09462_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_54_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10538__A _10707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12440_ _09169_/Y _12435_/Y _12439_/X vssd1 vssd1 vccd1 vccd1 _12440_/X sky130_fd_sc_hd__a21o_1
XANTENNA__06735__B _06963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08048__A1 _08752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08599__A2 _08732_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11052__B1 _10570_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12371_ _12372_/A _12371_/B vssd1 vssd1 vccd1 vccd1 _12371_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_34_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11322_ _10371_/B _10862_/A _11320_/Y _11321_/X vssd1 vssd1 vccd1 vccd1 _11323_/B
+ sky130_fd_sc_hd__a31o_4
XFILLER_0_22_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11253_ curr_PC[15] _11253_/B vssd1 vssd1 vccd1 vccd1 _11357_/C sky130_fd_sc_hd__and2_1
X_10204_ _10205_/A _10205_/B vssd1 vssd1 vccd1 vccd1 _10204_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__08220__A1 _07885_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11184_ _11182_/X _11184_/B vssd1 vssd1 vccd1 vccd1 _11185_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__08220__B2 _08721_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10135_ _09830_/A _10119_/X _10134_/X _10113_/Y vssd1 vssd1 vccd1 vccd1 _10135_/X
+ sky130_fd_sc_hd__a211o_1
X_10066_ _10418_/A _07087_/X fanout66/X _09745_/B vssd1 vssd1 vccd1 vccd1 _10067_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09720__B2 _07688_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09720__A1 fanout30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07731__B1 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10968_ _10967_/B _10967_/C _10967_/A vssd1 vssd1 vccd1 vccd1 _10969_/B sky130_fd_sc_hd__a21oi_1
X_12707_ reg1_val[16] _12741_/B vssd1 vssd1 vccd1 vccd1 _12709_/A sky130_fd_sc_hd__nor2_1
XANTENNA__10448__A _10448_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10899_ _07074_/A _12404_/A _10896_/Y _10898_/Y vssd1 vssd1 vccd1 vccd1 _10899_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__06645__B _07166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12638_ reg1_val[3] _12639_/B vssd1 vssd1 vccd1 vccd1 _12638_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_26_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09236__B1 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11043__B1 _11163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10397__A2 _09354_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12569_ _12581_/A _12581_/B _12582_/B vssd1 vssd1 vccd1 vccd1 _12570_/B sky130_fd_sc_hd__nand3_1
XANTENNA__07798__B1 _10413_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold217 hold217/A vssd1 vssd1 vccd1 vccd1 hold217/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold206 hold206/A vssd1 vssd1 vccd1 vccd1 hold206/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold239 hold239/A vssd1 vssd1 vccd1 vccd1 hold239/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold228 hold228/A vssd1 vssd1 vccd1 vccd1 hold228/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11279__A _12073_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08800_ _08801_/A _08801_/B vssd1 vssd1 vccd1 vccd1 _08853_/A sky130_fd_sc_hd__and2_1
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13099__B2 _06572_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06992_ _06992_/A _06992_/B vssd1 vssd1 vccd1 vccd1 _06993_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_56_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09780_ _11261_/A _09780_/B vssd1 vssd1 vccd1 vccd1 _09782_/B sky130_fd_sc_hd__xnor2_2
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08731_ _08731_/A _08731_/B vssd1 vssd1 vccd1 vccd1 _08735_/A sky130_fd_sc_hd__xnor2_2
X_08662_ _08728_/A _08662_/B vssd1 vssd1 vccd1 vccd1 _08683_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_56_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07613_ _07992_/A _07992_/B vssd1 vssd1 vccd1 vccd1 _07993_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07722__B1 _10022_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12838__A _12838_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08593_ _08594_/A _08594_/B vssd1 vssd1 vccd1 vccd1 _08593_/Y sky130_fd_sc_hd__nand2_1
XANTENNA_fanout166_A _08584_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07544_ _07545_/A _07545_/B vssd1 vssd1 vccd1 vccd1 _09212_/B sky130_fd_sc_hd__and2b_1
X_07475_ _10165_/A _07475_/B vssd1 vssd1 vccd1 vccd1 _07477_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_91_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09214_ _09214_/A _09214_/B vssd1 vssd1 vccd1 vccd1 _09260_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_17_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09145_ _09137_/X _09144_/X _09974_/A vssd1 vssd1 vccd1 vccd1 _09145_/X sky130_fd_sc_hd__mux2_1
X_09076_ _12426_/B _12426_/C vssd1 vssd1 vccd1 vccd1 _09543_/A sky130_fd_sc_hd__and2_1
XFILLER_0_31_135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08027_ _08027_/A _08027_/B vssd1 vssd1 vccd1 vccd1 _08081_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_31_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08202__A1 _11564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09978_ _10119_/S _09977_/Y _09973_/X vssd1 vssd1 vccd1 vccd1 _09978_/X sky130_fd_sc_hd__a21o_1
XANTENNA__09093__S _09108_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08929_ _08929_/A _08929_/B vssd1 vssd1 vccd1 vccd1 _08930_/B sky130_fd_sc_hd__xor2_4
XANTENNA_fanout79_A _12832_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11940_ _11940_/A _11940_/B vssd1 vssd1 vccd1 vccd1 _11943_/C sky130_fd_sc_hd__or2_1
XFILLER_0_67_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11871_ _11985_/A vssd1 vssd1 vccd1 vccd1 _11872_/C sky130_fd_sc_hd__inv_2
XFILLER_0_79_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11652__A _11908_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10822_ _10971_/B _10822_/B _10822_/C vssd1 vssd1 vccd1 vccd1 _10823_/A sky130_fd_sc_hd__or3_1
X_10753_ _10752_/A _10752_/B _10752_/Y _09156_/Y vssd1 vssd1 vccd1 vccd1 _10753_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_94_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_638 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10684_ _11294_/A fanout30/X fanout27/X _10418_/A vssd1 vssd1 vccd1 vccd1 _10685_/B
+ sky130_fd_sc_hd__o22a_1
X_12423_ _12423_/A _12423_/B vssd1 vssd1 vccd1 vccd1 _12423_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_63_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11576__A1 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12354_ hold268/A _11341_/B _12396_/B _12353_/Y _09837_/A vssd1 vssd1 vccd1 vccd1
+ _12354_/X sky130_fd_sc_hd__a311o_1
XANTENNA__07244__A2 _09568_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11576__B2 fanout27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11305_ _11198_/A _11197_/B _11197_/A vssd1 vssd1 vccd1 vccd1 _11306_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_22_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12285_ _12380_/B _12285_/B vssd1 vssd1 vccd1 vccd1 _12383_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_31_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11236_ hold228/A _11236_/B vssd1 vssd1 vccd1 vccd1 _11346_/B sky130_fd_sc_hd__or2_1
XANTENNA__08744__A2 _08744_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11167_ _11168_/A _11168_/B vssd1 vssd1 vccd1 vccd1 _11292_/B sky130_fd_sc_hd__and2_1
XANTENNA__11827__A _12317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10118_ _09367_/Y _11118_/B _11118_/A vssd1 vssd1 vccd1 vccd1 _10118_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_89_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11098_ _11098_/A _11098_/B vssd1 vssd1 vccd1 vccd1 _11318_/A sky130_fd_sc_hd__and2_2
XFILLER_0_117_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10049_ fanout94/X fanout48/X _10930_/B _10941_/A vssd1 vssd1 vccd1 vccd1 _10050_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10877__S _12174_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07260_ _12076_/A _07263_/B _10928_/A vssd1 vssd1 vccd1 vccd1 _07262_/A sky130_fd_sc_hd__o21ba_1
XFILLER_0_115_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07191_ _07191_/A _07191_/B vssd1 vssd1 vccd1 vccd1 _07191_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07235__A2 _09440_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09901_ _10445_/A _10571_/B fanout51/X _10706_/B2 vssd1 vssd1 vccd1 vccd1 _09902_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10790__A2 _12150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09832_ _10391_/A2 _10120_/C hold187/A vssd1 vssd1 vccd1 vccd1 _09832_/Y sky130_fd_sc_hd__a21oi_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07155__A1_N _07149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09763_ _09764_/A _09764_/B vssd1 vssd1 vccd1 vccd1 _09763_/X sky130_fd_sc_hd__and2_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06975_ _10707_/A _06975_/B vssd1 vssd1 vccd1 vccd1 _06992_/A sky130_fd_sc_hd__xnor2_1
X_08714_ _08382_/Y _08715_/B vssd1 vssd1 vccd1 vccd1 _08714_/X sky130_fd_sc_hd__and2b_1
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09694_ _11118_/A _06939_/Y _09354_/B _06791_/B _09693_/X vssd1 vssd1 vccd1 vccd1
+ _09694_/X sky130_fd_sc_hd__o221a_1
X_08645_ _08645_/A _08645_/B vssd1 vssd1 vccd1 vccd1 _08655_/A sky130_fd_sc_hd__xnor2_2
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08576_ _08586_/A _08586_/B vssd1 vssd1 vccd1 vccd1 _08589_/B sky130_fd_sc_hd__or2_1
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11472__A _11472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07527_ _07527_/A _07527_/B vssd1 vssd1 vccd1 vccd1 _07577_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_37_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07474__A2 _09567_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07458_ _07459_/B _07459_/A vssd1 vssd1 vccd1 vccd1 _09287_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__08671__B2 _08671_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08671__A1 _08730_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11270__A3 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07389_ _07389_/A _07389_/B vssd1 vssd1 vccd1 vccd1 _07396_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_45_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09128_ _09126_/X _09127_/X _09330_/S vssd1 vssd1 vccd1 vccd1 _09128_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09088__S _09108_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_731 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09620__B1 _08752_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09059_ _09059_/A _09059_/B _12238_/A vssd1 vssd1 vccd1 vccd1 _09061_/A sky130_fd_sc_hd__or3_2
XFILLER_0_20_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12070_ fanout56/X fanout15/X fanout36/X _12316_/A vssd1 vssd1 vccd1 vccd1 _12071_/B
+ sky130_fd_sc_hd__o22a_1
X_11021_ _09527_/B _09354_/B _11021_/S vssd1 vssd1 vccd1 vccd1 _11021_/X sky130_fd_sc_hd__mux2_1
XANTENNA__11730__B2 _12254_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10533__A2 _10500_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12972_ hold185/X _13016_/A2 _13016_/B1 hold157/X vssd1 vssd1 vccd1 vccd1 hold186/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12478__A _12649_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07860__A _08740_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10297__A1 _10948_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10297__B2 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11923_ _11923_/A _12412_/B vssd1 vssd1 vccd1 vccd1 _11927_/A sky130_fd_sc_hd__or2_1
XFILLER_0_86_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11854_ _11854_/A _11854_/B vssd1 vssd1 vccd1 vccd1 _11856_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__11246__B1 _11243_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10805_ _10575_/A fanout48/X _10930_/B _10574_/A vssd1 vssd1 vccd1 vccd1 _10806_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10049__A1 fanout94/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10049__B2 _10941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12443__C1 _12455_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11785_ _11785_/A _11866_/A vssd1 vssd1 vccd1 vccd1 _11787_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_28_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10736_ _10737_/A _10737_/B vssd1 vssd1 vccd1 vccd1 _10736_/X sky130_fd_sc_hd__and2_1
XFILLER_0_12_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10667_ _10959_/A _10668_/B vssd1 vssd1 vccd1 vccd1 _10669_/B sky130_fd_sc_hd__nand2_1
X_12406_ _12400_/Y _12401_/X _12405_/X vssd1 vssd1 vccd1 vccd1 _12406_/X sky130_fd_sc_hd__o21a_1
XANTENNA__11549__B2 _09163_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07100__A _07100_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13386_ instruction[12] vssd1 vssd1 vccd1 vccd1 loadstore_dest[1] sky130_fd_sc_hd__buf_12
X_10598_ _10460_/B _10476_/B _10458_/Y vssd1 vssd1 vccd1 vccd1 _10608_/A sky130_fd_sc_hd__a21oi_2
XANTENNA__10445__B _10941_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_466 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12337_ _12287_/A _12383_/A _12287_/B _12170_/A vssd1 vssd1 vccd1 vccd1 _12337_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_10_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12268_ fanout16/X fanout8/X _12138_/A vssd1 vssd1 vccd1 vccd1 _12268_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_120_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11219_ _11218_/A _11650_/C _11707_/A vssd1 vssd1 vccd1 vccd1 _11219_/X sky130_fd_sc_hd__o21a_1
XANTENNA__11557__A _11557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12199_ _06924_/X _12186_/X _12190_/X _12198_/Y vssd1 vssd1 vccd1 vccd1 _12199_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_37_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06760_ reg1_val[7] _07080_/A vssd1 vssd1 vccd1 vccd1 _06760_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__09678__B1 _11886_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06691_ reg1_val[18] _06691_/B vssd1 vssd1 vccd1 vccd1 _06693_/B sky130_fd_sc_hd__nor2_1
XANTENNA__07153__A1 _07343_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08430_ _08798_/B2 fanout87/X fanout82/X _08646_/B2 vssd1 vssd1 vccd1 vccd1 _08431_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_53_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08350__B1 _09568_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08361_ _08436_/A _08727_/A2 _08673_/B fanout99/X vssd1 vssd1 vccd1 vccd1 _08362_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_18_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07312_ fanout30/X _09423_/B2 _12802_/A _07688_/B vssd1 vssd1 vccd1 vccd1 _07313_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_46_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08292_ _08298_/A _08298_/B _08283_/Y vssd1 vssd1 vccd1 vccd1 _08340_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_34_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07243_ _07241_/A _07241_/B _07242_/X vssd1 vssd1 vccd1 vccd1 _07269_/A sky130_fd_sc_hd__o21bai_2
XFILLER_0_61_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout129_A _10167_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07174_ _07174_/A _07174_/B vssd1 vssd1 vccd1 vccd1 _07233_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_5_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07945__A _08722_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout302 _06578_/Y vssd1 vssd1 vccd1 vccd1 _13242_/A sky130_fd_sc_hd__buf_2
XFILLER_0_111_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09905__A1 fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09905__B2 _08304_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09815_ _09653_/A _08988_/A _08988_/B _09163_/X vssd1 vssd1 vccd1 vccd1 _09815_/X
+ sky130_fd_sc_hd__a31o_1
X_06958_ _11118_/A _09974_/A _09669_/S _09336_/S vssd1 vssd1 vccd1 vccd1 _07050_/C
+ sky130_fd_sc_hd__and4_1
X_09746_ _09746_/A _09746_/B _09746_/C vssd1 vssd1 vccd1 vccd1 _09751_/A sky130_fd_sc_hd__nand3_1
XANTENNA__12268__A2 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09677_ _09675_/X _09676_/Y _09673_/X vssd1 vssd1 vccd1 vccd1 _09677_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_69_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10279__A1 fanout94/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10279__B2 _10941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06889_ _06771_/A _06589_/X _09170_/A instruction[4] _06887_/Y vssd1 vssd1 vccd1
+ vccd1 _12790_/B sky130_fd_sc_hd__a221o_1
XFILLER_0_96_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08628_ _08628_/A _08628_/B vssd1 vssd1 vccd1 vccd1 _08637_/B sky130_fd_sc_hd__xor2_2
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08559_ _08557_/Y _08577_/B _08554_/Y vssd1 vssd1 vccd1 vccd1 _08567_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_77_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08644__B2 _09598_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08644__A1 _12626_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07447__A2 _12804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11570_ _11570_/A _11570_/B vssd1 vssd1 vccd1 vccd1 _11582_/A sky130_fd_sc_hd__xor2_1
X_10521_ _06749_/Y _09158_/Y _09154_/Y vssd1 vssd1 vccd1 vccd1 _10521_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_92_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13240_ hold166/X _06892_/B _12784_/Y _06572_/A vssd1 vssd1 vccd1 vccd1 hold300/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10452_ _10452_/A _10452_/B vssd1 vssd1 vccd1 vccd1 _10454_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_17_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13171_ hold292/A _13170_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13171_/X sky130_fd_sc_hd__mux2_1
X_10383_ _10381_/Y _10383_/B vssd1 vssd1 vccd1 vccd1 _10384_/B sky130_fd_sc_hd__nand2b_1
X_12122_ _12122_/A _12122_/B vssd1 vssd1 vccd1 vccd1 _12122_/X sky130_fd_sc_hd__or2_1
XFILLER_0_20_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12053_ _12044_/Y _12045_/X _12048_/X _12052_/Y vssd1 vssd1 vccd1 vccd1 _12053_/Y
+ sky130_fd_sc_hd__o211ai_2
X_11004_ _11004_/A _11004_/B vssd1 vssd1 vccd1 vccd1 _11004_/X sky130_fd_sc_hd__or2_1
X_12955_ _13224_/B _13225_/A _12861_/X vssd1 vssd1 vccd1 vccd1 _13229_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__11467__B1 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11906_ _12210_/A _11906_/B vssd1 vssd1 vccd1 vccd1 _11908_/B sky130_fd_sc_hd__xnor2_1
X_12886_ hold279/X hold13/X vssd1 vssd1 vccd1 vccd1 _13159_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__07686__A2 _07752_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11219__B1 _11707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11837_ _07033_/A fanout6/X _11836_/X vssd1 vssd1 vccd1 vccd1 _11839_/B sky130_fd_sc_hd__o21ba_2
XANTENNA__10690__A1 fanout23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10690__B2 _11171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11768_ _11768_/A _11768_/B _11766_/X vssd1 vssd1 vccd1 vccd1 _11769_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_28_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10719_ _10601_/A _10601_/B _10604_/A vssd1 vssd1 vccd1 vccd1 _10727_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_126_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11699_ _11507_/Y _11700_/B _11700_/C vssd1 vssd1 vccd1 vccd1 _11699_/Y sky130_fd_sc_hd__o21bai_1
XANTENNA__12195__A1 _09354_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13369_ _13371_/CLK _13369_/D vssd1 vssd1 vccd1 vccd1 hold246/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07930_ _07940_/A _07940_/B vssd1 vssd1 vccd1 vccd1 _07930_/X sky130_fd_sc_hd__and2b_1
X_07861_ _07862_/A _07862_/B vssd1 vssd1 vccd1 vccd1 _07861_/Y sky130_fd_sc_hd__nor2_1
X_06812_ _06870_/C _06811_/X _06781_/X vssd1 vssd1 vccd1 vccd1 _06812_/X sky130_fd_sc_hd__a21o_1
X_09600_ _07026_/X fanout9/A fanout5/X _12802_/A vssd1 vssd1 vccd1 vccd1 _09601_/B
+ sky130_fd_sc_hd__o22a_1
X_07792_ _08742_/A _07792_/B vssd1 vssd1 vccd1 vccd1 _07881_/B sky130_fd_sc_hd__xnor2_2
X_06743_ _10644_/S _06743_/B vssd1 vssd1 vccd1 vccd1 _10629_/A sky130_fd_sc_hd__nor2_1
X_09531_ _09974_/A _11343_/B _09529_/Y _09530_/X vssd1 vssd1 vccd1 vccd1 _09531_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08596__A _08645_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08323__B1 _10022_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06674_ reg1_val[21] _07135_/D vssd1 vssd1 vccd1 vccd1 _06675_/B sky130_fd_sc_hd__and2b_1
X_09462_ _09462_/A _09462_/B vssd1 vssd1 vccd1 vccd1 _09463_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__12846__A _12846_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09393_ _09393_/A _09393_/B vssd1 vssd1 vccd1 vccd1 _09467_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__07005__A _09669_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06885__B1 _06881_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08413_ _08413_/A _08413_/B vssd1 vssd1 vccd1 vccd1 _08414_/B sky130_fd_sc_hd__and2_1
XFILLER_0_19_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08344_ _08344_/A vssd1 vssd1 vccd1 vccd1 _09028_/A sky130_fd_sc_hd__inv_2
XFILLER_0_74_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08275_ _08275_/A _08275_/B vssd1 vssd1 vccd1 vccd1 _08332_/A sky130_fd_sc_hd__xor2_1
X_07226_ _07226_/A _07226_/B vssd1 vssd1 vccd1 vccd1 _07226_/X sky130_fd_sc_hd__and2_1
Xclkbuf_4_1_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13371_/CLK sky130_fd_sc_hd__clkbuf_8
X_07157_ reg1_val[4] _07160_/B _07200_/A vssd1 vssd1 vccd1 vccd1 _07159_/B sky130_fd_sc_hd__o21a_2
XFILLER_0_100_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07088_ _06964_/A _06964_/B _07074_/B vssd1 vssd1 vccd1 vccd1 _07089_/B sky130_fd_sc_hd__o21a_1
Xfanout121 _08432_/B vssd1 vssd1 vccd1 vccd1 _10706_/B2 sky130_fd_sc_hd__clkbuf_8
Xfanout110 _07009_/X vssd1 vssd1 vccd1 vccd1 _09716_/A sky130_fd_sc_hd__buf_8
Xfanout165 _08979_/X vssd1 vssd1 vccd1 vccd1 _10391_/A2 sky130_fd_sc_hd__buf_4
Xfanout154 _06946_/X vssd1 vssd1 vccd1 vccd1 _08722_/A sky130_fd_sc_hd__buf_12
Xfanout132 _07189_/X vssd1 vssd1 vccd1 vccd1 _09567_/B sky130_fd_sc_hd__buf_8
Xfanout143 _12802_/A vssd1 vssd1 vccd1 vccd1 _07955_/A sky130_fd_sc_hd__buf_6
Xfanout198 _12791_/Y vssd1 vssd1 vccd1 vccd1 _13077_/A2 sky130_fd_sc_hd__buf_2
Xfanout187 _09431_/A vssd1 vssd1 vccd1 vccd1 _08740_/A sky130_fd_sc_hd__buf_12
XANTENNA__08562__B1 _09568_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout176 _09444_/A vssd1 vssd1 vccd1 vccd1 _08727_/A2 sky130_fd_sc_hd__clkbuf_8
XANTENNA__11925__A _12317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11161__A2 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09729_ _09730_/A _09730_/B vssd1 vssd1 vccd1 vccd1 _09869_/A sky130_fd_sc_hd__nor2_1
XANTENNA_fanout61_A _12214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06738__B _06799_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12740_ _12737_/A _12739_/B _12737_/B vssd1 vssd1 vccd1 vccd1 _12742_/A sky130_fd_sc_hd__a21bo_1
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12671_ _12671_/A _12671_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[9] sky130_fd_sc_hd__xor2_4
XFILLER_0_127_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11622_ _11623_/B _11623_/C _11623_/A vssd1 vssd1 vccd1 vccd1 _11624_/B sky130_fd_sc_hd__a21oi_1
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11660__A _11751_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11248__A1_N _12254_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11553_ _11361_/B _11428_/Y _11518_/Y _11874_/A vssd1 vssd1 vccd1 vccd1 _11614_/A
+ sky130_fd_sc_hd__o31a_1
XANTENNA__08093__A2 _08744_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10504_ _10748_/A _10503_/B _10503_/C vssd1 vssd1 vccd1 vccd1 _10504_/Y sky130_fd_sc_hd__o21ai_1
X_11484_ fanout27/X _11989_/A _11923_/A fanout29/X vssd1 vssd1 vccd1 vccd1 _11485_/B
+ sky130_fd_sc_hd__o22a_1
X_13223_ _13235_/A hold267/X vssd1 vssd1 vccd1 vccd1 _13375_/D sky130_fd_sc_hd__and2_1
XANTENNA__12491__A _12659_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10435_ _10959_/A _10435_/B vssd1 vssd1 vccd1 vccd1 _10439_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__10188__B1 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13154_ _12887_/X _13154_/B vssd1 vssd1 vccd1 vccd1 _13155_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_110_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07053__B1 _12802_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11924__A1 _12150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11924__B2 _12213_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12105_ _12031_/B _12031_/C _12031_/A vssd1 vssd1 vccd1 vccd1 _12106_/B sky130_fd_sc_hd__a21oi_1
X_10366_ _10617_/A _10741_/A vssd1 vssd1 vccd1 vccd1 _10366_/Y sky130_fd_sc_hd__nor2_1
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13085_ _07508_/B _12798_/B hold84/X vssd1 vssd1 vccd1 vccd1 hold85/A sky130_fd_sc_hd__a21oi_1
XANTENNA__06800__B1 _06799_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10297_ _10948_/B2 _12214_/A fanout51/X fanout74/X vssd1 vssd1 vccd1 vccd1 _10298_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_20_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12036_ _06648_/D _12034_/X _12035_/Y vssd1 vssd1 vccd1 vccd1 _12036_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_18_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11152__A2 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11835__A _12073_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07108__B2 _09423_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07108__A1 fanout30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12938_ hold293/A hold15/X vssd1 vssd1 vccd1 vccd1 _12939_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_87_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07659__A2 _10574_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12869_ hold41/X hold254/X vssd1 vssd1 vccd1 vccd1 _12869_/X sky130_fd_sc_hd__and2b_1
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13062__C1 _13128_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08060_ _08060_/A _08060_/B vssd1 vssd1 vccd1 vccd1 _08067_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_114_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07011_ _09716_/A _07013_/B vssd1 vssd1 vccd1 vccd1 _07017_/A sky130_fd_sc_hd__and2_1
XFILLER_0_12_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08962_ _08962_/A _08962_/B vssd1 vssd1 vccd1 vccd1 _08965_/B sky130_fd_sc_hd__xor2_2
X_08893_ _08893_/A _08893_/B vssd1 vssd1 vccd1 vccd1 _08895_/B sky130_fd_sc_hd__xnor2_1
X_07913_ _07913_/A _07913_/B _07913_/C vssd1 vssd1 vccd1 vccd1 _07916_/A sky130_fd_sc_hd__and3_1
XANTENNA_fanout196_A _07220_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11143__A2 _10871_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07844_ _07816_/A _07816_/C _07816_/B vssd1 vssd1 vccd1 vccd1 _07846_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07775_ _07776_/A _07776_/B vssd1 vssd1 vccd1 vccd1 _07781_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_91_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09514_ reg1_val[2] curr_PC[2] vssd1 vssd1 vccd1 vccd1 _09514_/Y sky130_fd_sc_hd__nor2_1
X_06726_ reg2_val[12] _06799_/B vssd1 vssd1 vccd1 vccd1 _06726_/X sky130_fd_sc_hd__and2_1
XANTENNA__10103__B1 _11707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06657_ _06686_/A _12659_/B vssd1 vssd1 vccd1 vccd1 _06657_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_78_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09445_ _09445_/A _09445_/B vssd1 vssd1 vccd1 vccd1 _09446_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__10654__A1 _11876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13171__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06588_ instruction[1] instruction[2] instruction[0] pred_val vssd1 vssd1 vccd1 vccd1
+ _06897_/B sky130_fd_sc_hd__and4bb_2
XFILLER_0_74_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09376_ _09542_/A _09543_/A _09542_/B _12426_/A vssd1 vssd1 vccd1 vccd1 _09376_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__10406__A1 _11142_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06574__A _12626_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10096__A _10096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08327_ _08327_/A _08327_/B vssd1 vssd1 vccd1 vccd1 _08349_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_117_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07283__B1 _10570_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08258_ _08752_/A fanout75/X _08304_/B _08798_/B2 vssd1 vssd1 vccd1 vccd1 _08259_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_7_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_758 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07209_ _07131_/B _06961_/Y _06966_/Y _07129_/X _07223_/B vssd1 vssd1 vccd1 vccd1
+ _07210_/B sky130_fd_sc_hd__a41o_1
XFILLER_0_61_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09096__S _09108_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10220_ _10220_/A _10220_/B vssd1 vssd1 vccd1 vccd1 _10221_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_15_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08189_ _08189_/A _08242_/A vssd1 vssd1 vccd1 vccd1 _08200_/B sky130_fd_sc_hd__and2_1
XFILLER_0_30_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10151_ _10928_/A _10151_/B vssd1 vssd1 vccd1 vccd1 _10155_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__11382__A2 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10082_ _09885_/A _09885_/B _09883_/Y vssd1 vssd1 vccd1 vccd1 _10085_/A sky130_fd_sc_hd__a21boi_2
XANTENNA__08535__B1 _08564_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10984_ _10985_/B _10985_/A vssd1 vssd1 vccd1 vccd1 _11097_/B sky130_fd_sc_hd__and2b_1
XANTENNA__10645__A1 _12307_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12723_ _12723_/A _12725_/D vssd1 vssd1 vccd1 vccd1 loadstore_address[19] sky130_fd_sc_hd__xnor2_4
XFILLER_0_29_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12654_ reg1_val[6] _12654_/B vssd1 vssd1 vccd1 vccd1 _12655_/B sky130_fd_sc_hd__and2_1
XFILLER_0_127_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12585_ _12595_/A _12585_/B vssd1 vssd1 vccd1 vccd1 new_PC[20] sky130_fd_sc_hd__xnor2_4
XFILLER_0_65_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11605_ _11511_/A _11507_/Y _11509_/B vssd1 vssd1 vccd1 vccd1 _11605_/Y sky130_fd_sc_hd__o21ai_2
X_11536_ hold277/A hold292/A _11536_/C vssd1 vssd1 vccd1 vccd1 _11635_/B sky130_fd_sc_hd__or3_1
XFILLER_0_53_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10948__A2 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13206_ _12869_/X _13206_/B vssd1 vssd1 vccd1 vccd1 _13207_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_110_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11467_ _09613_/A _12213_/A fanout56/X _09614_/A vssd1 vssd1 vccd1 vccd1 _11468_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_0_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11398_ _11398_/A _11398_/B vssd1 vssd1 vccd1 vccd1 _11412_/A sky130_fd_sc_hd__xnor2_2
X_10418_ _10418_/A _11171_/A vssd1 vssd1 vccd1 vccd1 _10419_/C sky130_fd_sc_hd__or2_1
XFILLER_0_29_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13137_ hold269/X _12789_/B _13136_/X _12790_/A vssd1 vssd1 vccd1 vccd1 hold270/A
+ sky130_fd_sc_hd__a22o_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10349_ _10178_/A _10178_/C _10178_/B vssd1 vssd1 vccd1 vccd1 _10352_/A sky130_fd_sc_hd__o21ba_1
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13068_ hold123/X _12791_/A _13080_/B1 hold116/X _13113_/A vssd1 vssd1 vccd1 vccd1
+ hold127/A sky130_fd_sc_hd__o221a_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10581__B1 _10930_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12019_ _12017_/X _12019_/B vssd1 vssd1 vccd1 vccd1 _12162_/A sky130_fd_sc_hd__nand2b_2
XFILLER_0_29_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10396__A1_N _07089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07560_ _07560_/A _07560_/B vssd1 vssd1 vccd1 vccd1 _07597_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_45_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07491_ _07491_/A _07491_/B vssd1 vssd1 vccd1 vccd1 _07492_/B sky130_fd_sc_hd__nand2_1
X_09230_ _09231_/A _09231_/B vssd1 vssd1 vccd1 vccd1 _09232_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_48_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09161_ _12403_/A1 _09160_/X _06865_/Y vssd1 vssd1 vccd1 vccd1 _09161_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__13050__A2 _12788_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09092_ reg1_val[7] reg1_val[24] _09108_/S vssd1 vssd1 vccd1 vccd1 _09092_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_43_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08112_ _10537_/A1 _08723_/B1 _07885_/B _08432_/B vssd1 vssd1 vccd1 vccd1 _08113_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_28_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08043_ _08727_/A2 _11472_/A _11558_/A _08727_/B1 vssd1 vssd1 vccd1 vccd1 _08044_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__06841__B _07140_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout111_A _12076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10363__B _10364_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09994_ _09156_/Y _09964_/X _09968_/Y _09111_/S _09993_/X vssd1 vssd1 vccd1 vccd1
+ _09994_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_86_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12313__A1 _07343_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08945_ _08930_/A _08930_/B _08928_/Y vssd1 vssd1 vccd1 vccd1 _08946_/B sky130_fd_sc_hd__a21oi_2
X_08876_ _08876_/A _08876_/B vssd1 vssd1 vccd1 vccd1 _08878_/B sky130_fd_sc_hd__xor2_2
X_07827_ _11385_/A _07827_/B vssd1 vssd1 vccd1 vccd1 _07831_/A sky130_fd_sc_hd__xnor2_1
X_07758_ _12073_/A _07758_/B vssd1 vssd1 vccd1 vccd1 _07759_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_94_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06709_ _06805_/A _06587_/X _06686_/A _06708_/X vssd1 vssd1 vccd1 vccd1 _06988_/A
+ sky130_fd_sc_hd__a31o_4
XFILLER_0_109_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07689_ _11673_/A _07689_/B vssd1 vssd1 vccd1 vccd1 _07691_/B sky130_fd_sc_hd__xnor2_1
X_09428_ _09428_/A _09428_/B vssd1 vssd1 vccd1 vccd1 _09429_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_66_269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09359_ _09523_/A _09154_/Y _09346_/X _12394_/A vssd1 vssd1 vccd1 vccd1 _09359_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_19_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08048__A2 _09614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12370_ _12372_/B vssd1 vssd1 vccd1 vccd1 _12371_/B sky130_fd_sc_hd__inv_2
XFILLER_0_34_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11052__B2 _10574_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11052__A1 _10575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11321_ _10868_/A _11320_/Y _11319_/Y _11317_/Y vssd1 vssd1 vccd1 vccd1 _11321_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_35_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06751__B _06799_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11252_ curr_PC[15] _11253_/B vssd1 vssd1 vccd1 vccd1 _11252_/X sky130_fd_sc_hd__or2_1
XFILLER_0_30_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11183_ _11183_/A _11183_/B vssd1 vssd1 vccd1 vccd1 _11184_/B sky130_fd_sc_hd__or2_1
X_10203_ _10205_/A _10205_/B vssd1 vssd1 vccd1 vccd1 _10206_/A sky130_fd_sc_hd__and2_1
XFILLER_0_101_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10134_ _12244_/S _09172_/B _10133_/Y _10128_/X _10123_/Y vssd1 vssd1 vccd1 vccd1
+ _10134_/X sky130_fd_sc_hd__a311o_1
XANTENNA__08220__A2 _08744_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11385__A _11385_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10065_ _11172_/A _10065_/B vssd1 vssd1 vccd1 vccd1 _10069_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09720__A2 _10413_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07731__B2 _08732_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07731__A1 _08741_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_79 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10967_ _10967_/A _10967_/B _10967_/C vssd1 vssd1 vccd1 vccd1 _10969_/A sky130_fd_sc_hd__and3_1
XFILLER_0_127_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10898_ _12307_/B1 _10897_/X _06731_/B vssd1 vssd1 vccd1 vccd1 _10898_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__07495__B1 _09440_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12706_ _12706_/A _12706_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[15] sky130_fd_sc_hd__nor2_8
XFILLER_0_38_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09236__A1 _09444_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07103__A _11269_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12637_ _12636_/A _12633_/Y _12635_/B vssd1 vssd1 vccd1 vccd1 _12641_/A sky130_fd_sc_hd__o21a_2
XANTENNA__13032__A2 _06572_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09236__B2 _09236_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11043__A1 _10448_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12568_ _12581_/B _12582_/B _12581_/A vssd1 vssd1 vccd1 vccd1 _12575_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_80_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12663__B _12664_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold207 hold207/A vssd1 vssd1 vccd1 vccd1 hold207/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12499_ _12664_/B _12499_/B vssd1 vssd1 vccd1 vccd1 _12500_/B sky130_fd_sc_hd__or2_1
XFILLER_0_80_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11519_ _11519_/A _11649_/C vssd1 vssd1 vccd1 vccd1 _11519_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__10464__A _11269_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold218 hold218/A vssd1 vssd1 vccd1 vccd1 hold218/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold229 hold229/A vssd1 vssd1 vccd1 vccd1 hold229/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10003__C1 _10959_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13099__A2 _06892_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06773__A2 _06771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06991_ _06992_/A _06992_/B vssd1 vssd1 vccd1 vccd1 _07374_/A sky130_fd_sc_hd__or2_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10306__B1 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08730_ _08730_/A1 _08038_/B _08038_/C _08038_/A _11558_/A vssd1 vssd1 vccd1 vccd1
+ _08731_/B sky130_fd_sc_hd__o32a_1
X_08661_ _08673_/A _08661_/A2 _08673_/B _08671_/B2 vssd1 vssd1 vccd1 vccd1 _08662_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_56_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07722__A1 _10927_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07612_ _11269_/A _07612_/B vssd1 vssd1 vccd1 vccd1 _07992_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07722__B2 _11367_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08592_ _08613_/A _08592_/B vssd1 vssd1 vccd1 vccd1 _08594_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_76_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07543_ _10422_/A _07543_/B vssd1 vssd1 vccd1 vccd1 _07545_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__13015__A _13214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07474_ _12844_/A _09567_/B _09568_/B _12846_/A vssd1 vssd1 vccd1 vccd1 _07475_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_119_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09213_ _09211_/X _09213_/B vssd1 vssd1 vccd1 vccd1 _09214_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_17_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07013__A _11172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12854__A _12854_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09144_ _09140_/X _09143_/X _09663_/S vssd1 vssd1 vccd1 vccd1 _09144_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_72_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12231__B1 _11707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09075_ _09075_/A _09075_/B vssd1 vssd1 vccd1 vccd1 _12426_/C sky130_fd_sc_hd__xnor2_2
XFILLER_0_4_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1 fanout2/X vssd1 vssd1 vccd1 vccd1 fanout1/X sky130_fd_sc_hd__clkbuf_8
X_08026_ _08026_/A _08026_/B vssd1 vssd1 vccd1 vccd1 _08081_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_31_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09977_ _11010_/S _09975_/Y _09976_/X vssd1 vssd1 vccd1 vccd1 _09977_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__07410__B1 _10948_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08928_ _08929_/A _08929_/B vssd1 vssd1 vccd1 vccd1 _08928_/Y sky130_fd_sc_hd__nor2_1
X_08859_ _08859_/A _08859_/B vssd1 vssd1 vccd1 vccd1 _08861_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__13247__C1 _13242_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11870_ _12165_/A _11870_/B vssd1 vssd1 vccd1 vccd1 _11985_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_39_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10821_ _10821_/A _10821_/B vssd1 vssd1 vccd1 vccd1 _10822_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_109_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10752_ _10752_/A _10752_/B vssd1 vssd1 vccd1 vccd1 _10752_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_55_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12422_ _12389_/A _12387_/X _12423_/A _12402_/S vssd1 vssd1 vccd1 vccd1 _12422_/X
+ sky130_fd_sc_hd__a211o_1
X_10683_ _10695_/B vssd1 vssd1 vccd1 vccd1 _10683_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_62_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07858__A _08742_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12353_ _11341_/B _12396_/B hold268/A vssd1 vssd1 vccd1 vccd1 _12353_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_50_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11576__A2 _11989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12284_ _12161_/Y _12281_/B _12282_/Y _12028_/B _12283_/Y vssd1 vssd1 vccd1 vccd1
+ _12285_/B sky130_fd_sc_hd__o221a_1
XANTENNA__10784__B1 _10941_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11304_ _11304_/A _11304_/B vssd1 vssd1 vccd1 vccd1 _11306_/A sky130_fd_sc_hd__nand2_1
X_11235_ _11886_/A _11230_/Y _11234_/Y _09172_/B vssd1 vssd1 vccd1 vccd1 _11250_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_31_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11166_ _11470_/A _11166_/B vssd1 vssd1 vccd1 vccd1 _11168_/B sky130_fd_sc_hd__xnor2_1
Xclkbuf_4_14_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13383_/CLK sky130_fd_sc_hd__clkbuf_8
X_10117_ _09505_/X _09508_/X _10250_/S vssd1 vssd1 vccd1 vccd1 _11118_/B sky130_fd_sc_hd__mux2_1
X_11097_ _11097_/A _11097_/B _11097_/C vssd1 vssd1 vccd1 vccd1 _11098_/B sky130_fd_sc_hd__or3_1
X_10048_ _09864_/B _09867_/B _09864_/A vssd1 vssd1 vccd1 vccd1 _10059_/A sky130_fd_sc_hd__o21ba_1
XFILLER_0_26_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold90 hold90/A vssd1 vssd1 vccd1 vccd1 hold90/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12658__B _12659_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11999_ fanout29/X _12316_/A fanout12/X fanout27/X vssd1 vssd1 vccd1 vccd1 _12000_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_85_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07190_ _07220_/C _07134_/Y _07074_/B vssd1 vssd1 vccd1 vccd1 _07191_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_54_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07640__B1 _12802_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09900_ _09900_/A _09900_/B vssd1 vssd1 vccd1 vccd1 _09913_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_111_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09831_ hold234/A hold238/A hold248/A hold290/A vssd1 vssd1 vccd1 vccd1 _10120_/C
+ sky130_fd_sc_hd__or4_2
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06974_ _10445_/A _12826_/A _10706_/B2 _10418_/A vssd1 vssd1 vccd1 vccd1 _06975_/B
+ sky130_fd_sc_hd__o22a_1
X_09762_ _09889_/A _09762_/B vssd1 vssd1 vccd1 vccd1 _09764_/B sky130_fd_sc_hd__or2_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12819__A2 _12818_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08713_ _08425_/X _08715_/B _08382_/Y vssd1 vssd1 vccd1 vccd1 _08713_/Y sky130_fd_sc_hd__a21oi_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09693_ hold284/A _09691_/X _09692_/Y vssd1 vssd1 vccd1 vccd1 _09693_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08644_ _12626_/A _08632_/A _08632_/B _08632_/C _09598_/A vssd1 vssd1 vccd1 vccd1
+ _08645_/B sky130_fd_sc_hd__a32o_1
XFILLER_0_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08575_ _08575_/A _08575_/B vssd1 vssd1 vccd1 vccd1 _08586_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_49_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11472__B _12214_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07526_ _07526_/A _07526_/B vssd1 vssd1 vccd1 vccd1 _07527_/B sky130_fd_sc_hd__nor2_1
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07457_ _09287_/A _07457_/B vssd1 vssd1 vccd1 vccd1 _07459_/B sky130_fd_sc_hd__nand2_2
XANTENNA__08671__A2 _07821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07388_ _07281_/A _07281_/B _07277_/Y vssd1 vssd1 vccd1 vccd1 _07396_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_51_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09127_ reg1_val[15] reg1_val[16] _09127_/S vssd1 vssd1 vccd1 vccd1 _09127_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_60_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09620__A1 _11065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09058_ _09058_/A _09058_/B vssd1 vssd1 vccd1 vccd1 _12238_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_60_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09620__B2 _11146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08009_ _07784_/A _07784_/B _07745_/Y vssd1 vssd1 vccd1 vccd1 _08019_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_32_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout91_A _11564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11020_ _11020_/A _12404_/A vssd1 vssd1 vccd1 vccd1 _11020_/Y sky130_fd_sc_hd__nand2_1
X_12971_ _13009_/A hold188/X vssd1 vssd1 vccd1 vccd1 _13288_/D sky130_fd_sc_hd__and2_1
XFILLER_0_99_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07698__B1 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10297__A2 _12214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11922_ _12261_/A _11922_/B vssd1 vssd1 vccd1 vccd1 _11929_/A sky130_fd_sc_hd__xnor2_1
X_11853_ _11853_/A _11853_/B vssd1 vssd1 vccd1 vccd1 _11854_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__11246__A1 _06988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10804_ _10814_/B vssd1 vssd1 vccd1 vccd1 _10804_/Y sky130_fd_sc_hd__inv_2
XANTENNA__10049__A2 fanout48/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11784_ _11700_/B _11696_/Y _11698_/B vssd1 vssd1 vccd1 vccd1 _11784_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_125_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10735_ _10737_/A _10737_/B vssd1 vssd1 vccd1 vccd1 _10735_/X sky130_fd_sc_hd__or2_1
X_10666_ _10963_/A _10797_/B fanout4/X _10818_/A vssd1 vssd1 vccd1 vccd1 _10668_/B
+ sky130_fd_sc_hd__o22ai_1
XANTENNA__07870__B1 _11923_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12405_ _09127_/S _09341_/Y _12394_/B _09153_/Y _12404_/Y vssd1 vssd1 vccd1 vccd1
+ _12405_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_36_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13385_ instruction[11] vssd1 vssd1 vccd1 vccd1 loadstore_dest[0] sky130_fd_sc_hd__buf_12
XFILLER_0_106_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11954__C1 _11876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10597_ _10597_/A _10597_/B vssd1 vssd1 vccd1 vccd1 _10611_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_105_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06976__A2 _06994_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12336_ _12413_/A _12336_/B vssd1 vssd1 vccd1 vccd1 _12383_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_23_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06653__A_N _07194_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12267_ _12325_/B _12267_/B vssd1 vssd1 vccd1 vccd1 _12271_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_121_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12198_ _09111_/S _09978_/X _12194_/Y _12197_/Y vssd1 vssd1 vccd1 vccd1 _12198_/Y
+ sky130_fd_sc_hd__a211oi_1
X_11218_ _11218_/A _11650_/C vssd1 vssd1 vccd1 vccd1 _11218_/Y sky130_fd_sc_hd__nand2_1
X_11149_ _11150_/A _11150_/B vssd1 vssd1 vccd1 vccd1 _11303_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_128_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06690_ reg1_val[18] _06691_/B vssd1 vssd1 vccd1 vccd1 _11540_/A sky130_fd_sc_hd__and2_1
XFILLER_0_53_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08350__A1 _09768_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08350__B2 _07885_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08360_ _08364_/A _08364_/B vssd1 vssd1 vccd1 vccd1 _08360_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__10189__A _11163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07311_ _07269_/A _07269_/B _07268_/A vssd1 vssd1 vccd1 vccd1 _07325_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_53_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08291_ _08291_/A _08291_/B vssd1 vssd1 vccd1 vccd1 _08298_/B sky130_fd_sc_hd__xor2_1
X_07242_ _07302_/A _07302_/B vssd1 vssd1 vccd1 vccd1 _07242_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_6_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07173_ _07173_/A _07173_/B vssd1 vssd1 vccd1 vccd1 _07174_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_42_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13162__B2 _13246_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout303 _06577_/Y vssd1 vssd1 vccd1 vccd1 _12174_/S sky130_fd_sc_hd__clkbuf_8
XANTENNA__09218__A _10165_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09905__A2 _11847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09814_ _09653_/A _08988_/A _08988_/B vssd1 vssd1 vccd1 vccd1 _09814_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__11173__B1 _11172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06957_ _12341_/A _07064_/B vssd1 vssd1 vccd1 vccd1 _07223_/B sky130_fd_sc_hd__nand2_8
X_09745_ _09745_/A _09745_/B vssd1 vssd1 vccd1 vccd1 _09746_/C sky130_fd_sc_hd__or2_1
XTAP_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06888_ _06771_/A _06589_/X _09170_/A instruction[4] _06887_/Y vssd1 vssd1 vccd1
+ vccd1 _12791_/B sky130_fd_sc_hd__a221oi_4
XANTENNA__06577__A _12341_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09676_ reg1_val[3] curr_PC[3] vssd1 vssd1 vccd1 vccd1 _09676_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__10279__A2 _10571_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11483__A _12261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08627_ _08627_/A _08627_/B vssd1 vssd1 vccd1 vccd1 _08637_/A sky130_fd_sc_hd__xor2_2
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08558_ _08558_/A _08558_/B vssd1 vssd1 vccd1 vccd1 _08577_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_77_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08644__A2 _08632_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08489_ _08489_/A _08489_/B _08489_/C vssd1 vssd1 vccd1 vccd1 _08491_/B sky130_fd_sc_hd__nor3_1
X_07509_ _12138_/A _12316_/B _07508_/B vssd1 vssd1 vccd1 vccd1 _12366_/B sky130_fd_sc_hd__or3b_2
XFILLER_0_37_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10520_ hold232/A _11633_/B _10641_/B _11968_/B1 vssd1 vssd1 vccd1 vccd1 _10520_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__09400__B _10818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10451_ _10449_/X _10451_/B vssd1 vssd1 vccd1 vccd1 _10452_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_60_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13170_ _13170_/A _13170_/B vssd1 vssd1 vccd1 vccd1 _13170_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__09827__S _11118_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10382_ reg1_val[8] curr_PC[8] vssd1 vssd1 vccd1 vccd1 _10383_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_60_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12121_ hold261/A _11636_/B _12187_/B _12247_/C1 vssd1 vssd1 vccd1 vccd1 _12122_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_32_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12052_ _09111_/S _10252_/X _12051_/X vssd1 vssd1 vccd1 vccd1 _12052_/Y sky130_fd_sc_hd__a21oi_1
X_11003_ _11004_/A _11004_/B vssd1 vssd1 vccd1 vccd1 _11003_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__07871__A _08731_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12954_ _13220_/A _12953_/B _12863_/X vssd1 vssd1 vccd1 vccd1 _13225_/A sky130_fd_sc_hd__a21o_1
XANTENNA__11467__B2 _09614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11467__A1 _09613_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11905_ fanout29/X fanout56/X _12316_/A fanout27/X vssd1 vssd1 vccd1 vccd1 _11906_/B
+ sky130_fd_sc_hd__o22a_1
X_12885_ hold13/X hold279/X vssd1 vssd1 vccd1 vccd1 _12885_/X sky130_fd_sc_hd__and2b_1
XTAP_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11836_ _11261_/A _07037_/B fanout6/X _11180_/A vssd1 vssd1 vccd1 vccd1 _11836_/X
+ sky130_fd_sc_hd__o31a_1
XANTENNA__10690__A2 _09745_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11767_ _11768_/A _11768_/B _11766_/X vssd1 vssd1 vccd1 vccd1 _11767_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_28_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10718_ _10597_/A _10597_/B _10595_/Y vssd1 vssd1 vccd1 vccd1 _10729_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_70_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07111__A _11987_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11698_ _11698_/A _11698_/B vssd1 vssd1 vccd1 vccd1 _11866_/A sky130_fd_sc_hd__and2_1
X_10649_ _07100_/A _12404_/A _10645_/Y vssd1 vssd1 vccd1 vccd1 _10649_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_82_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13368_ _13371_/CLK _13368_/D vssd1 vssd1 vccd1 vccd1 hold252/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12319_ _12319_/A _12319_/B vssd1 vssd1 vccd1 vccd1 _12320_/B sky130_fd_sc_hd__and2_1
X_13299_ _13299_/CLK _13299_/D vssd1 vssd1 vccd1 vccd1 hold174/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07860_ _08740_/A _07860_/B vssd1 vssd1 vccd1 vccd1 _07862_/B sky130_fd_sc_hd__xnor2_1
X_06811_ _09686_/B _06810_/X _06788_/X vssd1 vssd1 vccd1 vccd1 _06811_/X sky130_fd_sc_hd__a21o_1
X_07791_ _11367_/A _08741_/A2 _08617_/B _11472_/A vssd1 vssd1 vccd1 vccd1 _07792_/B
+ sky130_fd_sc_hd__o22a_1
X_06742_ reg1_val[10] _07100_/A vssd1 vssd1 vccd1 vccd1 _06743_/B sky130_fd_sc_hd__nor2_1
X_09530_ hold240/A _09835_/B _09528_/X _09837_/A vssd1 vssd1 vccd1 vccd1 _09530_/X
+ sky130_fd_sc_hd__a31o_1
X_09461_ _09462_/A _09462_/B vssd1 vssd1 vccd1 vccd1 _09461_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__08323__A1 _07896_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08323__B2 _08723_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06673_ _07135_/D reg1_val[21] vssd1 vssd1 vccd1 vccd1 _11811_/S sky130_fd_sc_hd__and2b_1
XFILLER_0_93_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09392_ _09393_/B _09393_/A vssd1 vssd1 vccd1 vccd1 _09392_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_80_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08412_ _08443_/A _08443_/B vssd1 vssd1 vccd1 vccd1 _08444_/A sky130_fd_sc_hd__or2_1
XFILLER_0_59_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout141_A _12808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08343_ _08343_/A _08343_/B vssd1 vssd1 vccd1 vccd1 _08344_/A sky130_fd_sc_hd__xor2_1
XANTENNA__13023__A _13214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08274_ _08742_/A _08274_/B vssd1 vssd1 vccd1 vccd1 _08275_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_116_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07225_ _07074_/B _07220_/C _07223_/Y _07135_/D vssd1 vssd1 vccd1 vccd1 _07226_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_46_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08117__A _08724_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07156_ _08645_/A _07156_/B vssd1 vssd1 vccd1 vccd1 _07173_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07956__A _11564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07087_ _07087_/A _07087_/B vssd1 vssd1 vccd1 vccd1 _07087_/X sky130_fd_sc_hd__or2_4
Xfanout122 _06971_/Y vssd1 vssd1 vccd1 vccd1 _08432_/B sky130_fd_sc_hd__buf_6
Xfanout111 _12076_/A vssd1 vssd1 vccd1 vccd1 _12210_/A sky130_fd_sc_hd__clkbuf_16
Xfanout100 _11385_/A vssd1 vssd1 vccd1 vccd1 _11470_/A sky130_fd_sc_hd__clkbuf_16
Xfanout133 _09238_/B vssd1 vssd1 vccd1 vccd1 _08732_/A2 sky130_fd_sc_hd__buf_6
Xfanout144 _09766_/A vssd1 vssd1 vccd1 vccd1 _12802_/A sky130_fd_sc_hd__buf_8
Xfanout155 _12031_/A vssd1 vssd1 vccd1 vccd1 _11792_/A sky130_fd_sc_hd__buf_4
Xfanout199 _12790_/Y vssd1 vssd1 vccd1 vccd1 _12848_/B sky130_fd_sc_hd__buf_4
Xfanout188 _09153_/Y vssd1 vssd1 vccd1 vccd1 _12254_/A1 sky130_fd_sc_hd__buf_4
XANTENNA__08562__B2 _08646_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08562__A1 _08798_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout177 _09444_/A vssd1 vssd1 vccd1 vccd1 _08661_/A2 sky130_fd_sc_hd__clkbuf_4
Xfanout166 _08584_/A vssd1 vssd1 vccd1 vccd1 _08745_/A sky130_fd_sc_hd__clkbuf_16
X_09728_ _09575_/B _09578_/B _09575_/A vssd1 vssd1 vccd1 vccd1 _09730_/B sky130_fd_sc_hd__o21ba_1
X_07989_ _07989_/A _07989_/B vssd1 vssd1 vccd1 vccd1 _08008_/A sky130_fd_sc_hd__xnor2_2
XANTENNA_fanout54_A _12842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09659_ _09312_/X _09315_/X _09666_/S vssd1 vssd1 vccd1 vccd1 _09659_/X sky130_fd_sc_hd__mux2_1
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12670_ _12675_/B _12677_/A vssd1 vssd1 vccd1 vccd1 _12671_/B sky130_fd_sc_hd__nand2_2
X_11621_ _12423_/A _11621_/B vssd1 vssd1 vccd1 vccd1 _11623_/C sky130_fd_sc_hd__or2_1
XFILLER_0_77_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09411__A _09411_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11660__B _12261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06754__B _07089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11552_ _11142_/S _11549_/X _11734_/C _11551_/Y vssd1 vssd1 vccd1 vccd1 dest_val[18]
+ sky130_fd_sc_hd__o22ai_4
XFILLER_0_52_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10503_ _10748_/A _10503_/B _10503_/C vssd1 vssd1 vccd1 vccd1 _10503_/X sky130_fd_sc_hd__or3_1
XFILLER_0_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11483_ _12261_/A _11483_/B vssd1 vssd1 vccd1 vccd1 _11486_/A sky130_fd_sc_hd__xnor2_1
X_13222_ hold266/X _12789_/B _13221_/X _12790_/A vssd1 vssd1 vccd1 vccd1 hold267/A
+ sky130_fd_sc_hd__a22o_1
X_10434_ _10664_/A _10797_/B fanout5/X _10567_/A vssd1 vssd1 vccd1 vccd1 _10435_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10188__A1 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13153_ _13245_/A hold283/X vssd1 vssd1 vccd1 vccd1 _13360_/D sky130_fd_sc_hd__and2_1
XFILLER_0_60_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10365_ _10094_/X _10229_/X _10230_/X vssd1 vssd1 vccd1 vccd1 _10365_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__07053__B2 _11171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07053__A1 _09423_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11924__A2 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10188__B2 _10948_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12104_ _12103_/A _12103_/B _12290_/A vssd1 vssd1 vccd1 vccd1 _12104_/X sky130_fd_sc_hd__a21o_1
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13084_ hold83/X _06572_/A _06892_/B _06566_/Y rst vssd1 vssd1 vccd1 vccd1 hold84/A
+ sky130_fd_sc_hd__a221o_1
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10296_ _10448_/A _10296_/B vssd1 vssd1 vccd1 vccd1 _10413_/C sky130_fd_sc_hd__xnor2_1
X_12035_ _06648_/D _12034_/X _11624_/A vssd1 vssd1 vccd1 vccd1 _12035_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_18_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07108__A2 _12798_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12937_ _13179_/B _13180_/A _12878_/X vssd1 vssd1 vccd1 vccd1 _13184_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_88_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12868_ _12866_/X _12868_/B vssd1 vssd1 vccd1 vccd1 _13211_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__06945__A _07200_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11819_ curr_PC[21] _11819_/B vssd1 vssd1 vccd1 vccd1 _11982_/C sky130_fd_sc_hd__and2_1
XFILLER_0_126_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12799_ hold27/X _12798_/B _12798_/Y _13113_/A vssd1 vssd1 vccd1 vccd1 hold28/A sky130_fd_sc_hd__o211a_1
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06664__B _12649_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10467__A _11470_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09569__B1 _10165_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07010_ reg1_val[26] _07010_/B vssd1 vssd1 vccd1 vccd1 _07013_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_122_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_4_14_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13117__B2 _12790_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_86 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08961_ _08962_/B _08962_/A vssd1 vssd1 vccd1 vccd1 _08961_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_11_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08892_ _08893_/A _08893_/B vssd1 vssd1 vccd1 vccd1 _08901_/A sky130_fd_sc_hd__nand2_1
X_07912_ _07912_/A _07912_/B vssd1 vssd1 vccd1 vccd1 _07913_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__10930__A _11171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11143__A3 _10996_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07843_ _07810_/A _07810_/B _07808_/X vssd1 vssd1 vccd1 vccd1 _07846_/A sky130_fd_sc_hd__a21o_1
XANTENNA_fanout189_A _09127_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06839__B _07343_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07774_ _11758_/A _07774_/B vssd1 vssd1 vccd1 vccd1 _07776_/B sky130_fd_sc_hd__xnor2_1
X_06725_ _11021_/S _06725_/B vssd1 vssd1 vccd1 vccd1 _11004_/A sky130_fd_sc_hd__nor2_1
X_09513_ _09345_/A _09345_/B _09344_/A vssd1 vssd1 vccd1 vccd1 _09517_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_78_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06656_ instruction[32] _06694_/B vssd1 vssd1 vccd1 vccd1 _12659_/B sky130_fd_sc_hd__and2_4
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09444_ _09444_/A fanout7/X vssd1 vssd1 vccd1 vccd1 _09445_/B sky130_fd_sc_hd__nor2_1
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06587_ instruction[0] instruction[1] instruction[2] instruction[41] pred_val vssd1
+ vssd1 vccd1 vccd1 _06587_/X sky130_fd_sc_hd__o311a_4
X_09375_ _11142_/S _09373_/X _09374_/Y _09372_/Y vssd1 vssd1 vccd1 vccd1 dest_val[1]
+ sky130_fd_sc_hd__a31o_4
XFILLER_0_47_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10096__B _10096_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08326_ _08322_/A _08322_/B _08325_/Y vssd1 vssd1 vccd1 vccd1 _08349_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_19_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07283__B2 _09440_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07283__A1 _09238_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08257_ _08722_/A _08257_/B vssd1 vssd1 vccd1 vccd1 _08330_/A sky130_fd_sc_hd__xnor2_2
X_07208_ _07208_/A _07208_/B vssd1 vssd1 vccd1 vccd1 _07208_/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_62_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08188_ _08241_/A _08241_/B vssd1 vssd1 vccd1 vccd1 _08242_/A sky130_fd_sc_hd__or2_1
X_07139_ _07139_/A _07139_/B vssd1 vssd1 vccd1 vccd1 _07139_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__13108__B2 _06572_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06794__B1 _06792_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10150_ _10567_/A fanout15/X _07282_/B _10664_/A vssd1 vssd1 vccd1 vccd1 _10151_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_100_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10081_ _09871_/A _09871_/B _09870_/A vssd1 vssd1 vccd1 vccd1 _10086_/A sky130_fd_sc_hd__o21ai_2
XANTENNA__08535__B2 _08798_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08535__A1 _08673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06749__B _07095_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08310__A _08731_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10983_ _10983_/A _10983_/B vssd1 vssd1 vccd1 vccd1 _10985_/B sky130_fd_sc_hd__xnor2_1
X_12722_ reg1_val[19] _12741_/B vssd1 vssd1 vccd1 vccd1 _12725_/D sky130_fd_sc_hd__xnor2_4
XANTENNA__11842__A1 _11758_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12653_ reg1_val[6] _12654_/B vssd1 vssd1 vccd1 vccd1 _12655_/A sky130_fd_sc_hd__nor2_1
XANTENNA__10287__A _11269_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12584_ _12585_/B vssd1 vssd1 vccd1 vccd1 _12584_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_93_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08980__A _12423_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11604_ _11700_/B _11700_/C vssd1 vssd1 vccd1 vccd1 _11785_/A sky130_fd_sc_hd__nor2_1
X_11535_ _12394_/A _11024_/Y _11534_/Y _06924_/X vssd1 vssd1 vccd1 vccd1 _11535_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_80_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13205_ _13210_/A hold255/X vssd1 vssd1 vccd1 vccd1 _13371_/D sky130_fd_sc_hd__and2_1
XFILLER_0_33_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11466_ _11466_/A _11466_/B vssd1 vssd1 vccd1 vccd1 _11469_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_96_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08223__B1 _08617_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11397_ _11397_/A _11397_/B vssd1 vssd1 vccd1 vccd1 _11398_/B sky130_fd_sc_hd__nor2_1
X_10417_ _07048_/A _07048_/B _11294_/A vssd1 vssd1 vccd1 vccd1 _10419_/B sky130_fd_sc_hd__a21o_1
X_13136_ hold288/A _13135_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13136_/X sky130_fd_sc_hd__mux2_1
X_10348_ _10213_/A _10212_/B _10210_/X vssd1 vssd1 vccd1 vccd1 _10353_/A sky130_fd_sc_hd__a21o_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10581__A1 fanout66/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10030__B1 _07282_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13067_ _10422_/A _13087_/B2 hold124/X vssd1 vssd1 vccd1 vccd1 hold125/A sky130_fd_sc_hd__o21a_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10279_ fanout94/X _10571_/B _10570_/B _10941_/A vssd1 vssd1 vccd1 vccd1 _10280_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10581__B2 _07087_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12018_ _12093_/B _12016_/X _11935_/X _11940_/A vssd1 vssd1 vccd1 vccd1 _12019_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_76_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07490_ _07491_/A _07491_/B vssd1 vssd1 vccd1 vccd1 _09209_/B sky130_fd_sc_hd__or2_1
XFILLER_0_48_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13035__B1 _09897_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09160_ _11624_/A _12402_/A0 _08680_/A vssd1 vssd1 vccd1 vccd1 _09160_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_44_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09091_ _09087_/X _09090_/X _09666_/S vssd1 vssd1 vccd1 vccd1 _09091_/X sky130_fd_sc_hd__mux2_1
XANTENNA__08462__B1 _08564_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08111_ _08111_/A _08111_/B vssd1 vssd1 vccd1 vccd1 _08121_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_44_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08042_ _08042_/A _08042_/B _08042_/C vssd1 vssd1 vccd1 vccd1 _08046_/A sky130_fd_sc_hd__or3_2
XANTENNA__10925__A _11261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09993_ _09830_/A _09978_/X _09980_/Y _09169_/Y _09992_/X vssd1 vssd1 vccd1 vccd1
+ _09993_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_12_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08944_ _08944_/A _08944_/B vssd1 vssd1 vccd1 vccd1 _08946_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12313__A2 _12404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08875_ _08858_/A _08856_/Y _08855_/X vssd1 vssd1 vccd1 vccd1 _08876_/B sky130_fd_sc_hd__a21oi_2
X_07826_ fanout69/X _07885_/B _08721_/B1 _08216_/B vssd1 vssd1 vccd1 vccd1 _07827_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09660__S _09666_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07757_ _08752_/A fanout24/X _07819_/B _08798_/B2 vssd1 vssd1 vccd1 vccd1 _07758_/B
+ sky130_fd_sc_hd__o22a_1
X_06708_ reg2_val[15] _06720_/B vssd1 vssd1 vccd1 vccd1 _06708_/X sky130_fd_sc_hd__and2_1
XFILLER_0_79_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07688_ _08752_/A _07688_/B vssd1 vssd1 vccd1 vccd1 _07689_/B sky130_fd_sc_hd__nor2_1
X_06639_ _12195_/S _06639_/B vssd1 vssd1 vccd1 vccd1 _12176_/A sky130_fd_sc_hd__or2_2
X_09427_ _09427_/A _09427_/B vssd1 vssd1 vccd1 vccd1 _09428_/B sky130_fd_sc_hd__or2_1
X_09358_ _09837_/A _09356_/X _09357_/Y _06939_/Y _09663_/S vssd1 vssd1 vccd1 vccd1
+ _09358_/X sky130_fd_sc_hd__o32a_1
XANTENNA__09896__A _10449_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08309_ _08730_/A1 _08741_/B2 _08038_/A _12820_/A vssd1 vssd1 vccd1 vccd1 _08310_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout17_A _12852_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11052__A2 _11989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09289_ _07556_/A _07556_/B _07554_/X vssd1 vssd1 vccd1 vccd1 _09291_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_50_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11320_ _11320_/A _11514_/A vssd1 vssd1 vccd1 vccd1 _11320_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_50_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08305__A _08724_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11251_ _11218_/Y _11219_/X _11221_/Y _11876_/A _11250_/X vssd1 vssd1 vccd1 vccd1
+ _11251_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_101_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11182_ _11183_/A _11183_/B vssd1 vssd1 vccd1 vccd1 _11182_/X sky130_fd_sc_hd__and2_1
X_10202_ _11269_/A _10202_/B vssd1 vssd1 vccd1 vccd1 _10205_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_101_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10133_ _10133_/A _10133_/B vssd1 vssd1 vccd1 vccd1 _10133_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__11666__A _12317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10570__A _10570_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10064_ _11065_/A _11171_/A _10963_/A fanout24/X vssd1 vssd1 vccd1 vccd1 _10065_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07731__A2 fanout87/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10966_ _10966_/A _10966_/B vssd1 vssd1 vccd1 vccd1 _10967_/C sky130_fd_sc_hd__nand2_1
X_10897_ _09527_/B _09354_/B _10897_/S vssd1 vssd1 vccd1 vccd1 _10897_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_85_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07495__A1 _12848_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07495__B2 _10941_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12705_ _12705_/A _12705_/B _12705_/C vssd1 vssd1 vccd1 vccd1 _12706_/B sky130_fd_sc_hd__and3_2
XFILLER_0_127_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12636_ _12636_/A _12636_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[2] sky130_fd_sc_hd__xnor2_4
XFILLER_0_127_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09236__A2 _12854_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11043__A2 _06986_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12567_ _12554_/B _12559_/B _12623_/A vssd1 vssd1 vccd1 vccd1 _12582_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_81_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10745__A _10782_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold208 hold208/A vssd1 vssd1 vccd1 vccd1 hold208/X sky130_fd_sc_hd__dlygate4sd3_1
X_12498_ _12664_/B _12499_/B vssd1 vssd1 vccd1 vccd1 _12509_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_80_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11518_ _11649_/C vssd1 vssd1 vccd1 vccd1 _11518_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_40_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold219 hold219/A vssd1 vssd1 vccd1 vccd1 hold219/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11449_ hold174/A _11449_/B vssd1 vssd1 vccd1 vccd1 _11544_/B sky130_fd_sc_hd__or2_1
XFILLER_0_40_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10003__B1 _07035_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13119_ _12901_/X _13119_/B vssd1 vssd1 vccd1 vccd1 _13120_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__06758__B1 _06757_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06990_ _11163_/A _06990_/B vssd1 vssd1 vccd1 vccd1 _06992_/B sky130_fd_sc_hd__xnor2_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10306__B2 _10413_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10306__A1 _10567_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08660_ _08689_/A _08689_/B _08689_/C vssd1 vssd1 vccd1 vccd1 _08660_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__07722__A2 _10167_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07611_ _12810_/A _10570_/A _10571_/A _10413_/A vssd1 vssd1 vccd1 vccd1 _07612_/B
+ sky130_fd_sc_hd__o22a_1
X_08591_ _08591_/A _08591_/B vssd1 vssd1 vccd1 vccd1 _08594_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_49_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07542_ _10664_/A _11653_/A fanout66/X _07075_/Y vssd1 vssd1 vccd1 vccd1 _07543_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_49_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07473_ _10710_/A _07473_/B vssd1 vssd1 vccd1 vccd1 _07477_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_119_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09212_ _09212_/A _09212_/B _09210_/X vssd1 vssd1 vccd1 vccd1 _09213_/B sky130_fd_sc_hd__or3b_2
XFILLER_0_63_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07013__B _07013_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09143_ _09141_/X _09142_/X _09336_/S vssd1 vssd1 vccd1 vccd1 _09143_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout221_A _06890_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09074_ _09058_/B _09063_/X _09072_/Y _09073_/X _09071_/X vssd1 vssd1 vccd1 vccd1
+ _09075_/B sky130_fd_sc_hd__o311ai_4
XANTENNA__08125__A _08731_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout2 fanout2/A vssd1 vssd1 vccd1 vccd1 fanout2/X sky130_fd_sc_hd__buf_6
X_08025_ _07840_/A _07840_/C _07840_/B vssd1 vssd1 vccd1 vccd1 _08026_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_4_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07410__A1 _12826_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11742__B1 _12213_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09976_ _11118_/A _09976_/B vssd1 vssd1 vccd1 vccd1 _09976_/X sky130_fd_sc_hd__or2_1
XANTENNA__07410__B2 _12828_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06764__A3 _12659_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08927_ _08000_/A _08000_/B _08002_/B _08003_/X vssd1 vssd1 vccd1 vccd1 _08929_/B
+ sky130_fd_sc_hd__a31oi_4
X_08858_ _08858_/A _08858_/B vssd1 vssd1 vccd1 vccd1 _08859_/B sky130_fd_sc_hd__xnor2_2
X_07809_ _07809_/A _07809_/B vssd1 vssd1 vccd1 vccd1 _07810_/B sky130_fd_sc_hd__xnor2_1
X_08789_ _08780_/A _08780_/B _08782_/Y vssd1 vssd1 vccd1 vccd1 _08838_/A sky130_fd_sc_hd__o21ai_4
X_10820_ _10820_/A _10820_/B vssd1 vssd1 vccd1 vccd1 _10821_/B sky130_fd_sc_hd__xnor2_1
X_10751_ _06818_/X _10750_/X _12174_/S vssd1 vssd1 vccd1 vccd1 _10752_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_39_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12421_ _12411_/X _12419_/Y _12420_/Y vssd1 vssd1 vccd1 vccd1 _12421_/X sky130_fd_sc_hd__o21a_1
X_10682_ _10681_/A _10681_/B _10680_/X vssd1 vssd1 vccd1 vccd1 _10695_/B sky130_fd_sc_hd__o21bai_1
XFILLER_0_124_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10565__A _10959_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12352_ hold266/A _12352_/B vssd1 vssd1 vccd1 vccd1 _12396_/B sky130_fd_sc_hd__or2_1
XFILLER_0_105_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10784__A1 _10941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12283_ _12160_/A _12222_/Y _12224_/B vssd1 vssd1 vccd1 vccd1 _12283_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__10784__B2 fanout94/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11303_ _11303_/A _11303_/B _11303_/C vssd1 vssd1 vccd1 vccd1 _11304_/B sky130_fd_sc_hd__or3_1
X_11234_ _11886_/A _11234_/B vssd1 vssd1 vccd1 vccd1 _11234_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_105_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07874__A _08728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11165_ _10941_/A fanout12/X fanout8/X fanout94/X vssd1 vssd1 vccd1 vccd1 _11166_/B
+ sky130_fd_sc_hd__o22a_1
X_10116_ _10114_/X _10115_/X _11010_/S vssd1 vssd1 vccd1 vccd1 _10116_/X sky130_fd_sc_hd__mux2_1
X_11096_ _11097_/A _11097_/B _11097_/C vssd1 vssd1 vccd1 vccd1 _11098_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_117_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10047_ _10047_/A _10047_/B vssd1 vssd1 vccd1 vccd1 _10061_/A sky130_fd_sc_hd__xor2_1
Xhold80 hold80/A vssd1 vssd1 vccd1 vccd1 hold80/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold91 hold91/A vssd1 vssd1 vccd1 vccd1 hold91/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11998_ _12261_/A _11998_/B vssd1 vssd1 vccd1 vccd1 _12002_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_97_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10949_ _10949_/A _10949_/B vssd1 vssd1 vccd1 vccd1 _10950_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_42_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06953__A _10710_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12619_ _12612_/B _12614_/B _12612_/A vssd1 vssd1 vccd1 vccd1 _12620_/B sky130_fd_sc_hd__o21ba_2
XFILLER_0_53_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10775__A1 _12254_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11972__B1 _12247_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07640__A1 _12804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07640__B2 _09613_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09830_ _09830_/A vssd1 vssd1 vccd1 vccd1 _09830_/Y sky130_fd_sc_hd__inv_2
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06973_ _07130_/A _06973_/B vssd1 vssd1 vccd1 vccd1 _12828_/A sky130_fd_sc_hd__xnor2_4
X_09761_ _09761_/A _09761_/B vssd1 vssd1 vccd1 vccd1 _09762_/B sky130_fd_sc_hd__and2_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08712_ _08382_/A _08382_/B _08382_/C vssd1 vssd1 vccd1 vccd1 _08715_/B sky130_fd_sc_hd__o21ai_2
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09692_ hold284/A _09691_/X _09167_/Y vssd1 vssd1 vccd1 vccd1 _09692_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_83_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08643_ _08652_/A _08643_/B _08643_/C vssd1 vssd1 vccd1 vccd1 _08650_/A sky130_fd_sc_hd__nand3_1
XANTENNA_fanout171_A _09440_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout269_A _06770_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08574_ _08574_/A _08574_/B vssd1 vssd1 vccd1 vccd1 _08586_/A sky130_fd_sc_hd__or2_1
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07525_ _07526_/A _07526_/B vssd1 vssd1 vccd1 vccd1 _07527_/A sky130_fd_sc_hd__and2_1
XFILLER_0_49_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10463__B1 _10570_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07959__A _11758_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07456_ _07456_/A _07456_/B _07562_/A vssd1 vssd1 vccd1 vccd1 _07457_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_45_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10385__A _11118_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08408__B1 _08617_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07387_ _07116_/A _07116_/B _07112_/X vssd1 vssd1 vccd1 vccd1 _07389_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_106_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09126_ reg1_val[14] reg1_val[17] _09127_/S vssd1 vssd1 vccd1 vccd1 _09126_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_72_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09057_ _09065_/C _09065_/D _09055_/Y vssd1 vssd1 vccd1 vccd1 _09058_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_60_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09620__A2 _11653_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08008_ _08008_/A _08008_/B vssd1 vssd1 vccd1 vccd1 _08021_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_20_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09959_ _09958_/A _09958_/B _12290_/A vssd1 vssd1 vccd1 vccd1 _09959_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout84_A _12830_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12970_ hold187/X _13004_/A2 _13016_/B1 hold185/X vssd1 vssd1 vccd1 vccd1 hold188/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__06757__B _06799_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07698__A1 _08436_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07698__B2 _07149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11921_ _12067_/A fanout9/X fanout4/X _11989_/A vssd1 vssd1 vccd1 vccd1 _11922_/B
+ sky130_fd_sc_hd__o22a_1
X_11852_ _11853_/A _11853_/B vssd1 vssd1 vccd1 vccd1 _11852_/X sky130_fd_sc_hd__and2b_1
XANTENNA__11246__A2 _12404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12443__A1 _07064_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10803_ _10913_/C _10802_/C _10802_/A vssd1 vssd1 vccd1 vccd1 _10814_/B sky130_fd_sc_hd__a21o_1
XANTENNA__07869__A _08733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11783_ _11783_/A _11783_/B vssd1 vssd1 vccd1 vccd1 _12098_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_67_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10734_ _10612_/A _10610_/X _10609_/X vssd1 vssd1 vccd1 vccd1 _10737_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_27_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10665_ _10665_/A _10665_/B vssd1 vssd1 vccd1 vccd1 _10669_/A sky130_fd_sc_hd__xor2_1
XANTENNA__07870__B2 _08730_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07870__A1 _08038_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13384_ _13384_/CLK hold161/X vssd1 vssd1 vccd1 vccd1 hold160/A sky130_fd_sc_hd__dfxtp_1
X_12404_ _12404_/A _12404_/B vssd1 vssd1 vccd1 vccd1 _12404_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_88_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12335_ _12101_/B _12332_/Y _12333_/Y _12334_/Y vssd1 vssd1 vccd1 vccd1 _12336_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_2_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10596_ _10596_/A _10596_/B vssd1 vssd1 vccd1 vccd1 _10597_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_23_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12266_ _12266_/A _12266_/B vssd1 vssd1 vccd1 vccd1 _12267_/B sky130_fd_sc_hd__nand2_1
XANTENNA__11838__B _11839_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12197_ _07140_/B _11343_/B _12254_/A1 _09968_/A _12196_/X vssd1 vssd1 vccd1 vccd1
+ _12197_/Y sky130_fd_sc_hd__o221ai_1
XANTENNA__09375__A1 _11142_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11217_ _11421_/A _11217_/B vssd1 vssd1 vccd1 vccd1 _11650_/C sky130_fd_sc_hd__xor2_4
XANTENNA__07109__A _07522_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11148_ _11148_/A _11148_/B vssd1 vssd1 vccd1 vccd1 _11150_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_128_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12669__B _12669_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_78 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11079_ _11079_/A _11079_/B vssd1 vssd1 vccd1 vccd1 _11092_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__11890__C1 _12247_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06667__B _07220_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08350__A2 _09567_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07310_ _07602_/A _07602_/B _07272_/Y vssd1 vssd1 vccd1 vccd1 _07401_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_128_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_387 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08290_ _08290_/A _08346_/A vssd1 vssd1 vccd1 vccd1 _08298_/A sky130_fd_sc_hd__and2_1
X_07241_ _07241_/A _07241_/B vssd1 vssd1 vccd1 vccd1 _07302_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_73_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07172_ _07173_/A _07173_/B vssd1 vssd1 vccd1 vccd1 _07172_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_6_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_446 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13162__A2 _06890_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout304 _06577_/Y vssd1 vssd1 vccd1 vccd1 _12388_/S sky130_fd_sc_hd__buf_4
XFILLER_0_78_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09813_ _09704_/X _09853_/C _09812_/Y vssd1 vssd1 vccd1 vccd1 _09813_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__07019__A _11673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06956_ _12341_/A _07064_/B vssd1 vssd1 vccd1 vccd1 _07220_/B sky130_fd_sc_hd__and2_2
X_09744_ _07099_/A _07099_/B _10418_/A vssd1 vssd1 vccd1 vccd1 _09746_/B sky130_fd_sc_hd__a21o_1
XTAP_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06887_ instruction[6] instruction[5] instruction[4] vssd1 vssd1 vccd1 vccd1 _06887_/Y
+ sky130_fd_sc_hd__a21oi_2
X_09675_ reg1_val[3] curr_PC[3] vssd1 vssd1 vccd1 vccd1 _09675_/X sky130_fd_sc_hd__or2_1
XFILLER_0_69_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09234__A _09906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08626_ _08621_/A _08621_/B _08621_/C vssd1 vssd1 vccd1 vccd1 _08626_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__10684__B1 fanout27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13190__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08557_ _08577_/A vssd1 vssd1 vccd1 vccd1 _08557_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_37_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08488_ _08489_/A _08489_/B _08489_/C vssd1 vssd1 vccd1 vccd1 _09018_/A sky130_fd_sc_hd__o21a_1
XANTENNA__07689__A _11673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07508_ _10928_/A _07508_/B _10959_/A vssd1 vssd1 vccd1 vccd1 _07510_/A sky130_fd_sc_hd__or3_2
XANTENNA__10436__B1 _07688_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07439_ _07460_/B _07414_/B _07438_/B _07563_/A _07563_/B vssd1 vssd1 vccd1 vccd1
+ _07459_/A sky130_fd_sc_hd__a32o_2
XANTENNA__12189__B1 _12247_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10450_ _10449_/B _10449_/C _10449_/A vssd1 vssd1 vccd1 vccd1 _10451_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_17_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09109_ _09107_/X _09108_/X _09330_/S vssd1 vssd1 vccd1 vccd1 _09109_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_32_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10381_ reg1_val[8] curr_PC[8] vssd1 vssd1 vccd1 vccd1 _10381_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_20_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12120_ _11636_/B _12187_/B hold261/A vssd1 vssd1 vccd1 vccd1 _12122_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__08313__A _08728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09357__A1 hold260/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12051_ _07166_/A _12404_/A _09152_/Y _10246_/X _12050_/X vssd1 vssd1 vccd1 vccd1
+ _12051_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11002_ _06820_/X _11001_/X _12174_/S vssd1 vssd1 vccd1 vccd1 _11004_/B sky130_fd_sc_hd__mux2_1
XANTENNA__07368__B1 _07282_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12953_ _12863_/X _12953_/B vssd1 vssd1 vccd1 vccd1 _13220_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_99_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11467__A2 _12213_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11904_ _11872_/B _11872_/C _11874_/A vssd1 vssd1 vccd1 vccd1 _11951_/B sky130_fd_sc_hd__o21a_1
X_12884_ hold271/X hold17/X vssd1 vssd1 vccd1 vccd1 _13164_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_99_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11219__A2 _11650_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11835_ _12073_/A _11835_/B vssd1 vssd1 vccd1 vccd1 _11839_/A sky130_fd_sc_hd__xnor2_1
XTAP_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11766_ _11766_/A _12214_/B vssd1 vssd1 vccd1 vccd1 _11766_/X sky130_fd_sc_hd__or2_1
XFILLER_0_23_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10717_ _10717_/A _10717_/B vssd1 vssd1 vccd1 vccd1 _10731_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_126_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11697_ _11697_/A _11697_/B _11697_/C vssd1 vssd1 vccd1 vccd1 _11698_/B sky130_fd_sc_hd__nand3_1
X_10648_ hold269/A _09835_/B _10769_/B _10647_/Y _09837_/A vssd1 vssd1 vccd1 vccd1
+ _10648_/X sky130_fd_sc_hd__a311o_2
XFILLER_0_63_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13367_ _13376_/CLK _13367_/D vssd1 vssd1 vccd1 vccd1 hold275/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10579_ _10579_/A _10579_/B _10579_/C _10579_/D vssd1 vssd1 vccd1 vccd1 _10580_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_0_23_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13298_ _13299_/CLK _13298_/D vssd1 vssd1 vccd1 vccd1 hold183/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12318_ _12319_/A _12319_/B vssd1 vssd1 vccd1 vccd1 _12320_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_121_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12249_ _12434_/B1 _12304_/B hold195/A vssd1 vssd1 vccd1 vccd1 _12249_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_48_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10902__B2 _09111_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06810_ _09527_/A _06809_/X _06795_/X vssd1 vssd1 vccd1 vccd1 _06810_/X sky130_fd_sc_hd__a21o_1
XANTENNA__12104__B1 _12290_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07790_ _07790_/A _07790_/B vssd1 vssd1 vccd1 vccd1 _07881_/A sky130_fd_sc_hd__xnor2_2
X_06741_ reg1_val[10] _07100_/A vssd1 vssd1 vccd1 vccd1 _10644_/S sky130_fd_sc_hd__and2_1
XFILLER_0_78_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09460_ _09460_/A _09460_/B vssd1 vssd1 vccd1 vccd1 _09462_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__08323__A2 _08744_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10666__B1 fanout4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06672_ reg2_val[21] _06720_/B _06703_/B1 _06671_/Y vssd1 vssd1 vccd1 vccd1 _07135_/D
+ sky130_fd_sc_hd__o2bb2a_4
X_08411_ _08745_/A _08411_/B vssd1 vssd1 vccd1 vccd1 _08443_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07531__B1 _10963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09391_ _09391_/A _09391_/B vssd1 vssd1 vccd1 vccd1 _09393_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__06885__A2 _06921_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10928__A _10928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08342_ _08342_/A _08342_/B _08343_/B vssd1 vssd1 vccd1 vccd1 _08342_/X sky130_fd_sc_hd__and3_1
XFILLER_0_19_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08273_ _08721_/B1 _08741_/A2 _08617_/B _08739_/A1 vssd1 vssd1 vccd1 vccd1 _08274_/B
+ sky130_fd_sc_hd__o22a_1
X_07224_ _07220_/A _07220_/C _07074_/B _07135_/D vssd1 vssd1 vccd1 vccd1 _07226_/A
+ sky130_fd_sc_hd__o211ai_1
XFILLER_0_73_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout301_A _13242_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07155_ _07149_/A _12852_/A _08632_/C _12264_/A vssd1 vssd1 vccd1 vccd1 _07156_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_42_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10663__A _10928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09229__A _11385_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07086_ _11269_/A _07090_/B _11261_/A vssd1 vssd1 vccd1 vccd1 _07087_/B sky130_fd_sc_hd__a21oi_4
XANTENNA__08133__A _11385_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout101 _07485_/A vssd1 vssd1 vccd1 vccd1 _11385_/A sky130_fd_sc_hd__clkbuf_16
Xfanout112 _07522_/A vssd1 vssd1 vccd1 vccd1 _12076_/A sky130_fd_sc_hd__clkbuf_16
XANTENNA__13185__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout134 _07165_/X vssd1 vssd1 vccd1 vccd1 _09238_/B sky130_fd_sc_hd__buf_8
Xfanout145 _09768_/A1 vssd1 vssd1 vccd1 vccd1 _08723_/B1 sky130_fd_sc_hd__buf_6
Xfanout156 _10748_/A vssd1 vssd1 vccd1 vccd1 _12031_/A sky130_fd_sc_hd__clkbuf_4
Xfanout123 _10927_/A1 vssd1 vssd1 vccd1 vccd1 _11294_/A sky130_fd_sc_hd__buf_6
Xfanout189 _09127_/S vssd1 vssd1 vccd1 vccd1 _09142_/S sky130_fd_sc_hd__clkbuf_8
Xfanout167 _08584_/A vssd1 vssd1 vccd1 vccd1 _10449_/A sky130_fd_sc_hd__clkbuf_16
Xfanout178 _07128_/X vssd1 vssd1 vccd1 vccd1 _09444_/A sky130_fd_sc_hd__buf_4
XANTENNA__08562__A2 _09567_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07988_ _07989_/A _07989_/B vssd1 vssd1 vccd1 vccd1 _08925_/B sky130_fd_sc_hd__nand2b_1
X_06939_ _12423_/A _06939_/B vssd1 vssd1 vccd1 vccd1 _06939_/Y sky130_fd_sc_hd__nand2_4
X_09727_ _09619_/B _09622_/B _09617_/X vssd1 vssd1 vccd1 vccd1 _09730_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_97_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09658_ _12428_/A _09658_/B _09658_/C vssd1 vssd1 vccd1 vccd1 _09699_/B sky130_fd_sc_hd__and3_1
XFILLER_0_69_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout47_A _12838_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08609_ _08609_/A _08609_/B vssd1 vssd1 vccd1 vccd1 _08697_/B sky130_fd_sc_hd__xor2_1
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09589_ _09732_/B _09589_/B vssd1 vssd1 vccd1 vccd1 _09596_/A sky130_fd_sc_hd__or2_1
XANTENNA__13214__A _13214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11620_ _06866_/B _11526_/B _11540_/A vssd1 vssd1 vccd1 vccd1 _11621_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__13071__A1 _11987_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09275__B1 _08752_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07212__A _10710_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11551_ curr_PC[18] _11550_/B _11142_/S vssd1 vssd1 vccd1 vccd1 _11551_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__08308__A _08733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07825__A1 _12073_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10502_ _11792_/A _10410_/Y _10500_/Y _10501_/Y _11707_/A vssd1 vssd1 vccd1 vccd1
+ _10502_/X sky130_fd_sc_hd__o311a_1
XFILLER_0_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11482_ _11751_/A fanout9/X fanout4/X _11558_/A vssd1 vssd1 vccd1 vccd1 _11483_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_18_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11909__B1 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13221_ hold256/X _13220_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13221_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_100_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10433_ _10440_/A vssd1 vssd1 vccd1 vccd1 _10433_/Y sky130_fd_sc_hd__inv_2
XANTENNA__10188__A2 _10571_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13152_ hold282/X _06890_/Y _13151_/X _13246_/B2 vssd1 vssd1 vccd1 vccd1 hold283/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__07053__A2 fanout23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10364_ _10364_/A _10364_/B vssd1 vssd1 vccd1 vccd1 _10741_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_103_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12103_ _12103_/A _12103_/B vssd1 vssd1 vccd1 vccd1 _12103_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_103_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13083_ _09548_/A _12798_/B hold74/X vssd1 vssd1 vccd1 vccd1 hold75/A sky130_fd_sc_hd__a21oi_1
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10295_ _10445_/A fanout59/X _10941_/B _10706_/B2 vssd1 vssd1 vccd1 vccd1 _10296_/B
+ sky130_fd_sc_hd__o22a_1
X_12034_ _06836_/B _12033_/Y _12388_/S vssd1 vssd1 vccd1 vccd1 _12034_/X sky130_fd_sc_hd__mux2_1
XANTENNA__07761__B1 _12820_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12936_ _13174_/A _13175_/A _13174_/B vssd1 vssd1 vccd1 vccd1 _13180_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_88_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12867_ hold261/X hold29/X vssd1 vssd1 vccd1 vccd1 _12868_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__06945__B _06994_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11818_ curr_PC[21] _11819_/B vssd1 vssd1 vccd1 vccd1 _11820_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_8_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12798_ _12798_/A _12798_/B vssd1 vssd1 vccd1 vccd1 _12798_/Y sky130_fd_sc_hd__nand2_1
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07122__A _09343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12963__A _13214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11749_ _12317_/A _11749_/B vssd1 vssd1 vccd1 vccd1 _11750_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_119_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12174__S _12174_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06680__B _07210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13117__A2 _12789_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08960_ _08960_/A _08960_/B vssd1 vssd1 vccd1 vccd1 _08962_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_59_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07911_ _07911_/A _07911_/B _07911_/C vssd1 vssd1 vccd1 vccd1 _07913_/B sky130_fd_sc_hd__nand3_1
X_08891_ _08891_/A _08891_/B vssd1 vssd1 vccd1 vccd1 _08893_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__10930__B _10930_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07792__A _08742_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11143__A4 _11650_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07842_ _07836_/A _07836_/B _07837_/X vssd1 vssd1 vccd1 vccd1 _07847_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_75_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09512_ _09532_/B vssd1 vssd1 vccd1 vccd1 _09512_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_78_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07773_ _07955_/A _11653_/A _08752_/B _07896_/A vssd1 vssd1 vccd1 vccd1 _07774_/B
+ sky130_fd_sc_hd__o22a_1
X_06724_ reg1_val[13] _11020_/A vssd1 vssd1 vccd1 vccd1 _06725_/B sky130_fd_sc_hd__nor2_1
XANTENNA__10639__B1 _12244_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06655_ _11973_/A _06655_/B vssd1 vssd1 vccd1 vccd1 _11959_/A sky130_fd_sc_hd__nor2_1
X_09443_ _09593_/A _09443_/B vssd1 vssd1 vccd1 vccd1 _09446_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_66_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13053__A1 _06986_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09374_ curr_PC[0] curr_PC[1] vssd1 vssd1 vccd1 vccd1 _09374_/Y sky130_fd_sc_hd__nand2_1
X_06586_ instruction[0] instruction[1] instruction[2] pred_val vssd1 vssd1 vccd1 vccd1
+ _06586_/X sky130_fd_sc_hd__o31a_1
XFILLER_0_86_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07032__A _10422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08325_ _08373_/B _08373_/A vssd1 vssd1 vccd1 vccd1 _08325_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__08128__A _08728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07283__A2 fanout48/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08256_ _10537_/A1 _07821_/A _07752_/B _08432_/B vssd1 vssd1 vccd1 vccd1 _08257_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10811__B1 _10575_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07207_ _07131_/B _07205_/X _07206_/X _07220_/B vssd1 vssd1 vccd1 vccd1 _07207_/X
+ sky130_fd_sc_hd__a22o_1
X_08187_ _08187_/A _08187_/B vssd1 vssd1 vccd1 vccd1 _08241_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_104_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07138_ _07140_/B _07138_/B vssd1 vssd1 vccd1 vccd1 _07138_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_70_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13108__A2 _06892_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07069_ reg1_val[16] _07069_/B vssd1 vssd1 vccd1 vccd1 _07071_/D sky130_fd_sc_hd__xnor2_1
X_10080_ _09932_/A _09932_/B _09930_/X vssd1 vssd1 vccd1 vccd1 _10090_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_100_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08535__A2 _08744_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10982_ _10983_/A _10983_/B vssd1 vssd1 vccd1 vccd1 _11097_/A sky130_fd_sc_hd__and2_1
X_12721_ _12718_/A _12720_/B _12718_/B vssd1 vssd1 vccd1 vccd1 _12723_/A sky130_fd_sc_hd__a21bo_1
X_12652_ _12651_/A _12648_/Y _12650_/B vssd1 vssd1 vccd1 vccd1 _12656_/A sky130_fd_sc_hd__o21a_2
XFILLER_0_37_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11603_ _11603_/A _11603_/B _11603_/C vssd1 vssd1 vccd1 vccd1 _11700_/C sky130_fd_sc_hd__nor3_1
XANTENNA__08038__A _08038_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12583_ _12605_/A _12607_/A vssd1 vssd1 vccd1 vccd1 _12585_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_93_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12252__C1 _12455_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11534_ _11532_/Y _11533_/X _11886_/A vssd1 vssd1 vccd1 vccd1 _11534_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_53_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11465_ _11465_/A _11465_/B vssd1 vssd1 vccd1 vccd1 _11466_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_18_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13204_ hold254/X _13213_/A2 _13203_/X _13213_/B2 vssd1 vssd1 vccd1 vccd1 hold255/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08223__A1 _08739_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10416_ _10416_/A _10416_/B vssd1 vssd1 vccd1 vccd1 _10430_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_33_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08223__B2 _08436_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11396_ _11396_/A _11396_/B vssd1 vssd1 vccd1 vccd1 _11397_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_0_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10030__A1 _10413_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13135_ _13135_/A _13135_/B vssd1 vssd1 vccd1 vccd1 _13135_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_103_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12307__B1 _12307_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10347_ _10197_/B _10214_/B _10197_/A vssd1 vssd1 vccd1 vccd1 _10358_/A sky130_fd_sc_hd__o21ba_1
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10030__B2 _10567_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13066_ hold130/A _12791_/A _13080_/B1 hold123/X _13113_/A vssd1 vssd1 vccd1 vccd1
+ hold124/A sky130_fd_sc_hd__o221a_1
X_10278_ _10225_/A _10225_/B _10223_/Y vssd1 vssd1 vccd1 vccd1 _10361_/A sky130_fd_sc_hd__a21o_2
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10581__A2 fanout48/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11338__S _12244_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10242__S _12388_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10869__B1 _11100_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12017_ _11935_/X _11940_/A _12093_/B _12016_/X vssd1 vssd1 vccd1 vccd1 _12017_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_45_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06956__A _12341_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12919_ _13096_/B _13097_/A _12913_/X vssd1 vssd1 vccd1 vccd1 _13102_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_88_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13035__B2 _13087_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09239__B1 _09440_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09090_ _09088_/X _09089_/X _09336_/S vssd1 vssd1 vccd1 vccd1 _09090_/X sky130_fd_sc_hd__mux2_1
XANTENNA__08462__A1 _08646_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08462__B2 _09423_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08110_ _08110_/A _08110_/B vssd1 vssd1 vccd1 vccd1 _08111_/B sky130_fd_sc_hd__or2_1
XFILLER_0_16_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08041_ _08731_/A _08041_/B _08041_/C vssd1 vssd1 vccd1 vccd1 _08042_/C sky130_fd_sc_hd__and3_1
XFILLER_0_101_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09992_ _12429_/B _09172_/B _09991_/Y _09986_/Y vssd1 vssd1 vccd1 vccd1 _09992_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_3_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10941__A _10941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08943_ _08920_/A _08920_/B _08923_/A vssd1 vssd1 vccd1 vccd1 _08948_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_86_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08411__A _08745_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07725__B1 _11558_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08874_ _08874_/A _08874_/B vssd1 vssd1 vccd1 vccd1 _08876_/A sky130_fd_sc_hd__xnor2_2
X_07825_ _12073_/A _07824_/A _07824_/X vssd1 vssd1 vccd1 vccd1 _07838_/A sky130_fd_sc_hd__o21bai_1
X_07756_ _07856_/A _07856_/B _07753_/Y _07754_/X vssd1 vssd1 vccd1 vccd1 _07759_/B
+ sky130_fd_sc_hd__o211ai_2
X_06707_ _06705_/X _06707_/B vssd1 vssd1 vccd1 vccd1 _11332_/A sky130_fd_sc_hd__and2b_1
XANTENNA__09242__A _09593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06585__B _06771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09426_ _09427_/A _09427_/B vssd1 vssd1 vccd1 vccd1 _09426_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_66_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07687_ _11908_/A _07687_/B vssd1 vssd1 vccd1 vccd1 _07691_/A sky130_fd_sc_hd__xnor2_1
X_06638_ reg1_val[26] _07140_/B vssd1 vssd1 vccd1 vccd1 _06639_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_66_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06569_ hold79/X vssd1 vssd1 vccd1 vccd1 hold80/A sky130_fd_sc_hd__inv_2
X_09357_ hold260/A _09835_/B hold244/A vssd1 vssd1 vccd1 vccd1 _09357_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_47_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11037__B1 _10930_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11711__S _12174_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09288_ _07519_/A _07519_/B _07516_/Y vssd1 vssd1 vccd1 vccd1 _09291_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_74_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08308_ _08733_/A _08308_/B vssd1 vssd1 vccd1 vccd1 _08315_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_35_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08239_ _08282_/A _08237_/Y _08227_/Y vssd1 vssd1 vccd1 vccd1 _08249_/B sky130_fd_sc_hd__o21a_1
XANTENNA__11012__A _12394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11250_ _11250_/A _11250_/B _11250_/C vssd1 vssd1 vccd1 vccd1 _11250_/X sky130_fd_sc_hd__or3_2
XANTENNA__09402__B1 _11987_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11181_ _11181_/A _11181_/B vssd1 vssd1 vccd1 vccd1 _11183_/B sky130_fd_sc_hd__xnor2_1
X_10201_ _10570_/A _10575_/B _10930_/B _10571_/A vssd1 vssd1 vccd1 vccd1 _10202_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_101_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10132_ _10130_/Y _10132_/B vssd1 vssd1 vccd1 vccd1 _10133_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_30_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08321__A _08740_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10492__A_N _10493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10570__B _10570_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10063_ _09782_/A _09782_/B _09912_/B _09913_/B _09913_/A vssd1 vssd1 vccd1 vccd1
+ _10078_/A sky130_fd_sc_hd__a32oi_4
XANTENNA__09152__A _12423_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11276__B1 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12704_ _12705_/A _12705_/B _12705_/C vssd1 vssd1 vccd1 vccd1 _12706_/A sky130_fd_sc_hd__a21oi_4
XANTENNA__10298__A _11163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10965_ _10966_/A _10966_/B vssd1 vssd1 vccd1 vccd1 _10967_/B sky130_fd_sc_hd__or2_1
XANTENNA__08141__B1 _08038_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10896_ _10896_/A _10896_/B vssd1 vssd1 vccd1 vccd1 _10896_/Y sky130_fd_sc_hd__nor2_2
XANTENNA__07495__A2 _09238_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11028__B1 _11027_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12635_ _12633_/Y _12635_/B vssd1 vssd1 vccd1 vccd1 _12636_/B sky130_fd_sc_hd__and2b_2
XFILLER_0_26_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12566_ _12566_/A _12566_/B vssd1 vssd1 vccd1 vccd1 _12581_/B sky130_fd_sc_hd__or2_1
XFILLER_0_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11043__A3 _12412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11517_ _11700_/A _11517_/B vssd1 vssd1 vccd1 vccd1 _11649_/C sky130_fd_sc_hd__xor2_4
X_12497_ reg1_val[8] curr_PC[8] _12622_/S vssd1 vssd1 vccd1 vccd1 _12499_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_34_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold209 hold209/A vssd1 vssd1 vccd1 vccd1 hold209/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11448_ _09152_/Y _11443_/B _11447_/X vssd1 vssd1 vccd1 vccd1 _11448_/Y sky130_fd_sc_hd__a21oi_1
X_11379_ fanout24/X _11989_/A _12067_/A _07819_/B vssd1 vssd1 vccd1 vccd1 _11380_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_0_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13118_ _13128_/A hold243/X vssd1 vssd1 vccd1 vccd1 _13353_/D sky130_fd_sc_hd__and2_1
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08231__A _08724_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13049_ _06954_/B _12798_/B hold165/X vssd1 vssd1 vccd1 vccd1 _13327_/D sky130_fd_sc_hd__a21boi_1
XFILLER_0_56_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07707__B1 _10567_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10306__A2 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08590_ _09004_/A _08590_/B vssd1 vssd1 vccd1 vccd1 _09002_/A sky130_fd_sc_hd__and2_1
X_07610_ _07610_/A _07610_/B vssd1 vssd1 vccd1 vccd1 _07992_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_72_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07541_ _09212_/A _07541_/B vssd1 vssd1 vccd1 vccd1 _07545_/A sky130_fd_sc_hd__nand2b_2
XFILLER_0_88_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08132__B1 _08216_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07472_ _12838_/A _08507_/B _12836_/A _10589_/A vssd1 vssd1 vccd1 vccd1 _07473_/B
+ sky130_fd_sc_hd__o22a_1
X_09211_ _09212_/A _09212_/B _09210_/X vssd1 vssd1 vccd1 vccd1 _09211_/X sky130_fd_sc_hd__o21ba_1
X_09142_ reg1_val[7] reg1_val[24] _09142_/S vssd1 vssd1 vccd1 vccd1 _09142_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_56_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09073_ _09073_/A _09073_/B _09073_/C _09072_/B vssd1 vssd1 vccd1 vccd1 _09073_/X
+ sky130_fd_sc_hd__or4b_2
XFILLER_0_44_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08024_ _08024_/A _08024_/B vssd1 vssd1 vccd1 vccd1 _08909_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_102_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09237__A _09594_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11742__B2 fanout27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11742__A1 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07946__B1 _08216_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09975_ _10250_/S _09328_/X _09974_/X vssd1 vssd1 vccd1 vccd1 _09975_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__07410__A2 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08926_ _07991_/A _07991_/B _07997_/B _07996_/B _07996_/A vssd1 vssd1 vccd1 vccd1
+ _08929_/A sky130_fd_sc_hd__o32a_2
X_08857_ _08857_/A _08857_/B vssd1 vssd1 vccd1 vccd1 _08858_/B sky130_fd_sc_hd__xor2_1
X_07808_ _07808_/A _07808_/B _07809_/B vssd1 vssd1 vccd1 vccd1 _07808_/X sky130_fd_sc_hd__and3_1
X_08788_ _08788_/A _08788_/B vssd1 vssd1 vccd1 vccd1 _09036_/B sky130_fd_sc_hd__nor2_1
XANTENNA__11258__B1 _12067_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07739_ _07813_/A _07813_/B vssd1 vssd1 vccd1 vccd1 _07741_/C sky130_fd_sc_hd__or2_1
X_10750_ _10629_/A _10627_/Y _10644_/S vssd1 vssd1 vccd1 vccd1 _10750_/X sky130_fd_sc_hd__a21o_1
X_09409_ _09251_/A _12264_/B _09257_/B _09255_/X vssd1 vssd1 vccd1 vccd1 _09411_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_54_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10681_ _10681_/A _10681_/B _10680_/X vssd1 vssd1 vccd1 vccd1 _10844_/A sky130_fd_sc_hd__nor3b_1
XFILLER_0_109_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12420_ _12411_/X _12419_/Y _12290_/A vssd1 vssd1 vccd1 vccd1 _12420_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_118_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07220__A _07220_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12351_ _12394_/A _09497_/Y _12350_/X _06924_/X vssd1 vssd1 vccd1 vccd1 _12362_/C
+ sky130_fd_sc_hd__a211oi_1
X_12282_ _12380_/C vssd1 vssd1 vccd1 vccd1 _12282_/Y sky130_fd_sc_hd__inv_2
XANTENNA__10784__A2 fanout59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11302_ _11303_/A _11303_/B _11303_/C vssd1 vssd1 vccd1 vccd1 _11304_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_16_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11233_ _09182_/A _11232_/Y _11233_/S vssd1 vssd1 vccd1 vccd1 _11234_/B sky130_fd_sc_hd__mux2_2
XANTENNA__11733__B2 _09163_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11164_ _11164_/A _11164_/B vssd1 vssd1 vccd1 vccd1 _11168_/A sky130_fd_sc_hd__xnor2_1
X_10115_ _09501_/X _09506_/X _10250_/S vssd1 vssd1 vccd1 vccd1 _10115_/X sky130_fd_sc_hd__mux2_1
X_11095_ _11095_/A _11095_/B vssd1 vssd1 vccd1 vccd1 _11097_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_117_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10046_ _10046_/A _10046_/B vssd1 vssd1 vccd1 vccd1 _10047_/B sky130_fd_sc_hd__xnor2_2
Xhold81 hold81/A vssd1 vssd1 vccd1 vccd1 hold81/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold70 hold70/A vssd1 vssd1 vccd1 vccd1 hold70/X sky130_fd_sc_hd__buf_1
XANTENNA__07165__A1 _09441_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold92 hold92/A vssd1 vssd1 vccd1 vccd1 hold92/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13238__B2 _06572_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08114__B1 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11997_ _12150_/A fanout9/X fanout4/X _12067_/A vssd1 vssd1 vccd1 vccd1 _11998_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_85_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10948_ fanout74/X fanout13/X fanout6/X _10948_/B2 vssd1 vssd1 vccd1 vccd1 _10949_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_128_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09610__A _10418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10879_ _10879_/A _10879_/B vssd1 vssd1 vccd1 vccd1 _10879_/X sky130_fd_sc_hd__or2_1
XANTENNA__06953__B _06954_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12618_ _12618_/A _12618_/B vssd1 vssd1 vccd1 vccd1 _12620_/A sky130_fd_sc_hd__nor2_2
XANTENNA__07130__A _07130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12549_ _12556_/A _12549_/B vssd1 vssd1 vccd1 vccd1 _12551_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_81_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07640__A2 _09614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_1 _07178_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07928__B1 _09614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06972_ _11343_/A _06961_/Y _06966_/Y _07223_/B vssd1 vssd1 vccd1 vccd1 _06973_/B
+ sky130_fd_sc_hd__a31o_1
X_09760_ _09761_/A _09761_/B vssd1 vssd1 vccd1 vccd1 _09889_/A sky130_fd_sc_hd__nor2_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09691_ hold240/A hold244/A hold260/A _09835_/B vssd1 vssd1 vccd1 vccd1 _09691_/X
+ sky130_fd_sc_hd__o31a_1
X_08711_ _08711_/A _08711_/B vssd1 vssd1 vccd1 vccd1 _09023_/B sky130_fd_sc_hd__nand2_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06636__A2_N _06771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08642_ _09897_/A _08642_/B vssd1 vssd1 vccd1 vccd1 _08643_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__12437__C1 _12404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08573_ _08573_/A _08573_/B vssd1 vssd1 vccd1 vccd1 _08574_/B sky130_fd_sc_hd__and2_1
XFILLER_0_49_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07524_ _07524_/A _07524_/B vssd1 vssd1 vccd1 vccd1 _07526_/B sky130_fd_sc_hd__xnor2_1
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07455_ _07456_/B _07562_/A _07456_/A vssd1 vssd1 vccd1 vccd1 _09287_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_49_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10463__B2 _10571_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10463__A1 _10570_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08408__B2 _08723_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08408__A1 _12804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07386_ _07453_/A _07386_/B vssd1 vssd1 vccd1 vccd1 _07389_/A sky130_fd_sc_hd__nor2_1
X_09125_ _09123_/X _09124_/X _09330_/S vssd1 vssd1 vccd1 vccd1 _09125_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_60_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09666__S _09666_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09056_ _09056_/A _09056_/B vssd1 vssd1 vccd1 vccd1 _09065_/D sky130_fd_sc_hd__nand2_1
XFILLER_0_44_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08007_ _08007_/A _08007_/B vssd1 vssd1 vccd1 vccd1 _08008_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_102_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09958_ _09958_/A _09958_/B vssd1 vssd1 vccd1 vccd1 _09958_/X sky130_fd_sc_hd__or2_1
X_08909_ _08909_/A _08909_/B vssd1 vssd1 vccd1 vccd1 _08910_/B sky130_fd_sc_hd__nand2_1
XANTENNA_fanout77_A _09548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11436__S _12174_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09889_ _09889_/A _09889_/B vssd1 vssd1 vccd1 vccd1 _09891_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__12140__B2 _12076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07698__A2 _11989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11920_ _11833_/A _11918_/A _11832_/B _11840_/A _11840_/B vssd1 vssd1 vccd1 vccd1
+ _11934_/A sky130_fd_sc_hd__o32a_1
XFILLER_0_79_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11851_ _11853_/B _11853_/A vssd1 vssd1 vccd1 vccd1 _11851_/Y sky130_fd_sc_hd__nand2b_1
X_10802_ _10802_/A _10913_/C _10802_/C vssd1 vssd1 vccd1 vccd1 _10971_/A sky130_fd_sc_hd__and3_1
X_11782_ _11782_/A _11782_/B _11782_/C vssd1 vssd1 vccd1 vccd1 _11783_/B sky130_fd_sc_hd__and3_1
XANTENNA__12443__A2 _06939_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10733_ _10733_/A _10733_/B vssd1 vssd1 vccd1 vccd1 _10737_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_94_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10576__A _11180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11651__B1 fanout12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10664_ _10664_/A _12316_/B vssd1 vssd1 vccd1 vccd1 _10665_/B sky130_fd_sc_hd__or2_1
XANTENNA__07870__A2 _11847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13383_ _13383_/CLK hold54/X vssd1 vssd1 vccd1 vccd1 hold53/A sky130_fd_sc_hd__dfxtp_1
X_12403_ _12403_/A1 _12402_/X _06613_/B vssd1 vssd1 vccd1 vccd1 _12404_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_63_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10595_ _10596_/A _10596_/B vssd1 vssd1 vccd1 vccd1 _10595_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_23_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12334_ _12334_/A _12334_/B vssd1 vssd1 vccd1 vccd1 _12334_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__07885__A _08216_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13098__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12265_ _12266_/A _12266_/B vssd1 vssd1 vccd1 vccd1 _12325_/B sky130_fd_sc_hd__or2_1
XFILLER_0_31_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12196_ _12403_/A1 _12195_/X _06639_/B vssd1 vssd1 vccd1 vccd1 _12196_/X sky130_fd_sc_hd__a21o_1
X_11216_ _10744_/B _11215_/X _11214_/X vssd1 vssd1 vccd1 vccd1 _11217_/B sky130_fd_sc_hd__o21ba_1
XFILLER_0_128_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11147_ _11148_/A _11148_/B vssd1 vssd1 vccd1 vccd1 _11303_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12131__A1 _06924_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11078_ _11078_/A _11078_/B vssd1 vssd1 vccd1 vccd1 _11079_/B sky130_fd_sc_hd__xor2_1
X_10029_ _10029_/A _10029_/B vssd1 vssd1 vccd1 vccd1 _10046_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_58_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12685__B _12686_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07240_ _09445_/A _07240_/B vssd1 vssd1 vccd1 vccd1 _07302_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_116_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12198__A1 _09111_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07171_ _09441_/A _07171_/B vssd1 vssd1 vccd1 vccd1 _07173_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_54_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout305 _07149_/A vssd1 vssd1 vccd1 vccd1 _08730_/A1 sky130_fd_sc_hd__buf_6
XFILLER_0_1_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09812_ _09704_/X _09853_/C _09081_/X vssd1 vssd1 vccd1 vccd1 _09812_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_10_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09743_ _09743_/A _09743_/B vssd1 vssd1 vccd1 vccd1 _09765_/A sky130_fd_sc_hd__xor2_2
X_06955_ _06971_/B _06971_/A _10707_/A vssd1 vssd1 vccd1 vccd1 _06955_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout281_A _07200_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09674_ reg1_val[3] curr_PC[3] vssd1 vssd1 vccd1 vccd1 _09674_/Y sky130_fd_sc_hd__nor2_1
X_06886_ instruction[5] instruction[6] vssd1 vssd1 vccd1 vccd1 _09170_/A sky130_fd_sc_hd__nand2b_4
XTAP_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06888__B1 _09170_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07035__A _07036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08625_ _08625_/A _08625_/B vssd1 vssd1 vccd1 vccd1 _08995_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__10684__B2 _10418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10684__A1 _11294_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08556_ _08728_/A _08556_/B vssd1 vssd1 vccd1 vccd1 _08577_/A sky130_fd_sc_hd__xnor2_2
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07507_ _07417_/Y _07427_/B _07425_/Y vssd1 vssd1 vccd1 vccd1 _07514_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_76_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10436__A1 _11065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08487_ _08487_/A _08487_/B vssd1 vssd1 vccd1 vccd1 _08489_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_49_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10436__B2 _11146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07438_ _07438_/A _07438_/B vssd1 vssd1 vccd1 vccd1 _07563_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_9_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07369_ _09548_/A _07369_/B vssd1 vssd1 vccd1 vccd1 _07371_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_45_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09108_ reg1_val[10] reg1_val[21] _09108_/S vssd1 vssd1 vccd1 vccd1 _09108_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_32_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10380_ _10267_/A _10264_/Y _10266_/B vssd1 vssd1 vccd1 vccd1 _10384_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_32_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09039_ _11793_/A _11792_/B vssd1 vssd1 vccd1 vccd1 _11874_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_4_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11020__A _11020_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12050_ reg1_val[24] _07166_/A _09154_/Y _12049_/X vssd1 vssd1 vccd1 vccd1 _12050_/X
+ sky130_fd_sc_hd__o22a_1
X_11001_ _10879_/A _10876_/X _10897_/S vssd1 vssd1 vccd1 vccd1 _11001_/X sky130_fd_sc_hd__a21o_1
XANTENNA__07368__A1 _08671_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07368__B2 _12798_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06768__B _07036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12952_ hold256/X hold140/X vssd1 vssd1 vccd1 vccd1 _12953_/B sky130_fd_sc_hd__nand2b_1
X_11903_ _11142_/S _11900_/X _11902_/Y vssd1 vssd1 vccd1 vccd1 dest_val[22] sky130_fd_sc_hd__o21ai_4
X_12883_ hold17/X hold271/X vssd1 vssd1 vccd1 vccd1 _12883_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_87_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11834_ fanout24/X _12316_/A fanout12/X _07819_/B vssd1 vssd1 vccd1 vccd1 _11835_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11765_ _11677_/A _11677_/B _11664_/A vssd1 vssd1 vccd1 vccd1 _11775_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_126_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10716_ _10716_/A _10716_/B vssd1 vssd1 vccd1 vccd1 _10717_/B sky130_fd_sc_hd__xnor2_2
X_11696_ _11698_/A vssd1 vssd1 vccd1 vccd1 _11696_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_126_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10647_ _09835_/B _10769_/B hold269/A vssd1 vssd1 vccd1 vccd1 _10647_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_125_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13366_ _13376_/CLK _13366_/D vssd1 vssd1 vccd1 vccd1 hold293/A sky130_fd_sc_hd__dfxtp_2
XFILLER_0_51_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10578_ _10579_/A _10579_/B _10579_/C _10579_/D vssd1 vssd1 vccd1 vccd1 _10578_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_11_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13297_ _13299_/CLK _13297_/D vssd1 vssd1 vccd1 vccd1 hold228/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10658__D_N _10624_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12317_ _12317_/A _12317_/B vssd1 vssd1 vccd1 vccd1 _12319_/B sky130_fd_sc_hd__xnor2_1
X_12248_ hold223/A _12248_/B vssd1 vssd1 vccd1 vccd1 _12304_/B sky130_fd_sc_hd__or2_1
XFILLER_0_48_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12179_ _12170_/A _09059_/A _09059_/B _09163_/X vssd1 vssd1 vccd1 vccd1 _12180_/B
+ sky130_fd_sc_hd__a31o_1
XANTENNA__06678__B _12644_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06740_ _07100_/A reg1_val[10] vssd1 vssd1 vccd1 vccd1 _06740_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_64_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11458__A3 _11457_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06671_ _06702_/A _12654_/B vssd1 vssd1 vccd1 vccd1 _06671_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__10666__B2 _10818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10666__A1 _10963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08410_ _09423_/B2 _08744_/A2 _08564_/B _07955_/A vssd1 vssd1 vccd1 vccd1 _08411_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07531__A1 _07099_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09390_ _09214_/A _09213_/B _09211_/X vssd1 vssd1 vccd1 vccd1 _09391_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_80_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11615__B1 _12290_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08341_ _08343_/B _08343_/A vssd1 vssd1 vccd1 vccd1 _08341_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_117_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07295__B1 _11766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08272_ _08740_/A _08272_/B vssd1 vssd1 vccd1 vccd1 _08275_/A sky130_fd_sc_hd__xnor2_2
X_07223_ _07223_/A _07223_/B vssd1 vssd1 vccd1 vccd1 _07223_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_73_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout127_A _10022_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07154_ _07154_/A _07154_/B vssd1 vssd1 vccd1 vccd1 _07154_/X sky130_fd_sc_hd__and2_1
XFILLER_0_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07085_ _11269_/A _07090_/B _11261_/A vssd1 vssd1 vccd1 vccd1 _07087_/A sky130_fd_sc_hd__o21a_4
XFILLER_0_14_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout113 _08732_/A1 vssd1 vssd1 vccd1 vccd1 _11146_/A sky130_fd_sc_hd__buf_6
Xfanout102 _10422_/A vssd1 vssd1 vccd1 vccd1 _11261_/A sky130_fd_sc_hd__clkbuf_16
Xfanout146 _07036_/X vssd1 vssd1 vccd1 vccd1 _09768_/A1 sky130_fd_sc_hd__buf_8
Xfanout124 _12826_/A vssd1 vssd1 vccd1 vccd1 _10927_/A1 sky130_fd_sc_hd__clkbuf_8
Xfanout135 _12814_/A vssd1 vssd1 vccd1 vccd1 _10567_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout168 _07199_/Y vssd1 vssd1 vccd1 vccd1 _08584_/A sky130_fd_sc_hd__buf_8
Xfanout179 _09423_/B2 vssd1 vssd1 vccd1 vccd1 _07752_/B sky130_fd_sc_hd__buf_6
Xfanout157 _12426_/A vssd1 vssd1 vccd1 vccd1 _10748_/A sky130_fd_sc_hd__buf_2
X_07987_ _08925_/A _07987_/B vssd1 vssd1 vccd1 vccd1 _07989_/B sky130_fd_sc_hd__and2_1
X_06938_ _12423_/A _06939_/B vssd1 vssd1 vccd1 vccd1 _12404_/A sky130_fd_sc_hd__and2_4
X_09726_ _09726_/A _09726_/B vssd1 vssd1 vccd1 vccd1 _09791_/A sky130_fd_sc_hd__xnor2_4
X_06869_ _10752_/A _10629_/A _06869_/C _06869_/D vssd1 vssd1 vccd1 vccd1 _06873_/C
+ sky130_fd_sc_hd__or4_1
X_09657_ _12426_/A _09656_/C _09656_/B vssd1 vssd1 vccd1 vccd1 _09658_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_69_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13056__C1 _13128_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08608_ _08611_/A _08611_/B _08593_/Y vssd1 vssd1 vccd1 vccd1 _08697_/A sky130_fd_sc_hd__o21ai_1
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09588_ _09588_/A _09588_/B vssd1 vssd1 vccd1 vccd1 _09589_/B sky130_fd_sc_hd__and2_1
X_08539_ _08574_/A _08545_/B _08532_/X vssd1 vssd1 vccd1 vccd1 _08570_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_65_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09275__B2 _12820_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09275__A1 _07075_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11550_ curr_PC[18] _11550_/B vssd1 vssd1 vccd1 vccd1 _11734_/C sky130_fd_sc_hd__and2_2
XFILLER_0_108_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10501_ _11792_/A _10410_/Y _10500_/Y vssd1 vssd1 vccd1 vccd1 _10501_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout6_A fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13220_ _13220_/A _13220_/B vssd1 vssd1 vccd1 vccd1 _13220_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_80_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11481_ _12317_/A _11481_/B vssd1 vssd1 vccd1 vccd1 _11488_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__11909__A1 fanout24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11909__B2 _07819_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07038__B1 _09768_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08324__A _08745_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10432_ _10928_/A _10432_/B vssd1 vssd1 vccd1 vccd1 _10440_/A sky130_fd_sc_hd__xnor2_1
X_13151_ hold287/A _13150_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13151_/X sky130_fd_sc_hd__mux2_1
X_10363_ _10364_/A _10364_/B vssd1 vssd1 vccd1 vccd1 _10861_/D sky130_fd_sc_hd__or2_1
XFILLER_0_103_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13082_ hold73/X _06572_/A _06892_/B hold83/A rst vssd1 vssd1 vccd1 vccd1 hold74/A
+ sky130_fd_sc_hd__a221o_1
X_12102_ _12168_/B vssd1 vssd1 vccd1 vccd1 _12103_/B sky130_fd_sc_hd__inv_2
XFILLER_0_20_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12033_ _11959_/A _11956_/X _11973_/A vssd1 vssd1 vccd1 vccd1 _12033_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__06800__A3 _12634_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10294_ _10206_/B _10209_/B _10204_/Y vssd1 vssd1 vccd1 vccd1 _10303_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_18_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07761__B2 _10537_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07761__A1 _08432_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12935_ hold47/X hold277/X vssd1 vssd1 vccd1 vccd1 _13174_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_125_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12866_ hold29/X hold261/X vssd1 vssd1 vccd1 vccd1 _12866_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_87_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11817_ _11790_/Y _11791_/X _11793_/Y _09163_/X _11816_/X vssd1 vssd1 vccd1 vccd1
+ _11817_/X sky130_fd_sc_hd__o221a_1
X_12797_ _09251_/A _13077_/A2 hold133/X _13109_/A vssd1 vssd1 vccd1 vccd1 _13252_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11748_ _11989_/A fanout15/X fanout36/X _12067_/A vssd1 vssd1 vccd1 vccd1 _11749_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_83_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12455__S _12455_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11679_ _11575_/A _11575_/B _11580_/A vssd1 vssd1 vccd1 vccd1 _11685_/A sky130_fd_sc_hd__o21bai_2
XANTENNA__08234__A _08722_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13349_ _13383_/CLK _13349_/D vssd1 vssd1 vccd1 vccd1 hold240/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07910_ _07910_/A _07910_/B vssd1 vssd1 vccd1 vccd1 _07978_/B sky130_fd_sc_hd__xnor2_1
X_08890_ _08890_/A _08890_/B vssd1 vssd1 vccd1 vccd1 _08893_/A sky130_fd_sc_hd__and2_1
XFILLER_0_75_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07841_ _07840_/B _07840_/C _07840_/A vssd1 vssd1 vccd1 vccd1 _07910_/A sky130_fd_sc_hd__a21boi_1
X_07772_ _11385_/A _07772_/B vssd1 vssd1 vccd1 vccd1 _07776_/A sky130_fd_sc_hd__xnor2_1
X_06723_ reg1_val[13] _11020_/A vssd1 vssd1 vccd1 vccd1 _11021_/S sky130_fd_sc_hd__and2_1
X_09511_ _09504_/X _09510_/X _10119_/S vssd1 vssd1 vccd1 vccd1 _09532_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_79_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11836__B1 _11180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06654_ reg1_val[23] _07194_/A vssd1 vssd1 vccd1 vccd1 _06655_/B sky130_fd_sc_hd__and2b_1
X_09442_ _09442_/A _09443_/B vssd1 vssd1 vccd1 vccd1 _09442_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__08409__A _09433_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06585_ reg2_val[31] _06771_/A vssd1 vssd1 vccd1 vccd1 _06585_/X sky130_fd_sc_hd__and2_1
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09373_ curr_PC[0] curr_PC[1] vssd1 vssd1 vccd1 vccd1 _09373_/X sky130_fd_sc_hd__or2_1
XANTENNA__07313__A _07522_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13053__A2 _12818_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08324_ _08745_/A _08324_/B vssd1 vssd1 vccd1 vccd1 _08373_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07032__B _07037_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08255_ _08293_/A _08293_/B vssd1 vssd1 vccd1 vccd1 _08295_/B sky130_fd_sc_hd__and2_1
XANTENNA__10674__A _11261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10811__A1 fanout23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10811__B2 _11171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07206_ _07133_/A _07133_/B _07133_/C _06691_/B vssd1 vssd1 vccd1 vccd1 _07206_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08186_ _08742_/A _08186_/B vssd1 vssd1 vccd1 vccd1 _08241_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__08144__A _08728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07137_ _07169_/A _07140_/C _07142_/B _07142_/C _07223_/B vssd1 vssd1 vccd1 vccd1
+ _07138_/B sky130_fd_sc_hd__a41o_1
XFILLER_0_70_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07440__B1 _07282_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07068_ reg1_val[16] _07069_/B vssd1 vssd1 vccd1 vccd1 _07076_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_30_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09709_ _09486_/X _10097_/A _09708_/X vssd1 vssd1 vccd1 vccd1 _09810_/B sky130_fd_sc_hd__o21a_2
X_10981_ _10981_/A _10981_/B vssd1 vssd1 vccd1 vccd1 _10983_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_69_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12720_ _12725_/C _12720_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[18] sky130_fd_sc_hd__xnor2_4
XFILLER_0_85_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07223__A _07223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08319__A _08742_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12651_ _12651_/A _12651_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[5] sky130_fd_sc_hd__xor2_4
XANTENNA__10568__B _10959_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13044__A2 _12788_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11602_ _11603_/A _11603_/B _11603_/C vssd1 vssd1 vccd1 vccd1 _11700_/B sky130_fd_sc_hd__o21a_1
XANTENNA__08038__B _08038_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12582_ _12582_/A _12582_/B _12582_/C vssd1 vssd1 vccd1 vccd1 _12607_/A sky130_fd_sc_hd__and3_1
XANTENNA__12252__B1 _09354_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11533_ _11532_/A _11532_/B _11532_/C vssd1 vssd1 vccd1 vccd1 _11533_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_65_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11464_ _11465_/A _11465_/B vssd1 vssd1 vccd1 vccd1 _11466_/A sky130_fd_sc_hd__and2_1
XANTENNA__08054__A _08740_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13203_ hold265/A _13202_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13203_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_61_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10415_ _10415_/A _10415_/B vssd1 vssd1 vccd1 vccd1 _10416_/B sky130_fd_sc_hd__and2_1
XFILLER_0_110_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08223__A2 _08741_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11395_ _11396_/A _11396_/B vssd1 vssd1 vccd1 vccd1 _11397_/A sky130_fd_sc_hd__and2_1
XFILLER_0_0_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_534 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13134_ _12895_/X _13134_/B vssd1 vssd1 vccd1 vccd1 _13135_/B sky130_fd_sc_hd__nand2b_1
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10346_ _10346_/A _10346_/B vssd1 vssd1 vccd1 vccd1 _10360_/A sky130_fd_sc_hd__xor2_4
XANTENNA__10030__A2 fanout16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13065_ _07090_/B _13087_/B2 hold131/X vssd1 vssd1 vccd1 vccd1 _13335_/D sky130_fd_sc_hd__o21a_1
X_10277_ _10228_/A _10228_/B _10226_/X vssd1 vssd1 vccd1 vccd1 _10364_/A sky130_fd_sc_hd__a21o_2
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10318__B1 _08507_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12016_ _12093_/A _12014_/X _11932_/A _11933_/X vssd1 vssd1 vccd1 vccd1 _12016_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_45_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_0_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13285_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_88_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09613__A _09613_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12918_ _13092_/A _13092_/B _12915_/X vssd1 vssd1 vccd1 vccd1 _13097_/A sky130_fd_sc_hd__a21o_1
XANTENNA__06956__B _07064_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09239__A1 _07154_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08229__A _08740_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12849_ hold39/X _12848_/B _12848_/Y _13235_/A vssd1 vssd1 vccd1 vccd1 hold40/A sky130_fd_sc_hd__o211a_1
XFILLER_0_8_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06691__B _06691_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08462__A2 _08744_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08040_ _08041_/B _08041_/C _08731_/A vssd1 vssd1 vccd1 vccd1 _08042_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09991_ _09991_/A _09991_/B vssd1 vssd1 vccd1 vccd1 _09991_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_12_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10941__B _10941_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08942_ _08942_/A _08942_/B vssd1 vssd1 vccd1 vccd1 _08950_/A sky130_fd_sc_hd__xor2_4
XANTENNA__12214__A _12214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout194_A _09433_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07725__A1 _08741_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07725__B2 _08617_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08873_ _08847_/B _08849_/B _08847_/A vssd1 vssd1 vccd1 vccd1 _08878_/A sky130_fd_sc_hd__o21ba_1
XFILLER_0_98_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07824_ _07824_/A _07824_/B _07824_/C vssd1 vssd1 vccd1 vccd1 _07824_/X sky130_fd_sc_hd__and3_1
X_07755_ _07753_/Y _07754_/X _07856_/A _07856_/B vssd1 vssd1 vccd1 vccd1 _07759_/A
+ sky130_fd_sc_hd__a211o_1
X_06706_ reg1_val[16] _11343_/A vssd1 vssd1 vccd1 vccd1 _06707_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_79_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07686_ _09613_/A _07752_/B _07955_/A _09614_/A vssd1 vssd1 vccd1 vccd1 _07687_/B
+ sky130_fd_sc_hd__o22a_1
X_06637_ _07140_/B reg1_val[26] vssd1 vssd1 vccd1 vccd1 _12195_/S sky130_fd_sc_hd__and2b_1
XFILLER_0_79_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09425_ _09427_/A _09427_/B vssd1 vssd1 vccd1 vccd1 _09428_/A sky130_fd_sc_hd__nand2_1
XANTENNA__13026__A2 _12788_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11037__A1 _11171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09356_ hold244/A hold260/A _09835_/B vssd1 vssd1 vccd1 vccd1 _09356_/X sky130_fd_sc_hd__and3_1
X_06568_ hold72/X vssd1 vssd1 vccd1 vccd1 hold73/A sky130_fd_sc_hd__inv_2
XANTENNA__09669__S _09669_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11037__B2 fanout23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09287_ _09287_/A _09287_/B vssd1 vssd1 vccd1 vccd1 _09292_/A sky130_fd_sc_hd__nand2_4
XFILLER_0_74_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08307_ _08739_/A1 _08732_/A2 _08656_/B _08436_/A vssd1 vssd1 vccd1 vccd1 _08308_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_90_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07661__B1 _10022_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08238_ _08238_/A _08238_/B vssd1 vssd1 vccd1 vccd1 _08282_/B sky130_fd_sc_hd__xor2_1
XANTENNA__10796__B1 _07178_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11012__B _11012_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10200_ _11180_/A _10200_/B vssd1 vssd1 vccd1 vccd1 _10205_/A sky130_fd_sc_hd__xnor2_1
X_08169_ _08169_/A _08169_/B vssd1 vssd1 vccd1 vccd1 _08178_/A sky130_fd_sc_hd__xor2_1
X_11180_ _11180_/A _11180_/B vssd1 vssd1 vccd1 vccd1 _11181_/B sky130_fd_sc_hd__xnor2_1
X_10131_ reg1_val[6] curr_PC[6] vssd1 vssd1 vccd1 vccd1 _10132_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_100_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10062_ _10062_/A _10062_/B vssd1 vssd1 vccd1 vccd1 _10079_/A sky130_fd_sc_hd__nor2_2
XANTENNA__09433__A _09433_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06776__B _06960_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11276__A1 _10574_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11276__B2 _11751_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12703_ reg1_val[15] _12703_/B vssd1 vssd1 vccd1 vccd1 _12705_/C sky130_fd_sc_hd__xnor2_2
X_10964_ _10964_/A _10964_/B vssd1 vssd1 vccd1 vccd1 _10966_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__08141__B2 _10927_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08141__A1 _08730_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10895_ hold287/A _11341_/B _11017_/B _09837_/A vssd1 vssd1 vccd1 vccd1 _10896_/B
+ sky130_fd_sc_hd__a31o_1
XANTENNA__12794__A _12794_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11028__A1 _11876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12634_ reg1_val[2] _12634_/B vssd1 vssd1 vccd1 vccd1 _12635_/B sky130_fd_sc_hd__nand2_1
X_12565_ _12582_/A _12565_/B vssd1 vssd1 vccd1 vccd1 _12581_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_31_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11516_ _10622_/B _11102_/Y _11515_/B _11515_/X _11513_/X vssd1 vssd1 vccd1 vccd1
+ _11517_/B sky130_fd_sc_hd__a311o_4
XFILLER_0_25_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12496_ _12502_/B _12496_/B vssd1 vssd1 vccd1 vccd1 new_PC[7] sky130_fd_sc_hd__and2_4
XFILLER_0_80_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11447_ _06698_/X _11973_/B _11445_/Y _06700_/B _11446_/Y vssd1 vssd1 vccd1 vccd1
+ _11447_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_34_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10539__B1 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07404__B1 _12832_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11378_ _11378_/A _11378_/B vssd1 vssd1 vccd1 vccd1 _11381_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13117_ hold242/X _12789_/B _13116_/X _12790_/A vssd1 vssd1 vccd1 vccd1 hold243/A
+ sky130_fd_sc_hd__a22o_1
X_10329_ _10418_/A _10574_/A _10575_/A _11472_/A vssd1 vssd1 vccd1 vccd1 _10330_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13048_ hold134/X _12788_/A _13236_/B hold164/X _13109_/A vssd1 vssd1 vccd1 vccd1
+ hold165/A sky130_fd_sc_hd__o221a_1
XANTENNA__07707__A1 fanout69/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07707__B2 _08216_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06967__A _11020_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09343__A _09343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06686__B _12639_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07540_ _07540_/A _07540_/B _07540_/C _07540_/D vssd1 vssd1 vccd1 vccd1 _07541_/B
+ sky130_fd_sc_hd__or4_1
XANTENNA__08132__B2 _07752_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08132__A1 _07821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07471_ _09205_/B _07471_/B vssd1 vssd1 vccd1 vccd1 _07519_/A sky130_fd_sc_hd__and2_1
XFILLER_0_57_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09210_ _07478_/B _07481_/B _07478_/A vssd1 vssd1 vccd1 vccd1 _09210_/X sky130_fd_sc_hd__o21ba_1
XANTENNA__07891__B1 _08739_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09141_ reg1_val[6] reg1_val[25] _09142_/S vssd1 vssd1 vccd1 vccd1 _09141_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_8_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09072_ _09072_/A _09072_/B vssd1 vssd1 vccd1 vccd1 _09072_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__12209__A _12261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08023_ _08912_/A _08912_/B vssd1 vssd1 vccd1 vccd1 _08023_/X sky130_fd_sc_hd__or2_1
XANTENNA__07643__B1 _07819_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout4 fanout5/X vssd1 vssd1 vccd1 vccd1 fanout4/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_4_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09518__A _11886_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11742__A2 _12150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07946__B2 _08723_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07946__A1 _07896_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09974_ _09974_/A _09974_/B vssd1 vssd1 vccd1 vccd1 _09974_/X sky130_fd_sc_hd__or2_1
XFILLER_0_0_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08925_ _08925_/A _08925_/B vssd1 vssd1 vccd1 vccd1 _08930_/A sky130_fd_sc_hd__nand2_2
X_08856_ _08857_/A _08857_/B vssd1 vssd1 vccd1 vccd1 _08856_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_98_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07807_ _07807_/A _07807_/B vssd1 vssd1 vccd1 vccd1 _07809_/B sky130_fd_sc_hd__nand2_1
X_08787_ _08786_/B _08787_/B vssd1 vssd1 vccd1 vccd1 _08788_/B sky130_fd_sc_hd__and2b_1
XANTENNA__11258__A1 _09614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07738_ _07738_/A _07738_/B vssd1 vssd1 vccd1 vccd1 _07813_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__11258__B2 _09613_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07669_ _07669_/A _07669_/B vssd1 vssd1 vccd1 vccd1 _08944_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_48_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09408_ _09408_/A _09408_/B vssd1 vssd1 vccd1 vccd1 _09411_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_47_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07882__B1 _08436_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10680_ _10680_/A _10680_/B vssd1 vssd1 vccd1 vccd1 _10680_/X sky130_fd_sc_hd__xor2_1
XANTENNA_fanout22_A _07087_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09339_ _09332_/X _09338_/X _11010_/S vssd1 vssd1 vccd1 vccd1 _09339_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_82_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07220__B _07220_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12350_ _12429_/C _12349_/Y _12429_/B vssd1 vssd1 vccd1 vccd1 _12350_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_50_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12281_ _12281_/A _12281_/B vssd1 vssd1 vccd1 vccd1 _12380_/C sky130_fd_sc_hd__nor2_1
X_11301_ _11301_/A _11301_/B vssd1 vssd1 vccd1 vccd1 _11303_/C sky130_fd_sc_hd__xor2_1
X_11232_ _11232_/A vssd1 vssd1 vccd1 vccd1 _11232_/Y sky130_fd_sc_hd__inv_2
XANTENNA__09387__B1 _07089_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11163_ _11163_/A _11164_/B vssd1 vssd1 vccd1 vccd1 _11292_/A sky130_fd_sc_hd__and2_1
X_10114_ _09499_/X _09502_/X _10250_/S vssd1 vssd1 vccd1 vccd1 _10114_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_30_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11094_ _11095_/B _11095_/A vssd1 vssd1 vccd1 vccd1 _11210_/B sky130_fd_sc_hd__nand2b_1
X_10045_ _10046_/A _10046_/B vssd1 vssd1 vccd1 vccd1 _10045_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_26_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold60 hold60/A vssd1 vssd1 vccd1 vccd1 hold60/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 hold71/A vssd1 vssd1 vccd1 vccd1 hold71/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 hold82/A vssd1 vssd1 vccd1 vccd1 hold82/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13238__A2 _06892_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold93 hold93/A vssd1 vssd1 vccd1 vccd1 hold93/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_85_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08114__B2 _08739_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08114__A1 _08721_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11996_ _12317_/A _11996_/B vssd1 vssd1 vccd1 vccd1 _12005_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_98_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10947_ _10448_/A _10947_/B _10947_/C vssd1 vssd1 vccd1 vccd1 _10950_/B sky130_fd_sc_hd__nand3b_1
XANTENNA__07873__B1 _11766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10878_ _10879_/A _10879_/B vssd1 vssd1 vccd1 vccd1 _10878_/Y sky130_fd_sc_hd__nand2_1
X_12617_ _12623_/A _12617_/B vssd1 vssd1 vccd1 vccd1 _12618_/B sky130_fd_sc_hd__nor2_1
XANTENNA__08507__A _08673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07411__A _11163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12548_ _12703_/B _12548_/B vssd1 vssd1 vccd1 vccd1 _12549_/B sky130_fd_sc_hd__or2_1
XANTENNA__07130__B _11343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_2 _09984_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12479_ _12488_/A _12479_/B vssd1 vssd1 vccd1 vccd1 _12481_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_123_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10491__B _10493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07928__A1 _08752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07928__B2 _08798_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10932__B1 _12073_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06971_ _06971_/A _06971_/B vssd1 vssd1 vccd1 vccd1 _06971_/Y sky130_fd_sc_hd__nand2_2
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09690_ hold234/A _10391_/A2 _09688_/X _12401_/B1 vssd1 vssd1 vccd1 vccd1 _09690_/X
+ sky130_fd_sc_hd__a31o_1
X_08710_ _08710_/A _08710_/B vssd1 vssd1 vccd1 vccd1 _09021_/A sky130_fd_sc_hd__xnor2_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08641_ _08673_/A _09238_/B _09440_/B1 _08671_/B2 vssd1 vssd1 vccd1 vccd1 _08642_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_89_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08572_ _08572_/A _08572_/B vssd1 vssd1 vccd1 vccd1 _08589_/A sky130_fd_sc_hd__xnor2_1
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10012__A _10710_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07523_ _10574_/A _12810_/A _10413_/A _10575_/A vssd1 vssd1 vccd1 vccd1 _07524_/B
+ sky130_fd_sc_hd__o22a_1
X_07454_ _07561_/A _07561_/B vssd1 vssd1 vccd1 vccd1 _07562_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_36_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10463__A2 fanout48/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08408__A2 _08741_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07385_ _07385_/A _07385_/B vssd1 vssd1 vccd1 vccd1 _07386_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_115_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09124_ reg1_val[13] reg1_val[18] _09142_/S vssd1 vssd1 vccd1 vccd1 _09124_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_60_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_478 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09055_ _09055_/A vssd1 vssd1 vccd1 vccd1 _09055_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_44_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08006_ _08006_/A _08006_/B vssd1 vssd1 vccd1 vccd1 _08007_/B sky130_fd_sc_hd__and2_1
XFILLER_0_13_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08152__A _08722_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09957_ _09957_/A _09957_/B vssd1 vssd1 vccd1 vccd1 _09958_/B sky130_fd_sc_hd__nand2_2
X_08908_ _08904_/Y _09047_/B _08905_/X vssd1 vssd1 vccd1 vccd1 _09053_/A sky130_fd_sc_hd__o21ai_4
XANTENNA__09541__B1 _09538_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09888_ _09889_/A _09889_/B vssd1 vssd1 vccd1 vccd1 _10076_/A sky130_fd_sc_hd__nor2_1
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12140__A2 _12412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08839_ _09036_/B _09042_/A vssd1 vssd1 vccd1 vccd1 _08839_/X sky130_fd_sc_hd__and2_1
X_11850_ _11656_/Y _11769_/B _11767_/X vssd1 vssd1 vccd1 vccd1 _11853_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__09844__A1 _12394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10801_ _10800_/B _10800_/C _10800_/A vssd1 vssd1 vccd1 vccd1 _10802_/C sky130_fd_sc_hd__o21ai_1
X_11781_ _11781_/A vssd1 vssd1 vccd1 vccd1 _11783_/A sky130_fd_sc_hd__inv_2
XFILLER_0_67_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11651__A1 _09613_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10732_ _10733_/B _10733_/A vssd1 vssd1 vccd1 vccd1 _10858_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_48_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11651__B2 _09614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10663_ _10928_/A _10663_/B vssd1 vssd1 vccd1 vccd1 _10665_/A sky130_fd_sc_hd__xnor2_1
X_13382_ _13383_/CLK hold103/X vssd1 vssd1 vccd1 vccd1 hold101/A sky130_fd_sc_hd__dfxtp_1
X_12402_ _12402_/A0 _09165_/X _12402_/S vssd1 vssd1 vccd1 vccd1 _12402_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_51_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07607__B1 fanout66/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10594_ _10594_/A _10594_/B vssd1 vssd1 vccd1 vccd1 _10596_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_50_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12333_ _12222_/Y _12276_/X _12278_/B vssd1 vssd1 vccd1 vccd1 _12333_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__07885__B _07885_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09158__A _09168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12264_ _12264_/A _12264_/B vssd1 vssd1 vccd1 vccd1 _12266_/B sky130_fd_sc_hd__nand2_1
X_12195_ _12402_/A0 _09354_/B _12195_/S vssd1 vssd1 vccd1 vccd1 _12195_/X sky130_fd_sc_hd__mux2_1
X_11215_ _11215_/A _11423_/A vssd1 vssd1 vccd1 vccd1 _11215_/X sky130_fd_sc_hd__or2_1
XFILLER_0_128_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11146_ _11146_/A _12214_/B vssd1 vssd1 vccd1 vccd1 _11148_/B sky130_fd_sc_hd__or2_1
X_11077_ _11075_/X _11077_/B vssd1 vssd1 vccd1 vccd1 _11078_/B sky130_fd_sc_hd__and2b_1
X_10028_ _10147_/A _10028_/B vssd1 vssd1 vccd1 vccd1 _10029_/B sky130_fd_sc_hd__or2_1
XFILLER_0_53_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09621__A _10422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08099__B1 _08727_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11642__A1 _12247_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11979_ _09156_/Y _11958_/Y _11959_/X _11978_/Y _11954_/X vssd1 vssd1 vccd1 vccd1
+ _11979_/X sky130_fd_sc_hd__a311o_1
XFILLER_0_58_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07170_ _09238_/B _12842_/A _09440_/B1 _12844_/A vssd1 vssd1 vccd1 vccd1 _07171_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_42_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08271__B1 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13147__B2 _13246_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10905__B1 _10904_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout306 _06574_/Y vssd1 vssd1 vccd1 vccd1 _07149_/A sky130_fd_sc_hd__buf_8
X_09811_ _09811_/A _09811_/B vssd1 vssd1 vccd1 vccd1 _09853_/C sky130_fd_sc_hd__and2_1
XANTENNA__12107__C1 _09163_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09742_ _09742_/A _09742_/B vssd1 vssd1 vccd1 vccd1 _09743_/B sky130_fd_sc_hd__nand2_1
X_06954_ _10710_/A _06954_/B vssd1 vssd1 vccd1 vccd1 _06971_/B sky130_fd_sc_hd__nand2_1
X_09673_ _09517_/A _09514_/Y _09516_/B vssd1 vssd1 vccd1 vccd1 _09673_/X sky130_fd_sc_hd__o21a_1
X_06885_ dest_pred_val _06921_/B _06881_/X vssd1 vssd1 vccd1 vccd1 take_branch sky130_fd_sc_hd__a21o_4
XTAP_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06888__A1 _06771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08624_ _08625_/A _08625_/B vssd1 vssd1 vccd1 vccd1 _08624_/X sky130_fd_sc_hd__or2_1
XANTENNA__10684__A2 fanout30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08555_ _12804_/A _08661_/A2 _08673_/B _09768_/A1 vssd1 vssd1 vccd1 vccd1 _08556_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07506_ _09351_/B _12264_/B vssd1 vssd1 vccd1 vccd1 _07515_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_77_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07051__A _08632_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08486_ _08514_/A _08514_/B vssd1 vssd1 vccd1 vccd1 _08489_/B sky130_fd_sc_hd__and2b_1
XANTENNA__10436__A2 fanout30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_13_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13365_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_119_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07437_ _07437_/A _07437_/B vssd1 vssd1 vccd1 vccd1 _07563_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_18_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06890__A _12790_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07368_ _08671_/B2 fanout16/X _07282_/B _12798_/A vssd1 vssd1 vccd1 vccd1 _07369_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_18_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13199__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09107_ reg1_val[11] reg1_val[20] _09108_/S vssd1 vssd1 vccd1 vccd1 _09107_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_33_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07299_ _07999_/A _07999_/B vssd1 vssd1 vccd1 vccd1 _08000_/A sky130_fd_sc_hd__or2_4
XFILLER_0_102_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09038_ _09042_/A _09038_/B vssd1 vssd1 vccd1 vccd1 _11793_/A sky130_fd_sc_hd__xor2_2
XANTENNA__11020__B _12404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11000_ _11792_/A _10999_/B _10999_/C vssd1 vssd1 vccd1 vccd1 _11000_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__07368__A2 fanout16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12951_ _13215_/B _13216_/A _12864_/X vssd1 vssd1 vccd1 vccd1 _13220_/A sky130_fd_sc_hd__a21o_1
X_12882_ hold292/A hold25/X vssd1 vssd1 vccd1 vccd1 _13169_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_99_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11902_ curr_PC[22] _11982_/C _11901_/Y vssd1 vssd1 vccd1 vccd1 _11902_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_59_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09441__A _09441_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11833_ _11833_/A _11833_/B vssd1 vssd1 vccd1 vccd1 _11840_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_114_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07828__B1 _08752_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08057__A _08745_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11764_ _11764_/A _11764_/B vssd1 vssd1 vccd1 vccd1 _11777_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_28_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10715_ _10716_/A _10716_/B vssd1 vssd1 vccd1 vccd1 _10715_/Y sky130_fd_sc_hd__nand2b_1
X_11695_ _11697_/A _11697_/B _11697_/C vssd1 vssd1 vccd1 vccd1 _11698_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_126_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10646_ hold288/A _10646_/B vssd1 vssd1 vccd1 vccd1 _10769_/B sky130_fd_sc_hd__or2_1
XFILLER_0_70_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07896__A _07896_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13365_ _13365_/CLK _13365_/D vssd1 vssd1 vccd1 vccd1 hold263/A sky130_fd_sc_hd__dfxtp_1
X_10577_ _10576_/B _10576_/C _11180_/A vssd1 vssd1 vccd1 vccd1 _10579_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_24_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13296_ _13299_/CLK hold214/X vssd1 vssd1 vccd1 vccd1 hold212/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12316_ _12316_/A _12316_/B vssd1 vssd1 vccd1 vccd1 _12317_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_23_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12247_ hold256/A _09355_/X _12301_/B _12246_/Y _12247_/C1 vssd1 vssd1 vccd1 vccd1
+ _12247_/X sky130_fd_sc_hd__a311o_1
XFILLER_0_48_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09753__B1 _11751_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12178_ _12170_/A _09059_/A _09059_/B vssd1 vssd1 vccd1 vccd1 _12180_/A sky130_fd_sc_hd__a21oi_1
X_11129_ hold228/A _11450_/B _11236_/B _11968_/B1 vssd1 vssd1 vccd1 vccd1 _11129_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_3_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06670_ instruction[0] instruction[1] instruction[2] instruction[31] pred_val vssd1
+ vssd1 vccd1 vccd1 _12654_/B sky130_fd_sc_hd__o311a_4
XFILLER_0_64_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10666__A2 _10797_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09351__A _12388_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06975__A _10707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07531__A2 _07099_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08340_ _08340_/A _08340_/B vssd1 vssd1 vccd1 vccd1 _08343_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_117_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07295__B2 _09568_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07295__A1 _09567_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08271_ _07955_/A fanout87/X fanout82/X _07896_/A vssd1 vssd1 vccd1 vccd1 _08272_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_117_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07222_ _10321_/A _10320_/A vssd1 vssd1 vccd1 vccd1 _07222_/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_61_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07153_ _07343_/B _07223_/B _07151_/B _06838_/B vssd1 vssd1 vccd1 vccd1 _07154_/B
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__11379__B1 _12067_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11121__A _12394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07084_ reg1_val[20] _07084_/B vssd1 vssd1 vccd1 vccd1 _07090_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__10051__B1 _11751_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09744__B1 _10418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout103 _11758_/A vssd1 vssd1 vccd1 vccd1 _10422_/A sky130_fd_sc_hd__buf_12
XFILLER_0_1_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11551__B1 _11142_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout147 _12804_/A vssd1 vssd1 vccd1 vccd1 _07896_/A sky130_fd_sc_hd__buf_6
Xfanout125 _10537_/A1 vssd1 vssd1 vccd1 vccd1 _10445_/A sky130_fd_sc_hd__clkbuf_8
Xfanout136 _12814_/A vssd1 vssd1 vccd1 vccd1 _08436_/A sky130_fd_sc_hd__buf_6
Xfanout114 _12824_/A vssd1 vssd1 vccd1 vccd1 _08732_/A1 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout169 _09568_/B vssd1 vssd1 vccd1 vccd1 _08617_/B sky130_fd_sc_hd__buf_8
Xfanout158 _08980_/Y vssd1 vssd1 vccd1 vccd1 _12426_/A sky130_fd_sc_hd__clkbuf_4
X_07986_ _07986_/A _07986_/B _07986_/C vssd1 vssd1 vccd1 vccd1 _07987_/B sky130_fd_sc_hd__or3_1
X_06937_ _09163_/A _09159_/B vssd1 vssd1 vccd1 vccd1 _06939_/B sky130_fd_sc_hd__nor2_2
X_09725_ _09726_/B _09726_/A vssd1 vssd1 vccd1 vccd1 _09725_/Y sky130_fd_sc_hd__nand2b_1
X_09656_ _12426_/A _09656_/B _09656_/C vssd1 vssd1 vccd1 vccd1 _09658_/B sky130_fd_sc_hd__or3_1
X_06868_ _11224_/A _11111_/A _11004_/A _10879_/A vssd1 vssd1 vccd1 vccd1 _06869_/D
+ sky130_fd_sc_hd__or4_1
X_08607_ _08607_/A vssd1 vssd1 vccd1 vccd1 _08611_/B sky130_fd_sc_hd__inv_2
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06799_ reg2_val[1] _06799_/B vssd1 vssd1 vccd1 vccd1 _06799_/X sky130_fd_sc_hd__and2_2
XFILLER_0_77_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09587_ _09588_/A _09588_/B vssd1 vssd1 vccd1 vccd1 _09732_/B sky130_fd_sc_hd__nor2_1
X_08538_ _08538_/A _08538_/B vssd1 vssd1 vccd1 vccd1 _08545_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_77_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09275__A2 _11653_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10200__A _11180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08469_ _08469_/A _08469_/B vssd1 vssd1 vccd1 vccd1 _08483_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_49_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10500_ _10739_/A _10500_/B vssd1 vssd1 vccd1 vccd1 _10500_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_0_9_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07038__A1 _12804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11480_ _11766_/A fanout15/X fanout36/X _11847_/A vssd1 vssd1 vccd1 vccd1 _11481_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11909__A2 fanout12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07038__B2 _10575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10431_ _10818_/A fanout16/X _07282_/B _10963_/A vssd1 vssd1 vccd1 vccd1 _10432_/B
+ sky130_fd_sc_hd__o22a_1
X_13150_ _13150_/A _13150_/B vssd1 vssd1 vccd1 vccd1 _13150_/Y sky130_fd_sc_hd__xnor2_1
X_10362_ _10364_/A _10364_/B vssd1 vssd1 vccd1 vccd1 _10861_/C sky130_fd_sc_hd__nand2_1
X_13081_ _07263_/B _13087_/B2 hold129/X vssd1 vssd1 vccd1 vccd1 _13343_/D sky130_fd_sc_hd__o21a_1
XANTENNA__10870__A _11100_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12101_ _12226_/A _12101_/B vssd1 vssd1 vccd1 vccd1 _12168_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_21_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10293_ _10293_/A _10293_/B vssd1 vssd1 vccd1 vccd1 _10346_/A sky130_fd_sc_hd__and2_2
X_12032_ _12031_/A _12031_/B _12031_/C vssd1 vssd1 vccd1 vccd1 _12032_/Y sky130_fd_sc_hd__o21ai_1
Xhold190 hold190/A vssd1 vssd1 vccd1 vccd1 hold190/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07761__A2 _08741_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12934_ _13169_/B _13170_/A _12881_/X vssd1 vssd1 vccd1 vccd1 _13175_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_125_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12865_ hold281/A hold39/X vssd1 vssd1 vccd1 vccd1 _13215_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_34_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12796_ hold132/X _12798_/B vssd1 vssd1 vccd1 vccd1 hold133/A sky130_fd_sc_hd__or2_1
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11816_ _11624_/A _11797_/Y _11804_/X _11815_/X vssd1 vssd1 vccd1 vccd1 _11816_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_68_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11747_ _11750_/A vssd1 vssd1 vccd1 vccd1 _11747_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_126_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10281__B1 _10575_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09110__S _09111_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11678_ _11561_/Y _11570_/B _11583_/A vssd1 vssd1 vccd1 vccd1 _11689_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_126_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10629_ _10629_/A _10629_/B vssd1 vssd1 vccd1 vccd1 _10629_/Y sky130_fd_sc_hd__nand2_1
X_13348_ _13383_/CLK _13348_/D vssd1 vssd1 vccd1 vccd1 hold244/A sky130_fd_sc_hd__dfxtp_2
XANTENNA__10033__B1 _10148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11876__A _11876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13279_ _13357_/CLK _13279_/D vssd1 vssd1 vccd1 vccd1 hold140/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06689__B _07131_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07840_ _07840_/A _07840_/B _07840_/C vssd1 vssd1 vccd1 vccd1 _08026_/A sky130_fd_sc_hd__and3_1
X_07771_ fanout69/X _08721_/B1 _08739_/A1 _08216_/B vssd1 vssd1 vccd1 vccd1 _07772_/B
+ sky130_fd_sc_hd__o22a_1
X_06722_ _11020_/A reg1_val[13] vssd1 vssd1 vccd1 vccd1 _06722_/Y sky130_fd_sc_hd__nand2b_1
X_09510_ _09507_/X _09509_/X _11010_/S vssd1 vssd1 vccd1 vccd1 _09510_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_79_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11836__A1 _11261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06653_ _07194_/A reg1_val[23] vssd1 vssd1 vccd1 vccd1 _11973_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_91_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09441_ _09441_/A _09441_/B vssd1 vssd1 vccd1 vccd1 _09443_/B sky130_fd_sc_hd__xnor2_2
X_06584_ instruction[0] instruction[2] instruction[1] pred_val vssd1 vssd1 vccd1 vccd1
+ _06584_/X sky130_fd_sc_hd__or4bb_1
XFILLER_0_93_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09372_ _11142_/S _09372_/B vssd1 vssd1 vccd1 vccd1 _09372_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_117_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08465__B1 _09568_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08323_ _07896_/A _08744_/A2 _10022_/B1 _08723_/B1 vssd1 vssd1 vccd1 vccd1 _08324_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_19_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10811__A2 _10574_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08254_ _08254_/A _08254_/B vssd1 vssd1 vccd1 vccd1 _08293_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_105_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07205_ _06961_/Y _06966_/Y _07129_/X _07223_/B vssd1 vssd1 vccd1 vccd1 _07205_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_6_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08185_ _08436_/A _08741_/A2 _08617_/B fanout99/X vssd1 vssd1 vccd1 vccd1 _08186_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08217__A0 _11385_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07136_ _07142_/B _07142_/C _07223_/B vssd1 vssd1 vccd1 vccd1 _07166_/B sky130_fd_sc_hd__a21oi_1
X_07067_ _07067_/A _07067_/B vssd1 vssd1 vccd1 vccd1 _12816_/A sky130_fd_sc_hd__and2_4
XANTENNA__06779__B1 _06778_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07440__A1 _09423_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07440__B2 _12802_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06794__A3 _12639_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06599__B _07064_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09708_ _09482_/X _09645_/X _09646_/X vssd1 vssd1 vccd1 vccd1 _09708_/X sky130_fd_sc_hd__a21o_1
X_07969_ _07969_/A _07969_/B _07969_/C vssd1 vssd1 vccd1 vccd1 _07974_/A sky130_fd_sc_hd__or3_1
XFILLER_0_4_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10980_ _10981_/B _10981_/A vssd1 vssd1 vccd1 vccd1 _10980_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_85_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09639_ _09639_/A _09639_/B vssd1 vssd1 vccd1 vccd1 _09641_/B sky130_fd_sc_hd__xnor2_4
X_12650_ _12648_/Y _12650_/B vssd1 vssd1 vccd1 vccd1 _12651_/B sky130_fd_sc_hd__nand2b_2
XANTENNA__12252__A1 _07144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11601_ _11601_/A _11601_/B vssd1 vssd1 vccd1 vccd1 _11603_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__08038__C _08038_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12581_ _12581_/A _12581_/B _12581_/C vssd1 vssd1 vccd1 vccd1 _12605_/A sky130_fd_sc_hd__or3_1
XFILLER_0_93_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11532_ _11532_/A _11532_/B _11532_/C vssd1 vssd1 vccd1 vccd1 _11532_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_80_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11463_ _11758_/A _11463_/B vssd1 vssd1 vccd1 vccd1 _11465_/B sky130_fd_sc_hd__xnor2_1
X_13202_ _13202_/A _13202_/B vssd1 vssd1 vccd1 vccd1 _13202_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_61_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10414_ _10413_/A _12316_/B _10413_/C _10413_/D vssd1 vssd1 vccd1 vccd1 _10415_/B
+ sky130_fd_sc_hd__o22ai_1
X_13133_ _13235_/A hold289/X vssd1 vssd1 vccd1 vccd1 _13356_/D sky130_fd_sc_hd__and2_1
XFILLER_0_110_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_773 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11394_ _11394_/A _11394_/B vssd1 vssd1 vccd1 vccd1 _11396_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_21_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10345_ _10345_/A _10345_/B vssd1 vssd1 vccd1 vccd1 _10346_/B sky130_fd_sc_hd__nor2_2
X_13064_ hold99/X _12791_/A _13080_/B1 hold130/X _13128_/A vssd1 vssd1 vccd1 vccd1
+ hold131/A sky130_fd_sc_hd__o221a_1
X_10276_ _10658_/A _11033_/A vssd1 vssd1 vccd1 vccd1 _10410_/A sky130_fd_sc_hd__or2_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10318__B2 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10318__A1 _09568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12015_ _11932_/A _11933_/X _12093_/A _12014_/X vssd1 vssd1 vccd1 vccd1 _12093_/B
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__07195__B1 _09568_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10759__B _11886_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09613__B _10818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12917_ hold70/X hold59/X vssd1 vssd1 vccd1 vccd1 _13092_/B sky130_fd_sc_hd__nand2b_1
X_12848_ _12848_/A _12848_/B vssd1 vssd1 vccd1 vccd1 _12848_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_69_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09239__A2 _07154_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12779_ _12779_/A _12779_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[30] sky130_fd_sc_hd__xnor2_4
XFILLER_0_29_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09990_ _09988_/Y _09990_/B vssd1 vssd1 vccd1 vccd1 _09991_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_3_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08941_ _08932_/A _08932_/B _08933_/Y vssd1 vssd1 vccd1 vccd1 _08951_/A sky130_fd_sc_hd__o21ai_4
XFILLER_0_110_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12214__B _12214_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08872_ _08872_/A _08872_/B vssd1 vssd1 vccd1 vccd1 _08880_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__07725__A2 _11472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07823_ _07822_/B _07822_/C _11908_/A vssd1 vssd1 vccd1 vccd1 _07824_/C sky130_fd_sc_hd__a21o_1
XANTENNA_fanout187_A _09431_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07754_ _07753_/B _07753_/C _11908_/A vssd1 vssd1 vccd1 vccd1 _07754_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06705_ _11343_/A reg1_val[16] vssd1 vssd1 vccd1 vccd1 _06705_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_79_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07685_ _07685_/A _07685_/B vssd1 vssd1 vccd1 vccd1 _09706_/A sky130_fd_sc_hd__xnor2_4
X_06636_ reg2_val[26] _06771_/A _06596_/Y _06635_/Y vssd1 vssd1 vccd1 vccd1 _07140_/B
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_94_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09424_ _12264_/B _09424_/B vssd1 vssd1 vccd1 vccd1 _09427_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09355_ hold61/A _12341_/A vssd1 vssd1 vccd1 vccd1 _09355_/X sky130_fd_sc_hd__and2_1
X_06567_ hold82/X vssd1 vssd1 vccd1 vccd1 hold83/A sky130_fd_sc_hd__inv_2
XANTENNA__12234__A1 _12423_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08438__B1 _08731_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11037__A2 fanout48/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10685__A _12076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09286_ _07560_/A _07559_/B _07557_/Y vssd1 vssd1 vccd1 vccd1 _09296_/A sky130_fd_sc_hd__a21o_2
XFILLER_0_62_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07110__B1 _10575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08306_ _08370_/A _08370_/B vssd1 vssd1 vccd1 vccd1 _08327_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_34_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07661__A1 _11367_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08237_ _08238_/A _08238_/B vssd1 vssd1 vccd1 vccd1 _08237_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_105_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07661__B2 _09745_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08168_ _08253_/A _08253_/B _08160_/Y vssd1 vssd1 vccd1 vccd1 _08211_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_113_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07119_ reg1_val[3] _07120_/B vssd1 vssd1 vccd1 vccd1 _09594_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08099_ _10927_/A1 _08727_/A2 _08727_/B1 _11367_/A vssd1 vssd1 vccd1 vccd1 _08100_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_101_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10130_ reg1_val[6] curr_PC[6] vssd1 vssd1 vccd1 vccd1 _10130_/Y sky130_fd_sc_hd__nor2_1
X_10061_ _10061_/A _10061_/B vssd1 vssd1 vccd1 vccd1 _10062_/B sky130_fd_sc_hd__nor2_1
XANTENNA__09714__A _10928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11276__A2 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10963_ _10963_/A _12316_/B vssd1 vssd1 vccd1 vccd1 _10964_/B sky130_fd_sc_hd__or2_1
X_12702_ _12705_/B _12702_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[14] sky130_fd_sc_hd__and2_4
XANTENNA__08141__A2 _11367_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10894_ _11341_/B _11017_/B hold287/A vssd1 vssd1 vccd1 vccd1 _10896_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_38_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06792__B _06799_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12633_ reg1_val[2] _12634_/B vssd1 vssd1 vccd1 vccd1 _12633_/Y sky130_fd_sc_hd__nor2_1
X_12564_ _12623_/A _12564_/B vssd1 vssd1 vccd1 vccd1 _12565_/B sky130_fd_sc_hd__or2_1
XFILLER_0_65_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08065__A _08724_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11515_ _11515_/A _11515_/B vssd1 vssd1 vccd1 vccd1 _11515_/X sky130_fd_sc_hd__and2_1
XFILLER_0_25_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12495_ _12495_/A _12495_/B _12495_/C vssd1 vssd1 vccd1 vccd1 _12496_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_40_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11446_ _07130_/A _11343_/B _12455_/S vssd1 vssd1 vccd1 vccd1 _11446_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_1_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10539__A1 fanout94/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10539__B2 _10941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07404__B2 _10706_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07404__A1 _10445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12315__A _12316_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11377_ _11377_/A _11377_/B vssd1 vssd1 vccd1 vccd1 _11378_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_21_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13116_ hold258/A _13115_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13116_/X sky130_fd_sc_hd__mux2_1
XANTENNA__06758__A3 _12664_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10328_ _10328_/A _10328_/B vssd1 vssd1 vccd1 vccd1 _10341_/A sky130_fd_sc_hd__xnor2_1
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13047_ _10444_/A _13087_/B2 hold135/X vssd1 vssd1 vccd1 vccd1 hold136/A sky130_fd_sc_hd__o21a_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10259_ _07080_/A _12404_/A _12403_/A1 _06760_/Y vssd1 vssd1 vccd1 vccd1 _10259_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_56_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07707__A2 _10413_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06967__B _07074_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07144__A _07144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_56 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08132__A2 fanout69/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07470_ _07470_/A _07470_/B vssd1 vssd1 vccd1 vccd1 _07471_/B sky130_fd_sc_hd__or2_1
XANTENNA__06983__A _10448_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07891__A1 fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07891__B2 _08304_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09140_ _09138_/X _09139_/X _09336_/S vssd1 vssd1 vccd1 vccd1 _09140_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_57_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09071_ _08952_/Y _08963_/X _08964_/X vssd1 vssd1 vccd1 vccd1 _09071_/X sky130_fd_sc_hd__a21o_1
XANTENNA__07643__A1 _12798_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08022_ _08022_/A _08022_/B vssd1 vssd1 vccd1 vccd1 _08912_/B sky130_fd_sc_hd__xor2_2
XANTENNA__07643__B2 _09423_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout5 fanout5/A vssd1 vssd1 vccd1 vccd1 fanout5/X sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout102_A _10422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09973_ _11231_/S _09969_/X _09972_/Y _11233_/S vssd1 vssd1 vccd1 vccd1 _09973_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_40_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07946__A2 fanout69/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08924_ _08008_/A _08008_/B _08007_/A vssd1 vssd1 vccd1 vccd1 _08934_/A sky130_fd_sc_hd__a21o_1
X_08855_ _08853_/A _08853_/B _08857_/B vssd1 vssd1 vccd1 vccd1 _08855_/X sky130_fd_sc_hd__o21ba_1
X_08786_ _08787_/B _08786_/B vssd1 vssd1 vccd1 vccd1 _08786_/Y sky130_fd_sc_hd__nand2b_1
X_07806_ _07807_/A _07806_/B _07806_/C vssd1 vssd1 vccd1 vccd1 _07807_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_79_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07054__A _09716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07737_ _08722_/A _07737_/B vssd1 vssd1 vccd1 vccd1 _07813_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__11258__A2 _12150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10466__B1 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07668_ _07666_/A _07666_/B _07667_/X vssd1 vssd1 vccd1 vccd1 _08944_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_1_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06619_ _06621_/B vssd1 vssd1 vccd1 vccd1 _06619_/Y sky130_fd_sc_hd__inv_2
X_07599_ _07599_/A _07599_/B vssd1 vssd1 vccd1 vccd1 _07681_/A sky130_fd_sc_hd__xnor2_4
X_09407_ _10422_/A _09407_/B vssd1 vssd1 vccd1 vccd1 _09408_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_48_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07882__A1 _08432_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07882__B2 _10537_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09338_ _09334_/X _09974_/B _09974_/A vssd1 vssd1 vccd1 vccd1 _09338_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_63_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout15_A fanout16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07220__C _07220_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09269_ _09400_/A _10664_/A vssd1 vssd1 vccd1 vccd1 _09270_/C sky130_fd_sc_hd__or2_1
XANTENNA__11430__A2 _11649_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11300_ _11187_/A _11184_/B _11182_/X vssd1 vssd1 vccd1 vccd1 _11301_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_105_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12280_ _12280_/A _12414_/A vssd1 vssd1 vccd1 vccd1 _12281_/B sky130_fd_sc_hd__or2_1
XFILLER_0_15_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11231_ _10248_/X _10250_/X _11231_/S vssd1 vssd1 vccd1 vccd1 _11232_/A sky130_fd_sc_hd__mux2_1
XANTENNA__09387__A1 fanout30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09387__B2 _07688_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11162_ _11564_/A _11162_/B vssd1 vssd1 vccd1 vccd1 _11164_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_101_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10113_ _10113_/A _10113_/B vssd1 vssd1 vccd1 vccd1 _10113_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__12789__B _12789_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11093_ _10979_/A _10979_/B _10980_/X vssd1 vssd1 vccd1 vccd1 _11095_/B sky130_fd_sc_hd__o21ba_1
Xhold50 hold50/A vssd1 vssd1 vccd1 vccd1 hold50/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09444__A _09444_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10044_ _10192_/B _10044_/B vssd1 vssd1 vccd1 vccd1 _10046_/B sky130_fd_sc_hd__and2_1
Xhold61 hold61/A vssd1 vssd1 vccd1 vccd1 hold61/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 hold83/A vssd1 vssd1 vccd1 vccd1 hold83/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 hold72/A vssd1 vssd1 vccd1 vccd1 hold72/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09163__B _09170_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold94 hold94/A vssd1 vssd1 vccd1 vccd1 hold94/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07570__A0 _07504_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_49 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08114__A2 fanout87/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11995_ _12213_/A fanout15/X fanout36/X fanout56/X vssd1 vssd1 vccd1 vccd1 _11996_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_85_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10946_ _10947_/B _10947_/C _10448_/A vssd1 vssd1 vccd1 vccd1 _10950_/A sky130_fd_sc_hd__a21bo_1
X_10877_ _06819_/X _10876_/X _12174_/S vssd1 vssd1 vccd1 vccd1 _10879_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_39_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07873__B2 _08727_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07873__A1 _08727_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12616_ _12623_/A _12617_/B vssd1 vssd1 vccd1 vccd1 _12618_/A sky130_fd_sc_hd__and2_1
XANTENNA__08507__B _08507_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12547_ _12703_/B _12548_/B vssd1 vssd1 vccd1 vccd1 _12556_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_81_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_3 _10258_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12478_ _12649_/B _12478_/B vssd1 vssd1 vccd1 vccd1 _12479_/B sky130_fd_sc_hd__or2_1
XANTENNA__08523__A _08733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11429_ _11874_/A _11361_/B _11428_/Y _12290_/A vssd1 vssd1 vccd1 vccd1 _11429_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_6_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07928__A2 _09613_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06970_ _11343_/A _06968_/X _06969_/Y _07074_/B vssd1 vssd1 vccd1 vccd1 _12826_/A
+ sky130_fd_sc_hd__a22o_4
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06697__B _07130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08640_ _08636_/B _08636_/C _08636_/A vssd1 vssd1 vccd1 vccd1 _08643_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_83_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09838__C1 _09837_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08571_ _08571_/A _08571_/B _08571_/C vssd1 vssd1 vccd1 vccd1 _08703_/A sky130_fd_sc_hd__nor3_1
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07522_ _07522_/A _07522_/B vssd1 vssd1 vccd1 vccd1 _07526_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__11645__C1 _11644_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07453_ _07453_/A _07453_/B vssd1 vssd1 vccd1 vccd1 _07561_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_64_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09123_ reg1_val[12] reg1_val[19] _09142_/S vssd1 vssd1 vccd1 vccd1 _09123_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_84_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07384_ _07385_/A _07385_/B vssd1 vssd1 vccd1 vccd1 _07453_/A sky130_fd_sc_hd__and2_1
XFILLER_0_45_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10963__A _10963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09054_ _08910_/A _08903_/B _08910_/B vssd1 vssd1 vccd1 vccd1 _09055_/A sky130_fd_sc_hd__a21boi_1
XFILLER_0_32_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08005_ _08006_/A _08006_/B vssd1 vssd1 vccd1 vccd1 _08007_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_4_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09963__S _12388_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xmax_cap261 _09593_/A vssd1 vssd1 vccd1 vccd1 _08645_/A sky130_fd_sc_hd__buf_6
XFILLER_0_4_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09956_ _10496_/A _09956_/B _09956_/C vssd1 vssd1 vccd1 vccd1 _09957_/B sky130_fd_sc_hd__nand3_1
XANTENNA__09264__A _11065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09887_ _09755_/A _09755_/B _09752_/A vssd1 vssd1 vccd1 vccd1 _09889_/B sky130_fd_sc_hd__a21oi_2
X_08907_ _09033_/A _08839_/X _08886_/X _08887_/X _08906_/Y vssd1 vssd1 vccd1 vccd1
+ _09047_/B sky130_fd_sc_hd__a311oi_4
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08838_ _08838_/A _08838_/B vssd1 vssd1 vccd1 vccd1 _09042_/A sky130_fd_sc_hd__xor2_2
X_08769_ _08138_/A _08138_/B _08134_/Y vssd1 vssd1 vccd1 vccd1 _08775_/A sky130_fd_sc_hd__a21bo_1
X_10800_ _10800_/A _10800_/B _10800_/C vssd1 vssd1 vccd1 vccd1 _10913_/C sky130_fd_sc_hd__or3_2
X_11780_ _11782_/A _11782_/B _11782_/C vssd1 vssd1 vccd1 vccd1 _11781_/A sky130_fd_sc_hd__a21o_1
XANTENNA__09844__A2 _06924_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07512__A _12264_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10731_ _10731_/A _10731_/B vssd1 vssd1 vccd1 vccd1 _10733_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_94_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11651__A2 _12316_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12401_ hold215/A _12434_/B1 _12399_/X _12401_/B1 vssd1 vssd1 vccd1 vccd1 _12401_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_48_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10662_ _11065_/A fanout15/X fanout36/X _11146_/A vssd1 vssd1 vccd1 vccd1 _10663_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13381_ _13383_/CLK _13381_/D vssd1 vssd1 vccd1 vccd1 hold299/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07607__A1 _09768_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07607__B2 _12808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10593_ _10594_/A _10594_/B vssd1 vssd1 vccd1 vccd1 _10722_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_106_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12332_ _12332_/A _12334_/B vssd1 vssd1 vccd1 vccd1 _12332_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_106_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12263_ _12263_/A _12263_/B vssd1 vssd1 vccd1 vccd1 _12266_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_23_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11214_ _10988_/A _10988_/B _10989_/Y _11318_/A _11212_/Y vssd1 vssd1 vccd1 vccd1
+ _11214_/X sky130_fd_sc_hd__a41o_1
X_12194_ _12194_/A _12194_/B vssd1 vssd1 vccd1 vccd1 _12194_/Y sky130_fd_sc_hd__nor2_1
X_11145_ _11059_/A _11059_/B _11056_/A vssd1 vssd1 vccd1 vccd1 _11148_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__10127__C1 _10126_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07791__B1 _08617_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11076_ _11076_/A _11076_/B _11076_/C _11076_/D vssd1 vssd1 vccd1 vccd1 _11077_/B
+ sky130_fd_sc_hd__or4_1
XANTENNA__10678__B1 _12067_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10027_ _10027_/A _10027_/B vssd1 vssd1 vccd1 vccd1 _10028_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_53_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09902__A _10448_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11978_ _06924_/X _11965_/X _11977_/X vssd1 vssd1 vccd1 vccd1 _11978_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_98_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08099__B2 _11367_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08099__A1 _10927_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07422__A _09442_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10929_ _07048_/A _07048_/B _10575_/B vssd1 vssd1 vccd1 vccd1 _10931_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_128_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08271__A1 _07955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13147__A2 _06890_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08271__B2 _07896_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout307 reg1_val[1] vssd1 vssd1 vccd1 vccd1 _09343_/A sky130_fd_sc_hd__buf_8
X_09810_ _09810_/A _09810_/B _10368_/A vssd1 vssd1 vccd1 vccd1 _09811_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_10_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09084__A _12423_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09741_ _09741_/A _09741_/B vssd1 vssd1 vccd1 vccd1 _09742_/B sky130_fd_sc_hd__nand2_1
X_06953_ _10710_/A _06954_/B vssd1 vssd1 vccd1 vccd1 _06971_/A sky130_fd_sc_hd__or2_1
X_06884_ instruction[1] instruction[2] instruction[0] pred_val vssd1 vssd1 vccd1 vccd1
+ _06884_/Y sky130_fd_sc_hd__nand4b_4
XFILLER_0_118_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09672_ _09665_/X _09671_/X _10119_/S vssd1 vssd1 vccd1 vccd1 _09672_/X sky130_fd_sc_hd__mux2_2
XANTENNA__10023__A _10449_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08623_ _08625_/A _08625_/B vssd1 vssd1 vccd1 vccd1 _08623_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_27_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13083__A1 _09548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08554_ _08558_/A _08558_/B vssd1 vssd1 vccd1 vccd1 _08554_/Y sky130_fd_sc_hd__nor2_1
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout267_A _06881_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07505_ instruction[7] _07503_/X reg1_val[31] vssd1 vssd1 vccd1 vccd1 _12412_/B sky130_fd_sc_hd__a21bo_4
X_08485_ _08485_/A _08485_/B vssd1 vssd1 vccd1 vccd1 _08514_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_49_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07436_ _10449_/A _07436_/B vssd1 vssd1 vccd1 vccd1 _07437_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_9_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07367_ _12794_/A fanout9/A vssd1 vssd1 vccd1 vccd1 _07570_/S sky130_fd_sc_hd__nor2_1
XFILLER_0_33_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09106_ _09102_/X _09105_/X _09663_/S vssd1 vssd1 vccd1 vccd1 _09106_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_72_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07298_ _10449_/A _07298_/B vssd1 vssd1 vccd1 vccd1 _07999_/B sky130_fd_sc_hd__xnor2_1
X_09037_ _09032_/B _09036_/Y _09043_/A vssd1 vssd1 vccd1 vccd1 _09038_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_33_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_80 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout82_A _08507_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07773__B1 _08752_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09939_ _09939_/A _09939_/B vssd1 vssd1 vccd1 vccd1 _09940_/B sky130_fd_sc_hd__xor2_4
X_12950_ _12868_/B _13211_/B _12866_/X vssd1 vssd1 vccd1 vccd1 _13216_/A sky130_fd_sc_hd__a21o_1
X_12881_ hold25/X hold292/A vssd1 vssd1 vccd1 vccd1 _12881_/X sky130_fd_sc_hd__and2b_1
X_11901_ curr_PC[22] _11982_/C _12448_/S vssd1 vssd1 vccd1 vccd1 _11901_/Y sky130_fd_sc_hd__a21oi_1
X_11832_ _11918_/A _11832_/B vssd1 vssd1 vccd1 vccd1 _11833_/B sky130_fd_sc_hd__or2_1
XTAP_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07828__A1 _07752_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07828__B2 _07955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11763_ _11763_/A _11763_/B vssd1 vssd1 vccd1 vccd1 _11764_/B sky130_fd_sc_hd__or2_1
XTAP_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10714_ _10714_/A _10714_/B vssd1 vssd1 vccd1 vccd1 _10716_/B sky130_fd_sc_hd__xor2_2
X_11694_ _11782_/B _11694_/B vssd1 vssd1 vccd1 vccd1 _11697_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_126_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10645_ _12307_/B1 _10644_/X _06743_/B vssd1 vssd1 vccd1 vccd1 _10645_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__07896__B _09396_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13364_ _13365_/CLK _13364_/D vssd1 vssd1 vccd1 vccd1 hold277/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09169__A _09170_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12315_ _12316_/B _12315_/B vssd1 vssd1 vccd1 vccd1 _12319_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_2_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10576_ _11180_/A _10576_/B _10576_/C vssd1 vssd1 vccd1 vccd1 _10579_/C sky130_fd_sc_hd__and3_1
X_13295_ _13299_/CLK hold191/X vssd1 vssd1 vccd1 vccd1 _13295_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12246_ _09355_/X _12301_/B hold256/A vssd1 vssd1 vccd1 vccd1 _12246_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_121_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10899__B1 _10896_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12177_ _12176_/A _12175_/B _12175_/Y _11624_/A vssd1 vssd1 vccd1 vccd1 _12177_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_48_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09753__A1 _10941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09753__B2 fanout94/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11128_ _11450_/B _11236_/B hold228/A vssd1 vssd1 vccd1 vccd1 _11128_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__09108__S _09108_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06959__C _09666_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11059_ _11059_/A _11059_/B vssd1 vssd1 vccd1 vccd1 _11061_/B sky130_fd_sc_hd__xor2_1
XANTENNA__13065__A1 _07090_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09351__B _09351_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07295__A2 _11751_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08270_ _08330_/A _08330_/B _08280_/B vssd1 vssd1 vccd1 vccd1 _08270_/X sky130_fd_sc_hd__or3_1
XFILLER_0_27_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07221_ _08038_/B _08038_/C vssd1 vssd1 vccd1 vccd1 _07221_/X sky130_fd_sc_hd__or2_1
XFILLER_0_61_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07152_ _07144_/A _07343_/B _07141_/X _07223_/B _06838_/B vssd1 vssd1 vccd1 vccd1
+ _07154_/A sky130_fd_sc_hd__a311o_4
XFILLER_0_82_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11379__B2 _07819_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11379__A1 fanout24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10051__A1 _10570_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11121__B _11121_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09992__A1 _12429_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07083_ reg1_val[19] _07083_/B vssd1 vssd1 vccd1 vccd1 _07833_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_30_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10051__B2 _10571_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09807__A _09808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09744__A1 _07099_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout104 _07028_/X vssd1 vssd1 vccd1 vccd1 _11758_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_0_10_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12233__A _12341_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout115 _08304_/B vssd1 vssd1 vccd1 vccd1 _10948_/B2 sky130_fd_sc_hd__buf_6
Xfanout137 _12812_/A vssd1 vssd1 vccd1 vccd1 _10413_/A sky130_fd_sc_hd__buf_6
Xfanout126 _06955_/X vssd1 vssd1 vccd1 vccd1 _10537_/A1 sky130_fd_sc_hd__buf_8
XFILLER_0_1_195 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout159 _12170_/A vssd1 vssd1 vccd1 vccd1 _11874_/A sky130_fd_sc_hd__buf_4
X_07985_ _07986_/A _07986_/B _07986_/C vssd1 vssd1 vccd1 vccd1 _08925_/A sky130_fd_sc_hd__o21ai_1
Xfanout148 _07026_/X vssd1 vssd1 vccd1 vccd1 _12804_/A sky130_fd_sc_hd__buf_8
X_06936_ instruction[6] instruction[5] vssd1 vssd1 vccd1 vccd1 _09159_/B sky130_fd_sc_hd__nand2b_2
X_09724_ _09724_/A _09724_/B vssd1 vssd1 vccd1 vccd1 _09726_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__07046__B _11180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06867_ _10507_/A _06867_/B vssd1 vssd1 vccd1 vccd1 _06869_/C sky130_fd_sc_hd__nand2_1
X_09655_ _11707_/A _09655_/B _09655_/C vssd1 vssd1 vccd1 vccd1 _09699_/A sky130_fd_sc_hd__and3_1
X_08606_ _08606_/A _08615_/A vssd1 vssd1 vccd1 vccd1 _08607_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08180__B1 _08656_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06798_ _09684_/B _06798_/B vssd1 vssd1 vccd1 vccd1 _09527_/A sky130_fd_sc_hd__nand2b_2
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09586_ _09906_/A _09586_/B vssd1 vssd1 vccd1 vccd1 _09588_/B sky130_fd_sc_hd__xnor2_1
X_08537_ _08573_/A _08573_/B vssd1 vssd1 vccd1 vccd1 _08574_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_65_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08468_ _08495_/A _08495_/B _08464_/X vssd1 vssd1 vccd1 vccd1 _08483_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_92_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07419_ _07420_/A _07420_/B vssd1 vssd1 vccd1 vccd1 _12412_/A sky130_fd_sc_hd__nor2_4
XFILLER_0_80_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08399_ _08447_/A _08398_/B _08394_/X vssd1 vssd1 vccd1 vccd1 _08405_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_45_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10430_ _10430_/A _10430_/B vssd1 vssd1 vccd1 vccd1 _10441_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_18_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09432__B1 _09568_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07038__A2 _10574_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_1_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10361_ _10361_/A _10361_/B vssd1 vssd1 vccd1 vccd1 _10364_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_20_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13080_ hold113/X _12791_/A _13080_/B1 hold72/X _13113_/A vssd1 vssd1 vccd1 vccd1
+ hold129/A sky130_fd_sc_hd__o221a_1
X_12100_ _11427_/B _11787_/Y _12099_/B _12099_/X _12097_/X vssd1 vssd1 vccd1 vccd1
+ _12101_/B sky130_fd_sc_hd__a311oi_4
X_10292_ _10292_/A _10292_/B _10292_/C vssd1 vssd1 vccd1 vccd1 _10293_/B sky130_fd_sc_hd__or3_1
Xhold180 hold223/X vssd1 vssd1 vccd1 vccd1 hold180/X sky130_fd_sc_hd__dlygate4sd3_1
X_12031_ _12031_/A _12031_/B _12031_/C vssd1 vssd1 vccd1 vccd1 _12031_/X sky130_fd_sc_hd__or3_1
Xhold191 hold191/A vssd1 vssd1 vccd1 vccd1 hold191/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11542__A1 _07131_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12933_ _13164_/B _13165_/A _12883_/X vssd1 vssd1 vccd1 vccd1 _13170_/A sky130_fd_sc_hd__a21o_1
XANTENNA__10502__C1 _11707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12864_ hold39/X hold281/A vssd1 vssd1 vccd1 vccd1 _12864_/X sky130_fd_sc_hd__and2b_1
XANTENNA__13047__A1 _10444_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11815_ _11806_/Y _11807_/X _11810_/X _11814_/Y vssd1 vssd1 vccd1 vccd1 _11815_/X
+ sky130_fd_sc_hd__o211a_1
X_12795_ hold59/X _12798_/B _12794_/Y _13109_/A vssd1 vssd1 vccd1 vccd1 hold60/A sky130_fd_sc_hd__o211a_1
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10805__B1 _10930_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11746_ _11746_/A _11746_/B vssd1 vssd1 vccd1 vccd1 _11750_/A sky130_fd_sc_hd__and2_1
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10281__B2 fanout66/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10281__A1 _07087_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11677_ _11677_/A _11677_/B vssd1 vssd1 vccd1 vccd1 _11691_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_113_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10628_ _06817_/Y _10627_/Y _12174_/S vssd1 vssd1 vccd1 vccd1 _10629_/B sky130_fd_sc_hd__mux2_1
XANTENNA__09423__B1 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13347_ _13380_/CLK _13347_/D vssd1 vssd1 vccd1 vccd1 hold260/A sky130_fd_sc_hd__dfxtp_2
XFILLER_0_106_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10559_ _12076_/A _10559_/B vssd1 vssd1 vccd1 vccd1 _10560_/B sky130_fd_sc_hd__xnor2_1
X_13278_ _13378_/CLK hold40/X vssd1 vssd1 vccd1 vccd1 hold39/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12229_ _11949_/B _12228_/Y _12227_/Y vssd1 vssd1 vccd1 vccd1 _12230_/B sky130_fd_sc_hd__o21a_1
XANTENNA__07147__A _09594_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07770_ _07770_/A _07770_/B vssd1 vssd1 vccd1 vccd1 _07781_/A sky130_fd_sc_hd__xnor2_1
X_06721_ _06805_/A _06702_/A _12698_/B _06720_/X vssd1 vssd1 vccd1 vccd1 _11020_/A
+ sky130_fd_sc_hd__a31o_4
XANTENNA__06986__A _10707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09440_ _12852_/A _09238_/B _09440_/B1 _12854_/A vssd1 vssd1 vccd1 vccd1 _09441_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11836__A2 _07037_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06652_ reg2_val[23] _06720_/B _06703_/B1 _06651_/Y vssd1 vssd1 vccd1 vccd1 _07194_/A
+ sky130_fd_sc_hd__o2bb2a_2
XANTENNA__09081__B _09170_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06583_ instruction[0] instruction[2] instruction[1] pred_val vssd1 vssd1 vccd1 vccd1
+ _06596_/A sky130_fd_sc_hd__and4bb_4
X_09371_ _09371_/A _09371_/B _09371_/C vssd1 vssd1 vccd1 vccd1 _09372_/B sky130_fd_sc_hd__and3_1
XFILLER_0_47_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08465__A1 _12802_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08322_ _08322_/A _08322_/B vssd1 vssd1 vccd1 vccd1 _08373_/A sky130_fd_sc_hd__xor2_1
XANTENNA__08465__B2 _07896_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08253_ _08253_/A _08253_/B vssd1 vssd1 vccd1 vccd1 _08293_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_117_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07204_ _07208_/A _07208_/B _10444_/A vssd1 vssd1 vccd1 vccd1 _07204_/X sky130_fd_sc_hd__mux2_4
XFILLER_0_74_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08184_ _08187_/A _08187_/B vssd1 vssd1 vccd1 vccd1 _08189_/A sky130_fd_sc_hd__or2_1
XFILLER_0_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07135_ _07194_/A _07135_/B _07223_/A _07135_/D vssd1 vssd1 vccd1 vccd1 _07142_/C
+ sky130_fd_sc_hd__and4_2
XFILLER_0_42_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07066_ _07100_/B _07066_/B _06963_/A vssd1 vssd1 vccd1 vccd1 _07067_/B sky130_fd_sc_hd__or3b_2
XFILLER_0_113_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08441__A _09445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07440__A2 fanout16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07968_ _07968_/A _07968_/B vssd1 vssd1 vccd1 vccd1 _07969_/C sky130_fd_sc_hd__xnor2_1
X_06919_ instruction[28] _06921_/B vssd1 vssd1 vccd1 vccd1 _06919_/X sky130_fd_sc_hd__or2_1
X_09707_ _08977_/A _08977_/B _09706_/X vssd1 vssd1 vccd1 vccd1 _09810_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_4_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07899_ _07821_/A _07087_/A _07087_/B _08752_/B _07752_/B vssd1 vssd1 vccd1 vccd1
+ _07900_/B sky130_fd_sc_hd__o32a_1
XANTENNA__08153__B1 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09638_ _09474_/A _09474_/B _09472_/Y vssd1 vssd1 vccd1 vccd1 _09639_/B sky130_fd_sc_hd__a21boi_4
XFILLER_0_69_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout45_A _12840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09569_ _09570_/B _09570_/C _10165_/A vssd1 vssd1 vccd1 vccd1 _09573_/A sky130_fd_sc_hd__a21o_1
X_12580_ _12580_/A _12580_/B vssd1 vssd1 vccd1 vccd1 _12595_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_77_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11600_ _11601_/B _11601_/A vssd1 vssd1 vccd1 vccd1 _11697_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_108_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11531_ _11442_/A _11439_/Y _11441_/B vssd1 vssd1 vccd1 vccd1 _11532_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_93_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12252__A2 _11343_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12138__A _12138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11460__B1 _12067_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11042__A _11470_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11462_ _11653_/A _12316_/A fanout12/X _08752_/B vssd1 vssd1 vccd1 vccd1 _11463_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_18_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13201_ _13214_/A _13201_/B vssd1 vssd1 vccd1 vccd1 _13370_/D sky130_fd_sc_hd__and2_1
X_11393_ _11391_/Y _11393_/B vssd1 vssd1 vccd1 vccd1 _11394_/B sky130_fd_sc_hd__and2b_1
X_10413_ _10413_/A _12316_/B _10413_/C _10413_/D vssd1 vssd1 vccd1 vccd1 _10415_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_0_21_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12960__B1 fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13132_ hold288/X _12789_/B _13131_/X _12790_/A vssd1 vssd1 vccd1 vccd1 hold289/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10344_ _10344_/A _10344_/B vssd1 vssd1 vccd1 vccd1 _10345_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_104_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08351__A _08742_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07012__A_N _12076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13063_ _07833_/A _13087_/B2 hold100/X vssd1 vssd1 vccd1 vccd1 _13334_/D sky130_fd_sc_hd__o21a_1
X_10275_ _10275_/A _10275_/B _10275_/C _10275_/D vssd1 vssd1 vccd1 vccd1 _11033_/A
+ sky130_fd_sc_hd__nand4_2
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10318__A2 _10589_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09184__A2 _09152_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07195__A1 _09567_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12014_ _12089_/B _12013_/C _12013_/A vssd1 vssd1 vccd1 vccd1 _12014_/X sky130_fd_sc_hd__a21o_1
XANTENNA__08392__B1 _08645_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07195__B2 _12840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12916_ hold260/A hold132/X vssd1 vssd1 vccd1 vccd1 _13092_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_76_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12847_ hold29/X _12848_/B _12846_/Y _13210_/A vssd1 vssd1 vccd1 vccd1 hold30/A sky130_fd_sc_hd__o211a_1
XFILLER_0_29_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12778_ _12772_/B _12774_/B _12772_/A vssd1 vssd1 vccd1 vccd1 _12779_/B sky130_fd_sc_hd__a21bo_2
XFILLER_0_28_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11729_ _07223_/A _11343_/B _11728_/X _06669_/B vssd1 vssd1 vccd1 vccd1 _11729_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_126_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10791__A _11269_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07958__B1 _08752_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08940_ _08937_/A _08937_/B _08935_/X vssd1 vssd1 vccd1 vccd1 _08954_/A sky130_fd_sc_hd__a21o_2
X_08871_ _08859_/A _08859_/B _08860_/X vssd1 vssd1 vccd1 vccd1 _08882_/A sky130_fd_sc_hd__a21o_1
X_07822_ _11908_/A _07822_/B _07822_/C vssd1 vssd1 vccd1 vccd1 _07824_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_19_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07753_ _11908_/A _07753_/B _07753_/C vssd1 vssd1 vccd1 vccd1 _07753_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_126_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06704_ reg1_val[16] _11343_/A vssd1 vssd1 vccd1 vccd1 _06704_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__08686__A1 _09445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07684_ _07685_/A _07685_/B vssd1 vssd1 vccd1 vccd1 _09304_/A sky130_fd_sc_hd__and2_1
XANTENNA__10031__A _12138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06635_ _06635_/A _12680_/B vssd1 vssd1 vccd1 vccd1 _06635_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_79_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09423_ _12802_/A fanout9/A fanout5/X _09423_/B2 vssd1 vssd1 vccd1 vccd1 _09424_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_66_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09354_ _09663_/S _09354_/B _09343_/A vssd1 vssd1 vccd1 vccd1 _09354_/X sky130_fd_sc_hd__or3b_1
XFILLER_0_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06566_ hold295/X vssd1 vssd1 vccd1 vccd1 _06566_/Y sky130_fd_sc_hd__inv_2
XANTENNA__07340__A _09594_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08436__A _08436_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08305_ _08724_/A _08305_/B vssd1 vssd1 vccd1 vccd1 _08370_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09285_ _09285_/A _09285_/B vssd1 vssd1 vccd1 vccd1 _09298_/A sky130_fd_sc_hd__xor2_4
XANTENNA__07110__B2 _12808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07110__A1 _10574_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07661__A2 _10167_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08236_ _08287_/A _08287_/B _08232_/X vssd1 vssd1 vccd1 vccd1 _08282_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_28_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08167_ _08167_/A _08167_/B vssd1 vssd1 vccd1 vccd1 _08253_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_15_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07118_ _12626_/A _09343_/A reg1_val[2] _07200_/A vssd1 vssd1 vccd1 vccd1 _07120_/B
+ sky130_fd_sc_hd__o31a_2
X_08098_ _08098_/A _08098_/B vssd1 vssd1 vccd1 vccd1 _08110_/A sky130_fd_sc_hd__xor2_2
XANTENNA__08171__A _11385_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07049_ _07074_/B _06964_/A _09147_/S vssd1 vssd1 vccd1 vccd1 _08632_/A sky130_fd_sc_hd__a21o_2
XFILLER_0_30_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09166__A2 _11973_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10060_ _10061_/A _10061_/B vssd1 vssd1 vccd1 vccd1 _10062_/A sky130_fd_sc_hd__and2_1
XANTENNA__07177__A1 _07074_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10181__B1 fanout59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10962_ _10962_/A _10962_/B vssd1 vssd1 vccd1 vccd1 _10964_/A sky130_fd_sc_hd__nand2_1
X_12701_ _12701_/A _12701_/B _12701_/C vssd1 vssd1 vccd1 vccd1 _12702_/B sky130_fd_sc_hd__nand3_1
X_10893_ hold285/A _10893_/B vssd1 vssd1 vccd1 vccd1 _11017_/B sky130_fd_sc_hd__or2_1
XFILLER_0_66_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12632_ _12631_/A _12631_/B _12630_/A vssd1 vssd1 vccd1 vccd1 _12636_/A sky130_fd_sc_hd__o21a_2
X_12563_ _12623_/A _12564_/B vssd1 vssd1 vccd1 vccd1 _12582_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_93_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12494_ _12495_/A _12495_/B _12495_/C vssd1 vssd1 vccd1 vccd1 _12502_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_81_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11514_ _11514_/A _11702_/A vssd1 vssd1 vccd1 vccd1 _11515_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_25_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11445_ _06698_/X _09527_/B _12307_/B1 vssd1 vssd1 vccd1 vccd1 _11445_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_80_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10539__A2 _12214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09177__A _11118_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07404__A2 _12830_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11376_ _11377_/A _11377_/B vssd1 vssd1 vccd1 vccd1 _11378_/A sky130_fd_sc_hd__and2_1
X_13115_ _13115_/A _13115_/B vssd1 vssd1 vccd1 vccd1 _13115_/Y sky130_fd_sc_hd__xnor2_1
X_10327_ _10328_/A _10328_/B vssd1 vssd1 vccd1 vccd1 _10474_/B sky130_fd_sc_hd__nand2b_1
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10258_ hold294/A _09835_/B _10522_/C _09837_/A vssd1 vssd1 vccd1 vccd1 _10258_/X
+ sky130_fd_sc_hd__a31o_1
X_13046_ hold150/A _12788_/A _13236_/B hold134/X _13109_/A vssd1 vssd1 vccd1 vccd1
+ hold135/A sky130_fd_sc_hd__o221a_1
XFILLER_0_56_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10189_ _11163_/A _10189_/B vssd1 vssd1 vccd1 vccd1 _10190_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__09116__S _09142_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09865__B1 _10963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06983__B _10949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11672__B1 _12067_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07891__A2 _08721_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07160__A _07200_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11975__A1 _07194_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09070_ _09077_/A _09077_/B _12392_/A vssd1 vssd1 vccd1 vccd1 _12426_/B sky130_fd_sc_hd__and3_1
XFILLER_0_71_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08021_ _08021_/A _08021_/B vssd1 vssd1 vccd1 vccd1 _08022_/B sky130_fd_sc_hd__xor2_2
XANTENNA__07643__A2 fanout24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12506__A _12669_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout6 fanout8/X vssd1 vssd1 vccd1 vccd1 fanout6/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_40_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09972_ _11231_/S _09972_/B vssd1 vssd1 vccd1 vccd1 _09972_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_97_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08923_ _08923_/A _08923_/B vssd1 vssd1 vccd1 vccd1 _08936_/A sky130_fd_sc_hd__and2_2
XANTENNA_fanout297_A _13242_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08356__B1 _09440_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08854_ _08813_/A _08813_/C _08813_/B vssd1 vssd1 vccd1 vccd1 _08857_/B sky130_fd_sc_hd__a21boi_2
XANTENNA__10163__B1 _10710_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08785_ _08787_/B _08786_/B vssd1 vssd1 vccd1 vccd1 _08788_/A sky130_fd_sc_hd__and2b_1
X_07805_ _07805_/A _07805_/B _07805_/C vssd1 vssd1 vccd1 vccd1 _07806_/C sky130_fd_sc_hd__nand3_1
X_07736_ _10537_/A1 _12818_/A _12820_/A _08432_/B vssd1 vssd1 vccd1 vccd1 _07737_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11112__C1 _09156_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09550__A _09716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10466__A1 _10941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07667_ _08916_/B _08916_/A vssd1 vssd1 vccd1 vccd1 _07667_/X sky130_fd_sc_hd__and2b_1
XANTENNA__10466__B2 fanout94/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06618_ reg1_val[29] _06838_/B vssd1 vssd1 vccd1 vccd1 _06621_/B sky130_fd_sc_hd__or2_1
X_07598_ _07598_/A _07598_/B vssd1 vssd1 vccd1 vccd1 _07685_/A sky130_fd_sc_hd__xnor2_4
X_09406_ _11065_/A _07090_/Y _10963_/A _11653_/A vssd1 vssd1 vccd1 vccd1 _09407_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07882__A2 fanout99/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09337_ _09335_/X _09336_/X _09663_/S vssd1 vssd1 vccd1 vccd1 _09974_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_75_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09268_ _10574_/A _10567_/A vssd1 vssd1 vccd1 vccd1 _09270_/B sky130_fd_sc_hd__or2_1
XFILLER_0_35_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08219_ _08733_/A _08219_/B vssd1 vssd1 vccd1 vccd1 _08225_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09199_ _09199_/A _09199_/B vssd1 vssd1 vccd1 vccd1 _09200_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_62_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11230_ _11230_/A _11230_/B vssd1 vssd1 vccd1 vccd1 _11230_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__09387__A2 _12808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08595__B1 _08038_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11161_ _09609_/B fanout56/X _12316_/A _09396_/B vssd1 vssd1 vccd1 vccd1 _11162_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10112_ _10119_/S _10111_/X _09181_/X vssd1 vssd1 vccd1 vccd1 _10113_/B sky130_fd_sc_hd__o21ai_2
X_11092_ _11092_/A _11092_/B vssd1 vssd1 vccd1 vccd1 _11095_/A sky130_fd_sc_hd__xor2_1
Xhold40 hold40/A vssd1 vssd1 vccd1 vccd1 hold40/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09444__B fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10043_ _10042_/B _10042_/C _10042_/A vssd1 vssd1 vccd1 vccd1 _10044_/B sky130_fd_sc_hd__o21ai_1
Xhold62 hold62/A vssd1 vssd1 vccd1 vccd1 hold62/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 hold73/A vssd1 vssd1 vccd1 vccd1 hold73/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 hold51/A vssd1 vssd1 vccd1 vccd1 hold51/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07245__A _10165_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold95 hold95/A vssd1 vssd1 vccd1 vccd1 hold95/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 hold84/A vssd1 vssd1 vccd1 vccd1 hold84/X sky130_fd_sc_hd__dlygate4sd3_1
X_11994_ _11929_/A _11928_/B _11926_/Y vssd1 vssd1 vccd1 vccd1 _12009_/A sky130_fd_sc_hd__a21o_1
XANTENNA__12851__C1 _13128_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10945_ _10947_/B _10947_/C _10448_/A vssd1 vssd1 vccd1 vccd1 _11076_/C sky130_fd_sc_hd__a21boi_1
XFILLER_0_128_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10876_ _10752_/A _10750_/X _10767_/S vssd1 vssd1 vccd1 vccd1 _10876_/X sky130_fd_sc_hd__a21o_1
XANTENNA__07873__A2 _11751_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12615_ reg1_val[26] curr_PC[26] _12622_/S vssd1 vssd1 vccd1 vccd1 _12617_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_54_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11957__A1 _12174_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07086__B1 _11261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12546_ reg1_val[15] curr_PC[15] _12586_/S vssd1 vssd1 vccd1 vccd1 _12548_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_53_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_666 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12477_ _12649_/B _12478_/B vssd1 vssd1 vccd1 vccd1 _12488_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_81_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11428_ _11649_/B vssd1 vssd1 vccd1 vccd1 _11428_/Y sky130_fd_sc_hd__inv_2
XANTENNA_4 instruction[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11359_ _11550_/B _11358_/Y _11142_/S vssd1 vssd1 vccd1 vccd1 _11359_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13029_ _07127_/B _12798_/B hold105/X vssd1 vssd1 vccd1 vccd1 hold106/A sky130_fd_sc_hd__a21boi_1
XANTENNA__09354__B _09354_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08570_ _08570_/A _08570_/B vssd1 vssd1 vccd1 vccd1 _08571_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__09838__B1 _09354_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12437__A2 _07064_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07521_ _07688_/B _12804_/A _12802_/A fanout30/X vssd1 vssd1 vccd1 vccd1 _07522_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_13_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07452_ _07360_/A _07360_/B _07357_/A vssd1 vssd1 vccd1 vccd1 _07561_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_9_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07383_ _10422_/A _07383_/B vssd1 vssd1 vccd1 vccd1 _07385_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_57_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09122_ _09118_/X _09121_/X _09663_/S vssd1 vssd1 vccd1 vccd1 _09122_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_72_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07077__B1 _10818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12070__B1 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10963__B _12316_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout212_A _09445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09053_ _09053_/A _09056_/B vssd1 vssd1 vccd1 vccd1 _09059_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_44_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08004_ _08004_/A _08004_/B vssd1 vssd1 vccd1 vccd1 _08006_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_40_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_6_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09955_ _09956_/B _09956_/C _10496_/A vssd1 vssd1 vccd1 vccd1 _09957_/A sky130_fd_sc_hd__a21o_1
XANTENNA__09264__B _10570_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09886_ _09743_/A _09743_/B _09742_/A vssd1 vssd1 vccd1 vccd1 _09890_/B sky130_fd_sc_hd__o21ai_1
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08906_ _08867_/X _08884_/Y _08883_/X vssd1 vssd1 vccd1 vccd1 _08906_/Y sky130_fd_sc_hd__a21oi_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08837_ _08838_/A _08838_/B vssd1 vssd1 vccd1 vccd1 _09043_/B sky130_fd_sc_hd__nor2_1
XANTENNA__09829__B1 _09152_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08768_ _08111_/A _08111_/B _08121_/B _08139_/A _08139_/B vssd1 vssd1 vccd1 vccd1
+ _08779_/A sky130_fd_sc_hd__a32o_1
X_08699_ _08699_/A _08699_/B vssd1 vssd1 vccd1 vccd1 _09002_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_67_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07719_ _07719_/A _07719_/B vssd1 vssd1 vccd1 vccd1 _07746_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__09844__A3 _09843_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10730_ _10731_/A _10731_/B vssd1 vssd1 vccd1 vccd1 _10858_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_94_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10661_ _10606_/A _10606_/B _10607_/Y vssd1 vssd1 vccd1 vccd1 _10733_/A sky130_fd_sc_hd__o21ai_4
X_12400_ _08979_/X _12399_/X hold215/A vssd1 vssd1 vccd1 vccd1 _12400_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_75_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13380_ _13380_/CLK hold64/X vssd1 vssd1 vccd1 vccd1 hold297/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_105_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07607__A2 _07087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10592_ _10592_/A _10700_/A vssd1 vssd1 vccd1 vccd1 _10594_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_105_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12331_ _12414_/A _12414_/B vssd1 vssd1 vccd1 vccd1 _12334_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_121_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12262_ _12263_/A _12263_/B vssd1 vssd1 vccd1 vccd1 _12325_/A sky130_fd_sc_hd__nand2_1
XANTENNA__12364__A1 _12317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11213_ _11100_/B _11318_/A vssd1 vssd1 vccd1 vccd1 _11423_/A sky130_fd_sc_hd__nand2b_1
X_12193_ hold223/A _12434_/B1 _12248_/B _12401_/B1 vssd1 vssd1 vccd1 vccd1 _12194_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_120_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10375__B1 _09163_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09455__A _09906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11144_ _11090_/A _11090_/B _11089_/A vssd1 vssd1 vccd1 vccd1 _11207_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_128_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10127__B1 _11973_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07791__B2 _11472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11075_ _11076_/A _11076_/B _11076_/C _11076_/D vssd1 vssd1 vccd1 vccd1 _11075_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07791__A1 _11367_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10678__A1 _10570_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10678__B2 _10571_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10026_ _10027_/A _10027_/B vssd1 vssd1 vccd1 vccd1 _10147_/A sky130_fd_sc_hd__and2_1
X_11977_ _11971_/Y _11972_/X _11976_/X _11969_/X vssd1 vssd1 vccd1 vccd1 _11977_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_85_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08099__A2 _08727_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10928_ _10928_/A _10928_/B vssd1 vssd1 vccd1 vccd1 _10935_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__06740__A_N _07100_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10859_ _10859_/A _10859_/B vssd1 vssd1 vccd1 vccd1 _11100_/A sky130_fd_sc_hd__xor2_4
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08534__A _08742_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12529_ _12530_/A _12530_/B _12530_/C vssd1 vssd1 vccd1 vccd1 _12537_/B sky130_fd_sc_hd__a21o_1
XANTENNA__08271__A2 fanout87/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout308 reg1_val[0] vssd1 vssd1 vccd1 vccd1 _12626_/A sky130_fd_sc_hd__buf_8
XFILLER_0_1_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09740_ _09741_/A _09741_/B vssd1 vssd1 vccd1 vccd1 _09742_/A sky130_fd_sc_hd__or2_1
X_06952_ _10710_/A _06954_/B vssd1 vssd1 vccd1 vccd1 _06952_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_10_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
.ends

