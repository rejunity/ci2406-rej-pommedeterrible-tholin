VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO vliw
  CLASS BLOCK ;
  FOREIGN vliw ;
  ORIGIN 0.000 0.000 ;
  SIZE 2100.000 BY 640.000 ;
  PIN curr_PC[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.251000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 29.070 636.000 29.350 640.000 ;
    END
  END curr_PC[0]
  PIN curr_PC[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.877500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 107.270 636.000 107.550 640.000 ;
    END
  END curr_PC[10]
  PIN curr_PC[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.751500 ;
    ANTENNADIFFAREA 1.325700 ;
    PORT
      LAYER met2 ;
        RECT 115.090 636.000 115.370 640.000 ;
    END
  END curr_PC[11]
  PIN curr_PC[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.867500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 122.910 636.000 123.190 640.000 ;
    END
  END curr_PC[12]
  PIN curr_PC[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.372500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 130.730 636.000 131.010 640.000 ;
    END
  END curr_PC[13]
  PIN curr_PC[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.877500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 138.550 636.000 138.830 640.000 ;
    END
  END curr_PC[14]
  PIN curr_PC[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.630000 ;
    ANTENNADIFFAREA 1.760400 ;
    PORT
      LAYER met2 ;
        RECT 146.370 636.000 146.650 640.000 ;
    END
  END curr_PC[15]
  PIN curr_PC[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.246500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 154.190 636.000 154.470 640.000 ;
    END
  END curr_PC[16]
  PIN curr_PC[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.751500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 162.010 636.000 162.290 640.000 ;
    END
  END curr_PC[17]
  PIN curr_PC[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.877500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 169.830 636.000 170.110 640.000 ;
    END
  END curr_PC[18]
  PIN curr_PC[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.630000 ;
    ANTENNADIFFAREA 1.760400 ;
    PORT
      LAYER met2 ;
        RECT 177.650 636.000 177.930 640.000 ;
    END
  END curr_PC[19]
  PIN curr_PC[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.251000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 36.890 636.000 37.170 640.000 ;
    END
  END curr_PC[1]
  PIN curr_PC[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.877500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 185.470 636.000 185.750 640.000 ;
    END
  END curr_PC[20]
  PIN curr_PC[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.751500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 193.290 636.000 193.570 640.000 ;
    END
  END curr_PC[21]
  PIN curr_PC[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.877500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 201.110 636.000 201.390 640.000 ;
    END
  END curr_PC[22]
  PIN curr_PC[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.246500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 208.930 636.000 209.210 640.000 ;
    END
  END curr_PC[23]
  PIN curr_PC[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.751500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 216.750 636.000 217.030 640.000 ;
    END
  END curr_PC[24]
  PIN curr_PC[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.751500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 224.570 636.000 224.850 640.000 ;
    END
  END curr_PC[25]
  PIN curr_PC[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.069500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 232.390 636.000 232.670 640.000 ;
    END
  END curr_PC[26]
  PIN curr_PC[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.751500 ;
    ANTENNADIFFAREA 1.760400 ;
    PORT
      LAYER met2 ;
        RECT 240.210 636.000 240.490 640.000 ;
    END
  END curr_PC[27]
  PIN curr_PC[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.784500 ;
    ANTENNADIFFAREA 1.760400 ;
    PORT
      LAYER met2 ;
        RECT 44.710 636.000 44.990 640.000 ;
    END
  END curr_PC[2]
  PIN curr_PC[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.537000 ;
    ANTENNADIFFAREA 1.325700 ;
    PORT
      LAYER met2 ;
        RECT 52.530 636.000 52.810 640.000 ;
    END
  END curr_PC[3]
  PIN curr_PC[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.251000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 60.350 636.000 60.630 640.000 ;
    END
  END curr_PC[4]
  PIN curr_PC[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.838500 ;
    ANTENNADIFFAREA 1.760400 ;
    PORT
      LAYER met2 ;
        RECT 68.170 636.000 68.450 640.000 ;
    END
  END curr_PC[5]
  PIN curr_PC[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.658500 ;
    ANTENNADIFFAREA 1.325700 ;
    PORT
      LAYER met2 ;
        RECT 75.990 636.000 76.270 640.000 ;
    END
  END curr_PC[6]
  PIN curr_PC[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.494000 ;
    ANTENNADIFFAREA 1.760400 ;
    PORT
      LAYER met2 ;
        RECT 83.810 636.000 84.090 640.000 ;
    END
  END curr_PC[7]
  PIN curr_PC[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.877500 ;
    ANTENNADIFFAREA 1.325700 ;
    PORT
      LAYER met2 ;
        RECT 91.630 636.000 91.910 640.000 ;
    END
  END curr_PC[8]
  PIN curr_PC[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.372500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 99.450 636.000 99.730 640.000 ;
    END
  END curr_PC[9]
  PIN custom_settings[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 2000.630 0.000 2000.910 4.000 ;
    END
  END custom_settings[0]
  PIN custom_settings[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 2018.570 0.000 2018.850 4.000 ;
    END
  END custom_settings[1]
  PIN custom_settings[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.719500 ;
    PORT
      LAYER met2 ;
        RECT 2036.510 0.000 2036.790 4.000 ;
    END
  END custom_settings[2]
  PIN custom_settings[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.719500 ;
    PORT
      LAYER met2 ;
        RECT 2054.450 0.000 2054.730 4.000 ;
    END
  END custom_settings[3]
  PIN custom_settings[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2072.390 0.000 2072.670 4.000 ;
    END
  END custom_settings[4]
  PIN dest_idx0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.348000 ;
    PORT
      LAYER met2 ;
        RECT 592.110 636.000 592.390 640.000 ;
    END
  END dest_idx0[0]
  PIN dest_idx0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.348000 ;
    PORT
      LAYER met2 ;
        RECT 599.930 636.000 600.210 640.000 ;
    END
  END dest_idx0[1]
  PIN dest_idx0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.494000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 607.750 636.000 608.030 640.000 ;
    END
  END dest_idx0[2]
  PIN dest_idx0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.494000 ;
    PORT
      LAYER met2 ;
        RECT 615.570 636.000 615.850 640.000 ;
    END
  END dest_idx0[3]
  PIN dest_idx0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.494000 ;
    PORT
      LAYER met2 ;
        RECT 623.390 636.000 623.670 640.000 ;
    END
  END dest_idx0[4]
  PIN dest_idx1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.348000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 121.080 2100.000 121.680 ;
    END
  END dest_idx1[0]
  PIN dest_idx1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.348000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 123.800 2100.000 124.400 ;
    END
  END dest_idx1[1]
  PIN dest_idx1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 126.520 2100.000 127.120 ;
    END
  END dest_idx1[2]
  PIN dest_idx1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 129.240 2100.000 129.840 ;
    END
  END dest_idx1[3]
  PIN dest_idx1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.494000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 131.960 2100.000 132.560 ;
    END
  END dest_idx1[4]
  PIN dest_idx2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.618000 ;
    ANTENNADIFFAREA 6.955200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.080 4.000 121.680 ;
    END
  END dest_idx2[0]
  PIN dest_idx2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.618000 ;
    ANTENNADIFFAREA 16.953300 ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.800 4.000 124.400 ;
    END
  END dest_idx2[1]
  PIN dest_idx2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.780000 ;
    ANTENNADIFFAREA 6.085800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.520 4.000 127.120 ;
    END
  END dest_idx2[2]
  PIN dest_idx2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.780000 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END dest_idx2[3]
  PIN dest_idx2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.780000 ;
    ANTENNADIFFAREA 16.953300 ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.960 4.000 132.560 ;
    END
  END dest_idx2[4]
  PIN dest_mask0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.363500 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met2 ;
        RECT 576.470 636.000 576.750 640.000 ;
    END
  END dest_mask0[0]
  PIN dest_mask0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.621000 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met2 ;
        RECT 584.290 636.000 584.570 640.000 ;
    END
  END dest_mask0[1]
  PIN dest_mask1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.732500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 115.640 2100.000 116.240 ;
    END
  END dest_mask1[0]
  PIN dest_mask1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.732500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 118.360 2100.000 118.960 ;
    END
  END dest_mask1[1]
  PIN dest_mask2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.485000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END dest_mask2[0]
  PIN dest_mask2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.980000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.360 4.000 118.960 ;
    END
  END dest_mask2[1]
  PIN dest_pred0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.751500 ;
    ANTENNADIFFAREA 2.173500 ;
    PORT
      LAYER met2 ;
        RECT 654.670 636.000 654.950 640.000 ;
    END
  END dest_pred0[0]
  PIN dest_pred0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.882000 ;
    PORT
      LAYER met2 ;
        RECT 662.490 636.000 662.770 640.000 ;
    END
  END dest_pred0[1]
  PIN dest_pred0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.882000 ;
    ANTENNADIFFAREA 3.042900 ;
    PORT
      LAYER met2 ;
        RECT 670.310 636.000 670.590 640.000 ;
    END
  END dest_pred0[2]
  PIN dest_pred1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.868500 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 142.840 2100.000 143.440 ;
    END
  END dest_pred1[0]
  PIN dest_pred1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.251000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 145.560 2100.000 146.160 ;
    END
  END dest_pred1[1]
  PIN dest_pred1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.251000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 148.280 2100.000 148.880 ;
    END
  END dest_pred1[2]
  PIN dest_pred2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.994500 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END dest_pred2[0]
  PIN dest_pred2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.877500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.560 4.000 146.160 ;
    END
  END dest_pred2[1]
  PIN dest_pred2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.877500 ;
    ANTENNADIFFAREA 2.173500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.280 4.000 148.880 ;
    END
  END dest_pred2[2]
  PIN dest_pred_val0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.882000 ;
    PORT
      LAYER met2 ;
        RECT 678.130 636.000 678.410 640.000 ;
    END
  END dest_pred_val0
  PIN dest_pred_val1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.120500 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 151.000 2100.000 151.600 ;
    END
  END dest_pred_val1
  PIN dest_pred_val2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.003500 ;
    ANTENNADIFFAREA 3.042900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.000 4.000 151.600 ;
    END
  END dest_pred_val2
  PIN dest_val0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.673500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 326.230 636.000 326.510 640.000 ;
    END
  END dest_val0[0]
  PIN dest_val0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 404.430 636.000 404.710 640.000 ;
    END
  END dest_val0[10]
  PIN dest_val0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.673500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 412.250 636.000 412.530 640.000 ;
    END
  END dest_val0[11]
  PIN dest_val0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 420.070 636.000 420.350 640.000 ;
    END
  END dest_val0[12]
  PIN dest_val0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 427.890 636.000 428.170 640.000 ;
    END
  END dest_val0[13]
  PIN dest_val0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 435.710 636.000 435.990 640.000 ;
    END
  END dest_val0[14]
  PIN dest_val0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 443.530 636.000 443.810 640.000 ;
    END
  END dest_val0[15]
  PIN dest_val0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 451.350 636.000 451.630 640.000 ;
    END
  END dest_val0[16]
  PIN dest_val0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.673500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 459.170 636.000 459.450 640.000 ;
    END
  END dest_val0[17]
  PIN dest_val0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 466.990 636.000 467.270 640.000 ;
    END
  END dest_val0[18]
  PIN dest_val0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.673500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 474.810 636.000 475.090 640.000 ;
    END
  END dest_val0[19]
  PIN dest_val0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 334.050 636.000 334.330 640.000 ;
    END
  END dest_val0[1]
  PIN dest_val0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.673500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 482.630 636.000 482.910 640.000 ;
    END
  END dest_val0[20]
  PIN dest_val0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.673500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 490.450 636.000 490.730 640.000 ;
    END
  END dest_val0[21]
  PIN dest_val0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 498.270 636.000 498.550 640.000 ;
    END
  END dest_val0[22]
  PIN dest_val0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 506.090 636.000 506.370 640.000 ;
    END
  END dest_val0[23]
  PIN dest_val0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 513.910 636.000 514.190 640.000 ;
    END
  END dest_val0[24]
  PIN dest_val0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.639000 ;
    PORT
      LAYER met2 ;
        RECT 521.730 636.000 522.010 640.000 ;
    END
  END dest_val0[25]
  PIN dest_val0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.673500 ;
    PORT
      LAYER met2 ;
        RECT 529.550 636.000 529.830 640.000 ;
    END
  END dest_val0[26]
  PIN dest_val0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.673500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 537.370 636.000 537.650 640.000 ;
    END
  END dest_val0[27]
  PIN dest_val0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 545.190 636.000 545.470 640.000 ;
    END
  END dest_val0[28]
  PIN dest_val0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.673500 ;
    PORT
      LAYER met2 ;
        RECT 553.010 636.000 553.290 640.000 ;
    END
  END dest_val0[29]
  PIN dest_val0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 341.870 636.000 342.150 640.000 ;
    END
  END dest_val0[2]
  PIN dest_val0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 560.830 636.000 561.110 640.000 ;
    END
  END dest_val0[30]
  PIN dest_val0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 568.650 636.000 568.930 640.000 ;
    END
  END dest_val0[31]
  PIN dest_val0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 349.690 636.000 349.970 640.000 ;
    END
  END dest_val0[3]
  PIN dest_val0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 357.510 636.000 357.790 640.000 ;
    END
  END dest_val0[4]
  PIN dest_val0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.673500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 365.330 636.000 365.610 640.000 ;
    END
  END dest_val0[5]
  PIN dest_val0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.673500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 373.150 636.000 373.430 640.000 ;
    END
  END dest_val0[6]
  PIN dest_val0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.673500 ;
    PORT
      LAYER met2 ;
        RECT 380.970 636.000 381.250 640.000 ;
    END
  END dest_val0[7]
  PIN dest_val0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met2 ;
        RECT 388.790 636.000 389.070 640.000 ;
    END
  END dest_val0[8]
  PIN dest_val0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 396.610 636.000 396.890 640.000 ;
    END
  END dest_val0[9]
  PIN dest_val1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 28.600 2100.000 29.200 ;
    END
  END dest_val1[0]
  PIN dest_val1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 55.800 2100.000 56.400 ;
    END
  END dest_val1[10]
  PIN dest_val1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.673500 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 58.520 2100.000 59.120 ;
    END
  END dest_val1[11]
  PIN dest_val1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.168500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 61.240 2100.000 61.840 ;
    END
  END dest_val1[12]
  PIN dest_val1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.921000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 63.960 2100.000 64.560 ;
    END
  END dest_val1[13]
  PIN dest_val1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 66.680 2100.000 67.280 ;
    END
  END dest_val1[14]
  PIN dest_val1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 69.400 2100.000 70.000 ;
    END
  END dest_val1[15]
  PIN dest_val1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 72.120 2100.000 72.720 ;
    END
  END dest_val1[16]
  PIN dest_val1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.673500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 74.840 2100.000 75.440 ;
    END
  END dest_val1[17]
  PIN dest_val1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 77.560 2100.000 78.160 ;
    END
  END dest_val1[18]
  PIN dest_val1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 80.280 2100.000 80.880 ;
    END
  END dest_val1[19]
  PIN dest_val1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 31.320 2100.000 31.920 ;
    END
  END dest_val1[1]
  PIN dest_val1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.921000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 83.000 2100.000 83.600 ;
    END
  END dest_val1[20]
  PIN dest_val1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 85.720 2100.000 86.320 ;
    END
  END dest_val1[21]
  PIN dest_val1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 88.440 2100.000 89.040 ;
    END
  END dest_val1[22]
  PIN dest_val1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 2.173500 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 91.160 2100.000 91.760 ;
    END
  END dest_val1[23]
  PIN dest_val1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 93.880 2100.000 94.480 ;
    END
  END dest_val1[24]
  PIN dest_val1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.673500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 96.600 2100.000 97.200 ;
    END
  END dest_val1[25]
  PIN dest_val1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.673500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 99.320 2100.000 99.920 ;
    END
  END dest_val1[26]
  PIN dest_val1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.921000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 102.040 2100.000 102.640 ;
    END
  END dest_val1[27]
  PIN dest_val1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 104.760 2100.000 105.360 ;
    END
  END dest_val1[28]
  PIN dest_val1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 107.480 2100.000 108.080 ;
    END
  END dest_val1[29]
  PIN dest_val1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 34.040 2100.000 34.640 ;
    END
  END dest_val1[2]
  PIN dest_val1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 110.200 2100.000 110.800 ;
    END
  END dest_val1[30]
  PIN dest_val1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 112.920 2100.000 113.520 ;
    END
  END dest_val1[31]
  PIN dest_val1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 36.760 2100.000 37.360 ;
    END
  END dest_val1[3]
  PIN dest_val1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 39.480 2100.000 40.080 ;
    END
  END dest_val1[4]
  PIN dest_val1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 42.200 2100.000 42.800 ;
    END
  END dest_val1[5]
  PIN dest_val1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 44.920 2100.000 45.520 ;
    END
  END dest_val1[6]
  PIN dest_val1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.673500 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 47.640 2100.000 48.240 ;
    END
  END dest_val1[7]
  PIN dest_val1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 50.360 2100.000 50.960 ;
    END
  END dest_val1[8]
  PIN dest_val1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 53.080 2100.000 53.680 ;
    END
  END dest_val1[9]
  PIN dest_val2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.600 4.000 29.200 ;
    END
  END dest_val2[0]
  PIN dest_val2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 4.000 56.400 ;
    END
  END dest_val2[10]
  PIN dest_val2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 58.520 4.000 59.120 ;
    END
  END dest_val2[11]
  PIN dest_val2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END dest_val2[12]
  PIN dest_val2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 9.998099 ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.960 4.000 64.560 ;
    END
  END dest_val2[13]
  PIN dest_val2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.680 4.000 67.280 ;
    END
  END dest_val2[14]
  PIN dest_val2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.400 4.000 70.000 ;
    END
  END dest_val2[15]
  PIN dest_val2[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.120 4.000 72.720 ;
    END
  END dest_val2[16]
  PIN dest_val2[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END dest_val2[17]
  PIN dest_val2[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 77.560 4.000 78.160 ;
    END
  END dest_val2[18]
  PIN dest_val2[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.280 4.000 80.880 ;
    END
  END dest_val2[19]
  PIN dest_val2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.320 4.000 31.920 ;
    END
  END dest_val2[1]
  PIN dest_val2[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 4.000 83.600 ;
    END
  END dest_val2[20]
  PIN dest_val2[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.720 4.000 86.320 ;
    END
  END dest_val2[21]
  PIN dest_val2[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END dest_val2[22]
  PIN dest_val2[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.160 4.000 91.760 ;
    END
  END dest_val2[23]
  PIN dest_val2[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.880 4.000 94.480 ;
    END
  END dest_val2[24]
  PIN dest_val2[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.600 4.000 97.200 ;
    END
  END dest_val2[25]
  PIN dest_val2[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 99.320 4.000 99.920 ;
    END
  END dest_val2[26]
  PIN dest_val2[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END dest_val2[27]
  PIN dest_val2[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.760 4.000 105.360 ;
    END
  END dest_val2[28]
  PIN dest_val2[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 107.480 4.000 108.080 ;
    END
  END dest_val2[29]
  PIN dest_val2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END dest_val2[2]
  PIN dest_val2[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.200 4.000 110.800 ;
    END
  END dest_val2[30]
  PIN dest_val2[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.920 4.000 113.520 ;
    END
  END dest_val2[31]
  PIN dest_val2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.760 4.000 37.360 ;
    END
  END dest_val2[3]
  PIN dest_val2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 4.000 40.080 ;
    END
  END dest_val2[4]
  PIN dest_val2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.200 4.000 42.800 ;
    END
  END dest_val2[5]
  PIN dest_val2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.920 4.000 45.520 ;
    END
  END dest_val2[6]
  PIN dest_val2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.485000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END dest_val2[7]
  PIN dest_val2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.360 4.000 50.960 ;
    END
  END dest_val2[8]
  PIN dest_val2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.080 4.000 53.680 ;
    END
  END dest_val2[9]
  PIN eu0_busy
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met2 ;
        RECT 1241.170 636.000 1241.450 640.000 ;
    END
  END eu0_busy
  PIN eu0_instruction[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1248.990 636.000 1249.270 640.000 ;
    END
  END eu0_instruction[0]
  PIN eu0_instruction[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1327.190 636.000 1327.470 640.000 ;
    END
  END eu0_instruction[10]
  PIN eu0_instruction[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1335.010 636.000 1335.290 640.000 ;
    END
  END eu0_instruction[11]
  PIN eu0_instruction[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1342.830 636.000 1343.110 640.000 ;
    END
  END eu0_instruction[12]
  PIN eu0_instruction[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1350.650 636.000 1350.930 640.000 ;
    END
  END eu0_instruction[13]
  PIN eu0_instruction[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1358.470 636.000 1358.750 640.000 ;
    END
  END eu0_instruction[14]
  PIN eu0_instruction[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1366.290 636.000 1366.570 640.000 ;
    END
  END eu0_instruction[15]
  PIN eu0_instruction[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1374.110 636.000 1374.390 640.000 ;
    END
  END eu0_instruction[16]
  PIN eu0_instruction[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 1.325700 ;
    PORT
      LAYER met2 ;
        RECT 1381.930 636.000 1382.210 640.000 ;
    END
  END eu0_instruction[17]
  PIN eu0_instruction[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1389.750 636.000 1390.030 640.000 ;
    END
  END eu0_instruction[18]
  PIN eu0_instruction[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1397.570 636.000 1397.850 640.000 ;
    END
  END eu0_instruction[19]
  PIN eu0_instruction[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1256.810 636.000 1257.090 640.000 ;
    END
  END eu0_instruction[1]
  PIN eu0_instruction[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1405.390 636.000 1405.670 640.000 ;
    END
  END eu0_instruction[20]
  PIN eu0_instruction[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1413.210 636.000 1413.490 640.000 ;
    END
  END eu0_instruction[21]
  PIN eu0_instruction[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1421.030 636.000 1421.310 640.000 ;
    END
  END eu0_instruction[22]
  PIN eu0_instruction[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1428.850 636.000 1429.130 640.000 ;
    END
  END eu0_instruction[23]
  PIN eu0_instruction[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1436.670 636.000 1436.950 640.000 ;
    END
  END eu0_instruction[24]
  PIN eu0_instruction[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1444.490 636.000 1444.770 640.000 ;
    END
  END eu0_instruction[25]
  PIN eu0_instruction[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1452.310 636.000 1452.590 640.000 ;
    END
  END eu0_instruction[26]
  PIN eu0_instruction[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1460.130 636.000 1460.410 640.000 ;
    END
  END eu0_instruction[27]
  PIN eu0_instruction[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1467.950 636.000 1468.230 640.000 ;
    END
  END eu0_instruction[28]
  PIN eu0_instruction[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1475.770 636.000 1476.050 640.000 ;
    END
  END eu0_instruction[29]
  PIN eu0_instruction[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1264.630 636.000 1264.910 640.000 ;
    END
  END eu0_instruction[2]
  PIN eu0_instruction[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1483.590 636.000 1483.870 640.000 ;
    END
  END eu0_instruction[30]
  PIN eu0_instruction[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1491.410 636.000 1491.690 640.000 ;
    END
  END eu0_instruction[31]
  PIN eu0_instruction[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1499.230 636.000 1499.510 640.000 ;
    END
  END eu0_instruction[32]
  PIN eu0_instruction[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1507.050 636.000 1507.330 640.000 ;
    END
  END eu0_instruction[33]
  PIN eu0_instruction[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1514.870 636.000 1515.150 640.000 ;
    END
  END eu0_instruction[34]
  PIN eu0_instruction[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1522.690 636.000 1522.970 640.000 ;
    END
  END eu0_instruction[35]
  PIN eu0_instruction[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1530.510 636.000 1530.790 640.000 ;
    END
  END eu0_instruction[36]
  PIN eu0_instruction[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1538.330 636.000 1538.610 640.000 ;
    END
  END eu0_instruction[37]
  PIN eu0_instruction[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1546.150 636.000 1546.430 640.000 ;
    END
  END eu0_instruction[38]
  PIN eu0_instruction[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1553.970 636.000 1554.250 640.000 ;
    END
  END eu0_instruction[39]
  PIN eu0_instruction[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1272.450 636.000 1272.730 640.000 ;
    END
  END eu0_instruction[3]
  PIN eu0_instruction[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 2.629800 ;
    PORT
      LAYER met2 ;
        RECT 1561.790 636.000 1562.070 640.000 ;
    END
  END eu0_instruction[40]
  PIN eu0_instruction[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1569.610 636.000 1569.890 640.000 ;
    END
  END eu0_instruction[41]
  PIN eu0_instruction[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1280.270 636.000 1280.550 640.000 ;
    END
  END eu0_instruction[4]
  PIN eu0_instruction[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1288.090 636.000 1288.370 640.000 ;
    END
  END eu0_instruction[5]
  PIN eu0_instruction[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1295.910 636.000 1296.190 640.000 ;
    END
  END eu0_instruction[6]
  PIN eu0_instruction[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1303.730 636.000 1304.010 640.000 ;
    END
  END eu0_instruction[7]
  PIN eu0_instruction[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1311.550 636.000 1311.830 640.000 ;
    END
  END eu0_instruction[8]
  PIN eu0_instruction[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1319.370 636.000 1319.650 640.000 ;
    END
  END eu0_instruction[9]
  PIN eu1_busy
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 346.840 2100.000 347.440 ;
    END
  END eu1_busy
  PIN eu1_instruction[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 349.560 2100.000 350.160 ;
    END
  END eu1_instruction[0]
  PIN eu1_instruction[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 376.760 2100.000 377.360 ;
    END
  END eu1_instruction[10]
  PIN eu1_instruction[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 379.480 2100.000 380.080 ;
    END
  END eu1_instruction[11]
  PIN eu1_instruction[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 382.200 2100.000 382.800 ;
    END
  END eu1_instruction[12]
  PIN eu1_instruction[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 384.920 2100.000 385.520 ;
    END
  END eu1_instruction[13]
  PIN eu1_instruction[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 387.640 2100.000 388.240 ;
    END
  END eu1_instruction[14]
  PIN eu1_instruction[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 390.360 2100.000 390.960 ;
    END
  END eu1_instruction[15]
  PIN eu1_instruction[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 393.080 2100.000 393.680 ;
    END
  END eu1_instruction[16]
  PIN eu1_instruction[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 395.800 2100.000 396.400 ;
    END
  END eu1_instruction[17]
  PIN eu1_instruction[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 398.520 2100.000 399.120 ;
    END
  END eu1_instruction[18]
  PIN eu1_instruction[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 401.240 2100.000 401.840 ;
    END
  END eu1_instruction[19]
  PIN eu1_instruction[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 352.280 2100.000 352.880 ;
    END
  END eu1_instruction[1]
  PIN eu1_instruction[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 403.960 2100.000 404.560 ;
    END
  END eu1_instruction[20]
  PIN eu1_instruction[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 406.680 2100.000 407.280 ;
    END
  END eu1_instruction[21]
  PIN eu1_instruction[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 409.400 2100.000 410.000 ;
    END
  END eu1_instruction[22]
  PIN eu1_instruction[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 412.120 2100.000 412.720 ;
    END
  END eu1_instruction[23]
  PIN eu1_instruction[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 414.840 2100.000 415.440 ;
    END
  END eu1_instruction[24]
  PIN eu1_instruction[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 417.560 2100.000 418.160 ;
    END
  END eu1_instruction[25]
  PIN eu1_instruction[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 13.540500 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 420.280 2100.000 420.880 ;
    END
  END eu1_instruction[26]
  PIN eu1_instruction[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 8.397200 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 423.000 2100.000 423.600 ;
    END
  END eu1_instruction[27]
  PIN eu1_instruction[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 19.264700 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 425.720 2100.000 426.320 ;
    END
  END eu1_instruction[28]
  PIN eu1_instruction[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 10.062900 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 428.440 2100.000 429.040 ;
    END
  END eu1_instruction[29]
  PIN eu1_instruction[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 355.000 2100.000 355.600 ;
    END
  END eu1_instruction[2]
  PIN eu1_instruction[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 24.842699 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 431.160 2100.000 431.760 ;
    END
  END eu1_instruction[30]
  PIN eu1_instruction[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 13.540500 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 433.880 2100.000 434.480 ;
    END
  END eu1_instruction[31]
  PIN eu1_instruction[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 8.758800 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 436.600 2100.000 437.200 ;
    END
  END eu1_instruction[32]
  PIN eu1_instruction[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 13.540500 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 439.320 2100.000 439.920 ;
    END
  END eu1_instruction[33]
  PIN eu1_instruction[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 18.322199 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 442.040 2100.000 442.640 ;
    END
  END eu1_instruction[34]
  PIN eu1_instruction[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 20.568800 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 444.760 2100.000 445.360 ;
    END
  END eu1_instruction[35]
  PIN eu1_instruction[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 447.480 2100.000 448.080 ;
    END
  END eu1_instruction[36]
  PIN eu1_instruction[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 3.542400 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 450.200 2100.000 450.800 ;
    END
  END eu1_instruction[37]
  PIN eu1_instruction[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 452.920 2100.000 453.520 ;
    END
  END eu1_instruction[38]
  PIN eu1_instruction[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 12.671100 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 455.640 2100.000 456.240 ;
    END
  END eu1_instruction[39]
  PIN eu1_instruction[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 357.720 2100.000 358.320 ;
    END
  END eu1_instruction[3]
  PIN eu1_instruction[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 458.360 2100.000 458.960 ;
    END
  END eu1_instruction[40]
  PIN eu1_instruction[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 461.080 2100.000 461.680 ;
    END
  END eu1_instruction[41]
  PIN eu1_instruction[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 360.440 2100.000 361.040 ;
    END
  END eu1_instruction[4]
  PIN eu1_instruction[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 363.160 2100.000 363.760 ;
    END
  END eu1_instruction[5]
  PIN eu1_instruction[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 365.880 2100.000 366.480 ;
    END
  END eu1_instruction[6]
  PIN eu1_instruction[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 368.600 2100.000 369.200 ;
    END
  END eu1_instruction[7]
  PIN eu1_instruction[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 371.320 2100.000 371.920 ;
    END
  END eu1_instruction[8]
  PIN eu1_instruction[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 1.325700 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 374.040 2100.000 374.640 ;
    END
  END eu1_instruction[9]
  PIN eu2_busy
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.840 4.000 347.440 ;
    END
  END eu2_busy
  PIN eu2_instruction[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 349.560 4.000 350.160 ;
    END
  END eu2_instruction[0]
  PIN eu2_instruction[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 376.760 4.000 377.360 ;
    END
  END eu2_instruction[10]
  PIN eu2_instruction[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 379.480 4.000 380.080 ;
    END
  END eu2_instruction[11]
  PIN eu2_instruction[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 382.200 4.000 382.800 ;
    END
  END eu2_instruction[12]
  PIN eu2_instruction[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.920 4.000 385.520 ;
    END
  END eu2_instruction[13]
  PIN eu2_instruction[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 387.640 4.000 388.240 ;
    END
  END eu2_instruction[14]
  PIN eu2_instruction[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 390.360 4.000 390.960 ;
    END
  END eu2_instruction[15]
  PIN eu2_instruction[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 393.080 4.000 393.680 ;
    END
  END eu2_instruction[16]
  PIN eu2_instruction[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 395.800 4.000 396.400 ;
    END
  END eu2_instruction[17]
  PIN eu2_instruction[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 398.520 4.000 399.120 ;
    END
  END eu2_instruction[18]
  PIN eu2_instruction[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 401.240 4.000 401.840 ;
    END
  END eu2_instruction[19]
  PIN eu2_instruction[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 352.280 4.000 352.880 ;
    END
  END eu2_instruction[1]
  PIN eu2_instruction[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 403.960 4.000 404.560 ;
    END
  END eu2_instruction[20]
  PIN eu2_instruction[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 406.680 4.000 407.280 ;
    END
  END eu2_instruction[21]
  PIN eu2_instruction[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 409.400 4.000 410.000 ;
    END
  END eu2_instruction[22]
  PIN eu2_instruction[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 412.120 4.000 412.720 ;
    END
  END eu2_instruction[23]
  PIN eu2_instruction[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 414.840 4.000 415.440 ;
    END
  END eu2_instruction[24]
  PIN eu2_instruction[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 417.560 4.000 418.160 ;
    END
  END eu2_instruction[25]
  PIN eu2_instruction[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 420.280 4.000 420.880 ;
    END
  END eu2_instruction[26]
  PIN eu2_instruction[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 423.000 4.000 423.600 ;
    END
  END eu2_instruction[27]
  PIN eu2_instruction[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 425.720 4.000 426.320 ;
    END
  END eu2_instruction[28]
  PIN eu2_instruction[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 428.440 4.000 429.040 ;
    END
  END eu2_instruction[29]
  PIN eu2_instruction[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 355.000 4.000 355.600 ;
    END
  END eu2_instruction[2]
  PIN eu2_instruction[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 431.160 4.000 431.760 ;
    END
  END eu2_instruction[30]
  PIN eu2_instruction[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 433.880 4.000 434.480 ;
    END
  END eu2_instruction[31]
  PIN eu2_instruction[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 436.600 4.000 437.200 ;
    END
  END eu2_instruction[32]
  PIN eu2_instruction[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 439.320 4.000 439.920 ;
    END
  END eu2_instruction[33]
  PIN eu2_instruction[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 442.040 4.000 442.640 ;
    END
  END eu2_instruction[34]
  PIN eu2_instruction[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 444.760 4.000 445.360 ;
    END
  END eu2_instruction[35]
  PIN eu2_instruction[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 447.480 4.000 448.080 ;
    END
  END eu2_instruction[36]
  PIN eu2_instruction[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 450.200 4.000 450.800 ;
    END
  END eu2_instruction[37]
  PIN eu2_instruction[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 452.920 4.000 453.520 ;
    END
  END eu2_instruction[38]
  PIN eu2_instruction[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 455.640 4.000 456.240 ;
    END
  END eu2_instruction[39]
  PIN eu2_instruction[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.720 4.000 358.320 ;
    END
  END eu2_instruction[3]
  PIN eu2_instruction[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 458.360 4.000 458.960 ;
    END
  END eu2_instruction[40]
  PIN eu2_instruction[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 461.080 4.000 461.680 ;
    END
  END eu2_instruction[41]
  PIN eu2_instruction[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 360.440 4.000 361.040 ;
    END
  END eu2_instruction[4]
  PIN eu2_instruction[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.160 4.000 363.760 ;
    END
  END eu2_instruction[5]
  PIN eu2_instruction[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 365.880 4.000 366.480 ;
    END
  END eu2_instruction[6]
  PIN eu2_instruction[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 368.600 4.000 369.200 ;
    END
  END eu2_instruction[7]
  PIN eu2_instruction[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 371.320 4.000 371.920 ;
    END
  END eu2_instruction[8]
  PIN eu2_instruction[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.040 4.000 374.640 ;
    END
  END eu2_instruction[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 27.230 0.000 27.510 4.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.994500 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met2 ;
        RECT 206.630 0.000 206.910 4.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.751500 ;
    ANTENNADIFFAREA 2.608200 ;
    PORT
      LAYER met2 ;
        RECT 224.570 0.000 224.850 4.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.751500 ;
    ANTENNADIFFAREA 2.173500 ;
    PORT
      LAYER met2 ;
        RECT 242.510 0.000 242.790 4.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.751500 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met2 ;
        RECT 260.450 0.000 260.730 4.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.751500 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met2 ;
        RECT 278.390 0.000 278.670 4.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.751500 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met2 ;
        RECT 296.330 0.000 296.610 4.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.751500 ;
    ANTENNADIFFAREA 2.173500 ;
    PORT
      LAYER met2 ;
        RECT 314.270 0.000 314.550 4.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.246500 ;
    ANTENNADIFFAREA 3.477600 ;
    PORT
      LAYER met2 ;
        RECT 332.210 0.000 332.490 4.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.246500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 350.150 0.000 350.430 4.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.090 0.000 368.370 4.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.030 0.000 386.310 4.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.970 0.000 404.250 4.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 0.000 422.190 4.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.850 0.000 440.130 4.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.790 0.000 458.070 4.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.730 0.000 476.010 4.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER met2 ;
        RECT 493.670 0.000 493.950 4.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 511.610 0.000 511.890 4.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 529.550 0.000 529.830 4.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 547.490 0.000 547.770 4.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 63.110 0.000 63.390 4.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 565.430 0.000 565.710 4.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 583.370 0.000 583.650 4.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 601.310 0.000 601.590 4.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 619.250 0.000 619.530 4.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 637.190 0.000 637.470 4.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 655.130 0.000 655.410 4.000 ;
    END
  END io_in[35]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.994500 ;
    ANTENNADIFFAREA 2.608200 ;
    PORT
      LAYER met2 ;
        RECT 81.050 0.000 81.330 4.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.994500 ;
    ANTENNADIFFAREA 2.608200 ;
    PORT
      LAYER met2 ;
        RECT 98.990 0.000 99.270 4.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.994500 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met2 ;
        RECT 116.930 0.000 117.210 4.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.994500 ;
    ANTENNADIFFAREA 2.608200 ;
    PORT
      LAYER met2 ;
        RECT 134.870 0.000 135.150 4.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.994500 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met2 ;
        RECT 152.810 0.000 153.090 4.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.994500 ;
    ANTENNADIFFAREA 2.608200 ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 4.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.994500 ;
    ANTENNADIFFAREA 2.173500 ;
    PORT
      LAYER met2 ;
        RECT 188.690 0.000 188.970 4.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.484000 ;
    PORT
      LAYER met2 ;
        RECT 673.070 0.000 673.350 4.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 852.470 0.000 852.750 4.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 870.410 0.000 870.690 4.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 888.350 0.000 888.630 4.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 906.290 0.000 906.570 4.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 924.230 0.000 924.510 4.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 942.170 0.000 942.450 4.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 960.110 0.000 960.390 4.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 978.050 0.000 978.330 4.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 13.860000 ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 995.990 0.000 996.270 4.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.930 0.000 1014.210 4.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 691.010 0.000 691.290 4.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1031.870 0.000 1032.150 4.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1049.810 0.000 1050.090 4.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1067.750 0.000 1068.030 4.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1085.690 0.000 1085.970 4.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1103.630 0.000 1103.910 4.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1121.570 0.000 1121.850 4.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1139.510 0.000 1139.790 4.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1157.450 0.000 1157.730 4.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1175.390 0.000 1175.670 4.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1193.330 0.000 1193.610 4.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.484000 ;
    PORT
      LAYER met2 ;
        RECT 708.950 0.000 709.230 4.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 6.172200 ;
    PORT
      LAYER met2 ;
        RECT 1211.270 0.000 1211.550 4.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1229.210 0.000 1229.490 4.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1247.150 0.000 1247.430 4.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1265.090 0.000 1265.370 4.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1283.030 0.000 1283.310 4.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1300.970 0.000 1301.250 4.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 726.890 0.000 727.170 4.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 744.830 0.000 745.110 4.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 762.770 0.000 763.050 4.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 780.710 0.000 780.990 4.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 798.650 0.000 798.930 4.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 816.590 0.000 816.870 4.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 834.530 0.000 834.810 4.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1318.910 0.000 1319.190 4.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1498.310 0.000 1498.590 4.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1516.250 0.000 1516.530 4.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1534.190 0.000 1534.470 4.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1552.130 0.000 1552.410 4.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1570.070 0.000 1570.350 4.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1588.010 0.000 1588.290 4.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1605.950 0.000 1606.230 4.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1623.890 0.000 1624.170 4.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.484000 ;
    PORT
      LAYER met2 ;
        RECT 1641.830 0.000 1642.110 4.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1659.770 0.000 1660.050 4.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1336.850 0.000 1337.130 4.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1677.710 0.000 1677.990 4.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1695.650 0.000 1695.930 4.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1713.590 0.000 1713.870 4.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1731.530 0.000 1731.810 4.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.715500 ;
    PORT
      LAYER met2 ;
        RECT 1749.470 0.000 1749.750 4.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1767.410 0.000 1767.690 4.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1785.350 0.000 1785.630 4.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1803.290 0.000 1803.570 4.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1821.230 0.000 1821.510 4.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1839.170 0.000 1839.450 4.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1354.790 0.000 1355.070 4.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 10.454400 ;
    PORT
      LAYER met2 ;
        RECT 1857.110 0.000 1857.390 4.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1875.050 0.000 1875.330 4.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 3.499200 ;
    PORT
      LAYER met2 ;
        RECT 1892.990 0.000 1893.270 4.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 6.107400 ;
    PORT
      LAYER met2 ;
        RECT 1910.930 0.000 1911.210 4.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 12.236400 ;
    PORT
      LAYER met2 ;
        RECT 1928.870 0.000 1929.150 4.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1946.810 0.000 1947.090 4.000 ;
    END
  END io_out[35]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1372.730 0.000 1373.010 4.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1390.670 0.000 1390.950 4.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1408.610 0.000 1408.890 4.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1426.550 0.000 1426.830 4.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1444.490 0.000 1444.770 4.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1462.430 0.000 1462.710 4.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1480.370 0.000 1480.650 4.000 ;
    END
  END io_out[9]
  PIN is_load0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met2 ;
        RECT 936.190 636.000 936.470 640.000 ;
    END
  END is_load0
  PIN is_load1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.621000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 240.760 2100.000 241.360 ;
    END
  END is_load1
  PIN is_load2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.760 4.000 241.360 ;
    END
  END is_load2
  PIN is_store0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.237500 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met2 ;
        RECT 944.010 636.000 944.290 640.000 ;
    END
  END is_store0
  PIN is_store1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.868500 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 243.480 2100.000 244.080 ;
    END
  END is_store1
  PIN is_store2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 10.867499 ;
    PORT
      LAYER met3 ;
        RECT 0.000 243.480 4.000 244.080 ;
    END
  END is_store2
  PIN loadstore_address0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 685.950 636.000 686.230 640.000 ;
    END
  END loadstore_address0[0]
  PIN loadstore_address0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 764.150 636.000 764.430 640.000 ;
    END
  END loadstore_address0[10]
  PIN loadstore_address0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 771.970 636.000 772.250 640.000 ;
    END
  END loadstore_address0[11]
  PIN loadstore_address0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 779.790 636.000 780.070 640.000 ;
    END
  END loadstore_address0[12]
  PIN loadstore_address0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 787.610 636.000 787.890 640.000 ;
    END
  END loadstore_address0[13]
  PIN loadstore_address0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 795.430 636.000 795.710 640.000 ;
    END
  END loadstore_address0[14]
  PIN loadstore_address0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 803.250 636.000 803.530 640.000 ;
    END
  END loadstore_address0[15]
  PIN loadstore_address0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 811.070 636.000 811.350 640.000 ;
    END
  END loadstore_address0[16]
  PIN loadstore_address0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 818.890 636.000 819.170 640.000 ;
    END
  END loadstore_address0[17]
  PIN loadstore_address0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 826.710 636.000 826.990 640.000 ;
    END
  END loadstore_address0[18]
  PIN loadstore_address0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 834.530 636.000 834.810 640.000 ;
    END
  END loadstore_address0[19]
  PIN loadstore_address0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met2 ;
        RECT 693.770 636.000 694.050 640.000 ;
    END
  END loadstore_address0[1]
  PIN loadstore_address0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 842.350 636.000 842.630 640.000 ;
    END
  END loadstore_address0[20]
  PIN loadstore_address0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 850.170 636.000 850.450 640.000 ;
    END
  END loadstore_address0[21]
  PIN loadstore_address0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 857.990 636.000 858.270 640.000 ;
    END
  END loadstore_address0[22]
  PIN loadstore_address0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 865.810 636.000 866.090 640.000 ;
    END
  END loadstore_address0[23]
  PIN loadstore_address0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 873.630 636.000 873.910 640.000 ;
    END
  END loadstore_address0[24]
  PIN loadstore_address0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 881.450 636.000 881.730 640.000 ;
    END
  END loadstore_address0[25]
  PIN loadstore_address0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 889.270 636.000 889.550 640.000 ;
    END
  END loadstore_address0[26]
  PIN loadstore_address0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 897.090 636.000 897.370 640.000 ;
    END
  END loadstore_address0[27]
  PIN loadstore_address0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 904.910 636.000 905.190 640.000 ;
    END
  END loadstore_address0[28]
  PIN loadstore_address0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 912.730 636.000 913.010 640.000 ;
    END
  END loadstore_address0[29]
  PIN loadstore_address0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 701.590 636.000 701.870 640.000 ;
    END
  END loadstore_address0[2]
  PIN loadstore_address0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 920.550 636.000 920.830 640.000 ;
    END
  END loadstore_address0[30]
  PIN loadstore_address0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 928.370 636.000 928.650 640.000 ;
    END
  END loadstore_address0[31]
  PIN loadstore_address0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 709.410 636.000 709.690 640.000 ;
    END
  END loadstore_address0[3]
  PIN loadstore_address0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 717.230 636.000 717.510 640.000 ;
    END
  END loadstore_address0[4]
  PIN loadstore_address0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 725.050 636.000 725.330 640.000 ;
    END
  END loadstore_address0[5]
  PIN loadstore_address0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 732.870 636.000 733.150 640.000 ;
    END
  END loadstore_address0[6]
  PIN loadstore_address0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 740.690 636.000 740.970 640.000 ;
    END
  END loadstore_address0[7]
  PIN loadstore_address0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 748.510 636.000 748.790 640.000 ;
    END
  END loadstore_address0[8]
  PIN loadstore_address0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 756.330 636.000 756.610 640.000 ;
    END
  END loadstore_address0[9]
  PIN loadstore_address1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 153.720 2100.000 154.320 ;
    END
  END loadstore_address1[0]
  PIN loadstore_address1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 180.920 2100.000 181.520 ;
    END
  END loadstore_address1[10]
  PIN loadstore_address1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 183.640 2100.000 184.240 ;
    END
  END loadstore_address1[11]
  PIN loadstore_address1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 186.360 2100.000 186.960 ;
    END
  END loadstore_address1[12]
  PIN loadstore_address1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 20.430899 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 189.080 2100.000 189.680 ;
    END
  END loadstore_address1[13]
  PIN loadstore_address1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 20.430899 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 191.800 2100.000 192.400 ;
    END
  END loadstore_address1[14]
  PIN loadstore_address1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 9.998099 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 194.520 2100.000 195.120 ;
    END
  END loadstore_address1[15]
  PIN loadstore_address1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 20.430899 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 197.240 2100.000 197.840 ;
    END
  END loadstore_address1[16]
  PIN loadstore_address1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 22.169699 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 199.960 2100.000 200.560 ;
    END
  END loadstore_address1[17]
  PIN loadstore_address1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 9.998099 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 202.680 2100.000 203.280 ;
    END
  END loadstore_address1[18]
  PIN loadstore_address1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 205.400 2100.000 206.000 ;
    END
  END loadstore_address1[19]
  PIN loadstore_address1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 156.440 2100.000 157.040 ;
    END
  END loadstore_address1[1]
  PIN loadstore_address1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 208.120 2100.000 208.720 ;
    END
  END loadstore_address1[20]
  PIN loadstore_address1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 210.840 2100.000 211.440 ;
    END
  END loadstore_address1[21]
  PIN loadstore_address1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 30.863699 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 213.560 2100.000 214.160 ;
    END
  END loadstore_address1[22]
  PIN loadstore_address1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 8.694000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 216.280 2100.000 216.880 ;
    END
  END loadstore_address1[23]
  PIN loadstore_address1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 219.000 2100.000 219.600 ;
    END
  END loadstore_address1[24]
  PIN loadstore_address1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 221.720 2100.000 222.320 ;
    END
  END loadstore_address1[25]
  PIN loadstore_address1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 9.998099 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 224.440 2100.000 225.040 ;
    END
  END loadstore_address1[26]
  PIN loadstore_address1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 227.160 2100.000 227.760 ;
    END
  END loadstore_address1[27]
  PIN loadstore_address1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 229.880 2100.000 230.480 ;
    END
  END loadstore_address1[28]
  PIN loadstore_address1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 232.600 2100.000 233.200 ;
    END
  END loadstore_address1[29]
  PIN loadstore_address1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 159.160 2100.000 159.760 ;
    END
  END loadstore_address1[2]
  PIN loadstore_address1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 235.320 2100.000 235.920 ;
    END
  END loadstore_address1[30]
  PIN loadstore_address1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 238.040 2100.000 238.640 ;
    END
  END loadstore_address1[31]
  PIN loadstore_address1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 161.880 2100.000 162.480 ;
    END
  END loadstore_address1[3]
  PIN loadstore_address1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 164.600 2100.000 165.200 ;
    END
  END loadstore_address1[4]
  PIN loadstore_address1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 167.320 2100.000 167.920 ;
    END
  END loadstore_address1[5]
  PIN loadstore_address1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 170.040 2100.000 170.640 ;
    END
  END loadstore_address1[6]
  PIN loadstore_address1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 172.760 2100.000 173.360 ;
    END
  END loadstore_address1[7]
  PIN loadstore_address1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 9.998099 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 175.480 2100.000 176.080 ;
    END
  END loadstore_address1[8]
  PIN loadstore_address1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 178.200 2100.000 178.800 ;
    END
  END loadstore_address1[9]
  PIN loadstore_address2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.720 4.000 154.320 ;
    END
  END loadstore_address2[0]
  PIN loadstore_address2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.920 4.000 181.520 ;
    END
  END loadstore_address2[10]
  PIN loadstore_address2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END loadstore_address2[11]
  PIN loadstore_address2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 186.360 4.000 186.960 ;
    END
  END loadstore_address2[12]
  PIN loadstore_address2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 3.477600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.080 4.000 189.680 ;
    END
  END loadstore_address2[13]
  PIN loadstore_address2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 6.085800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.800 4.000 192.400 ;
    END
  END loadstore_address2[14]
  PIN loadstore_address2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 7.389900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 194.520 4.000 195.120 ;
    END
  END loadstore_address2[15]
  PIN loadstore_address2[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.347000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.240 4.000 197.840 ;
    END
  END loadstore_address2[16]
  PIN loadstore_address2[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 199.960 4.000 200.560 ;
    END
  END loadstore_address2[17]
  PIN loadstore_address2[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 3.912300 ;
    PORT
      LAYER met3 ;
        RECT 0.000 202.680 4.000 203.280 ;
    END
  END loadstore_address2[18]
  PIN loadstore_address2[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 205.400 4.000 206.000 ;
    END
  END loadstore_address2[19]
  PIN loadstore_address2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 3.912300 ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END loadstore_address2[1]
  PIN loadstore_address2[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 208.120 4.000 208.720 ;
    END
  END loadstore_address2[20]
  PIN loadstore_address2[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 3.912300 ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.840 4.000 211.440 ;
    END
  END loadstore_address2[21]
  PIN loadstore_address2[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.347000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 213.560 4.000 214.160 ;
    END
  END loadstore_address2[22]
  PIN loadstore_address2[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 3.912300 ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.280 4.000 216.880 ;
    END
  END loadstore_address2[23]
  PIN loadstore_address2[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 7.824600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.000 4.000 219.600 ;
    END
  END loadstore_address2[24]
  PIN loadstore_address2[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 3.912300 ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.720 4.000 222.320 ;
    END
  END loadstore_address2[25]
  PIN loadstore_address2[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.440 4.000 225.040 ;
    END
  END loadstore_address2[26]
  PIN loadstore_address2[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.160 4.000 227.760 ;
    END
  END loadstore_address2[27]
  PIN loadstore_address2[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.347000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.880 4.000 230.480 ;
    END
  END loadstore_address2[28]
  PIN loadstore_address2[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 232.600 4.000 233.200 ;
    END
  END loadstore_address2[29]
  PIN loadstore_address2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 3.912300 ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.160 4.000 159.760 ;
    END
  END loadstore_address2[2]
  PIN loadstore_address2[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 235.320 4.000 235.920 ;
    END
  END loadstore_address2[30]
  PIN loadstore_address2[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.040 4.000 238.640 ;
    END
  END loadstore_address2[31]
  PIN loadstore_address2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.347000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.880 4.000 162.480 ;
    END
  END loadstore_address2[3]
  PIN loadstore_address2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 164.600 4.000 165.200 ;
    END
  END loadstore_address2[4]
  PIN loadstore_address2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 167.320 4.000 167.920 ;
    END
  END loadstore_address2[5]
  PIN loadstore_address2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END loadstore_address2[6]
  PIN loadstore_address2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.760 4.000 173.360 ;
    END
  END loadstore_address2[7]
  PIN loadstore_address2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 175.480 4.000 176.080 ;
    END
  END loadstore_address2[8]
  PIN loadstore_address2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.200 4.000 178.800 ;
    END
  END loadstore_address2[9]
  PIN loadstore_dest0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 975.290 636.000 975.570 640.000 ;
    END
  END loadstore_dest0[0]
  PIN loadstore_dest0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met2 ;
        RECT 983.110 636.000 983.390 640.000 ;
    END
  END loadstore_dest0[1]
  PIN loadstore_dest0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met2 ;
        RECT 990.930 636.000 991.210 640.000 ;
    END
  END loadstore_dest0[2]
  PIN loadstore_dest0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met2 ;
        RECT 998.750 636.000 999.030 640.000 ;
    END
  END loadstore_dest0[3]
  PIN loadstore_dest0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met2 ;
        RECT 1006.570 636.000 1006.850 640.000 ;
    END
  END loadstore_dest0[4]
  PIN loadstore_dest1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 254.360 2100.000 254.960 ;
    END
  END loadstore_dest1[0]
  PIN loadstore_dest1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 257.080 2100.000 257.680 ;
    END
  END loadstore_dest1[1]
  PIN loadstore_dest1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.237500 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 259.800 2100.000 260.400 ;
    END
  END loadstore_dest1[2]
  PIN loadstore_dest1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.485000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 262.520 2100.000 263.120 ;
    END
  END loadstore_dest1[3]
  PIN loadstore_dest1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.485000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 265.240 2100.000 265.840 ;
    END
  END loadstore_dest1[4]
  PIN loadstore_dest2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 0.000 254.360 4.000 254.960 ;
    END
  END loadstore_dest2[0]
  PIN loadstore_dest2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 257.080 4.000 257.680 ;
    END
  END loadstore_dest2[1]
  PIN loadstore_dest2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.237500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.800 4.000 260.400 ;
    END
  END loadstore_dest2[2]
  PIN loadstore_dest2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.485000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 262.520 4.000 263.120 ;
    END
  END loadstore_dest2[3]
  PIN loadstore_dest2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.485000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.240 4.000 265.840 ;
    END
  END loadstore_dest2[4]
  PIN loadstore_size0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 959.650 636.000 959.930 640.000 ;
    END
  END loadstore_size0[0]
  PIN loadstore_size0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 967.470 636.000 967.750 640.000 ;
    END
  END loadstore_size0[1]
  PIN loadstore_size1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 248.920 2100.000 249.520 ;
    END
  END loadstore_size1[0]
  PIN loadstore_size1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 251.640 2100.000 252.240 ;
    END
  END loadstore_size1[1]
  PIN loadstore_size2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.920 4.000 249.520 ;
    END
  END loadstore_size2[0]
  PIN loadstore_size2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 9.998099 ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.640 4.000 252.240 ;
    END
  END loadstore_size2[1]
  PIN new_PC0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met2 ;
        RECT 1022.210 636.000 1022.490 640.000 ;
    END
  END new_PC0[0]
  PIN new_PC0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 5.216400 ;
    PORT
      LAYER met2 ;
        RECT 1100.410 636.000 1100.690 640.000 ;
    END
  END new_PC0[10]
  PIN new_PC0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1108.230 636.000 1108.510 640.000 ;
    END
  END new_PC0[11]
  PIN new_PC0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1116.050 636.000 1116.330 640.000 ;
    END
  END new_PC0[12]
  PIN new_PC0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1123.870 636.000 1124.150 640.000 ;
    END
  END new_PC0[13]
  PIN new_PC0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1131.690 636.000 1131.970 640.000 ;
    END
  END new_PC0[14]
  PIN new_PC0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 2.173500 ;
    PORT
      LAYER met2 ;
        RECT 1139.510 636.000 1139.790 640.000 ;
    END
  END new_PC0[15]
  PIN new_PC0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1147.330 636.000 1147.610 640.000 ;
    END
  END new_PC0[16]
  PIN new_PC0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.485000 ;
    PORT
      LAYER met2 ;
        RECT 1155.150 636.000 1155.430 640.000 ;
    END
  END new_PC0[17]
  PIN new_PC0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.485000 ;
    PORT
      LAYER met2 ;
        RECT 1162.970 636.000 1163.250 640.000 ;
    END
  END new_PC0[18]
  PIN new_PC0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 5.651100 ;
    PORT
      LAYER met2 ;
        RECT 1170.790 636.000 1171.070 640.000 ;
    END
  END new_PC0[19]
  PIN new_PC0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1030.030 636.000 1030.310 640.000 ;
    END
  END new_PC0[1]
  PIN new_PC0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.485000 ;
    PORT
      LAYER met2 ;
        RECT 1178.610 636.000 1178.890 640.000 ;
    END
  END new_PC0[20]
  PIN new_PC0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 5.651100 ;
    PORT
      LAYER met2 ;
        RECT 1186.430 636.000 1186.710 640.000 ;
    END
  END new_PC0[21]
  PIN new_PC0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met2 ;
        RECT 1194.250 636.000 1194.530 640.000 ;
    END
  END new_PC0[22]
  PIN new_PC0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 3.477600 ;
    PORT
      LAYER met2 ;
        RECT 1202.070 636.000 1202.350 640.000 ;
    END
  END new_PC0[23]
  PIN new_PC0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 5.651100 ;
    PORT
      LAYER met2 ;
        RECT 1209.890 636.000 1210.170 640.000 ;
    END
  END new_PC0[24]
  PIN new_PC0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.980000 ;
    PORT
      LAYER met2 ;
        RECT 1217.710 636.000 1217.990 640.000 ;
    END
  END new_PC0[25]
  PIN new_PC0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met2 ;
        RECT 1225.530 636.000 1225.810 640.000 ;
    END
  END new_PC0[26]
  PIN new_PC0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.304000 ;
    PORT
      LAYER met2 ;
        RECT 1233.350 636.000 1233.630 640.000 ;
    END
  END new_PC0[27]
  PIN new_PC0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1037.850 636.000 1038.130 640.000 ;
    END
  END new_PC0[2]
  PIN new_PC0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met2 ;
        RECT 1045.670 636.000 1045.950 640.000 ;
    END
  END new_PC0[3]
  PIN new_PC0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1053.490 636.000 1053.770 640.000 ;
    END
  END new_PC0[4]
  PIN new_PC0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 4.347000 ;
    PORT
      LAYER met2 ;
        RECT 1061.310 636.000 1061.590 640.000 ;
    END
  END new_PC0[5]
  PIN new_PC0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 7.389900 ;
    PORT
      LAYER met2 ;
        RECT 1069.130 636.000 1069.410 640.000 ;
    END
  END new_PC0[6]
  PIN new_PC0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1076.950 636.000 1077.230 640.000 ;
    END
  END new_PC0[7]
  PIN new_PC0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1084.770 636.000 1085.050 640.000 ;
    END
  END new_PC0[8]
  PIN new_PC0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 6.955200 ;
    PORT
      LAYER met2 ;
        RECT 1092.590 636.000 1092.870 640.000 ;
    END
  END new_PC0[9]
  PIN new_PC1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 270.680 2100.000 271.280 ;
    END
  END new_PC1[0]
  PIN new_PC1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 297.880 2100.000 298.480 ;
    END
  END new_PC1[10]
  PIN new_PC1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 5.216400 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 300.600 2100.000 301.200 ;
    END
  END new_PC1[11]
  PIN new_PC1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 303.320 2100.000 303.920 ;
    END
  END new_PC1[12]
  PIN new_PC1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 306.040 2100.000 306.640 ;
    END
  END new_PC1[13]
  PIN new_PC1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 5.216400 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 308.760 2100.000 309.360 ;
    END
  END new_PC1[14]
  PIN new_PC1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 311.480 2100.000 312.080 ;
    END
  END new_PC1[15]
  PIN new_PC1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 314.200 2100.000 314.800 ;
    END
  END new_PC1[16]
  PIN new_PC1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 316.920 2100.000 317.520 ;
    END
  END new_PC1[17]
  PIN new_PC1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 24.343199 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 319.640 2100.000 320.240 ;
    END
  END new_PC1[18]
  PIN new_PC1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 322.360 2100.000 322.960 ;
    END
  END new_PC1[19]
  PIN new_PC1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 273.400 2100.000 274.000 ;
    END
  END new_PC1[1]
  PIN new_PC1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 5.651100 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 325.080 2100.000 325.680 ;
    END
  END new_PC1[20]
  PIN new_PC1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 327.800 2100.000 328.400 ;
    END
  END new_PC1[21]
  PIN new_PC1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 330.520 2100.000 331.120 ;
    END
  END new_PC1[22]
  PIN new_PC1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 333.240 2100.000 333.840 ;
    END
  END new_PC1[23]
  PIN new_PC1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 335.960 2100.000 336.560 ;
    END
  END new_PC1[24]
  PIN new_PC1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 5.216400 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 338.680 2100.000 339.280 ;
    END
  END new_PC1[25]
  PIN new_PC1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 341.400 2100.000 342.000 ;
    END
  END new_PC1[26]
  PIN new_PC1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 19.126799 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 344.120 2100.000 344.720 ;
    END
  END new_PC1[27]
  PIN new_PC1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 276.120 2100.000 276.720 ;
    END
  END new_PC1[2]
  PIN new_PC1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 278.840 2100.000 279.440 ;
    END
  END new_PC1[3]
  PIN new_PC1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 281.560 2100.000 282.160 ;
    END
  END new_PC1[4]
  PIN new_PC1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 284.280 2100.000 284.880 ;
    END
  END new_PC1[5]
  PIN new_PC1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 287.000 2100.000 287.600 ;
    END
  END new_PC1[6]
  PIN new_PC1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 289.720 2100.000 290.320 ;
    END
  END new_PC1[7]
  PIN new_PC1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 292.440 2100.000 293.040 ;
    END
  END new_PC1[8]
  PIN new_PC1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 295.160 2100.000 295.760 ;
    END
  END new_PC1[9]
  PIN new_PC2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 3.477600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 270.680 4.000 271.280 ;
    END
  END new_PC2[0]
  PIN new_PC2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 297.880 4.000 298.480 ;
    END
  END new_PC2[10]
  PIN new_PC2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 300.600 4.000 301.200 ;
    END
  END new_PC2[11]
  PIN new_PC2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 303.320 4.000 303.920 ;
    END
  END new_PC2[12]
  PIN new_PC2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.040 4.000 306.640 ;
    END
  END new_PC2[13]
  PIN new_PC2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 308.760 4.000 309.360 ;
    END
  END new_PC2[14]
  PIN new_PC2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 311.480 4.000 312.080 ;
    END
  END new_PC2[15]
  PIN new_PC2[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 314.200 4.000 314.800 ;
    END
  END new_PC2[16]
  PIN new_PC2[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.920 4.000 317.520 ;
    END
  END new_PC2[17]
  PIN new_PC2[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 319.640 4.000 320.240 ;
    END
  END new_PC2[18]
  PIN new_PC2[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 322.360 4.000 322.960 ;
    END
  END new_PC2[19]
  PIN new_PC2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 273.400 4.000 274.000 ;
    END
  END new_PC2[1]
  PIN new_PC2[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 325.080 4.000 325.680 ;
    END
  END new_PC2[20]
  PIN new_PC2[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 327.800 4.000 328.400 ;
    END
  END new_PC2[21]
  PIN new_PC2[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 330.520 4.000 331.120 ;
    END
  END new_PC2[22]
  PIN new_PC2[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.240 4.000 333.840 ;
    END
  END new_PC2[23]
  PIN new_PC2[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 335.960 4.000 336.560 ;
    END
  END new_PC2[24]
  PIN new_PC2[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 338.680 4.000 339.280 ;
    END
  END new_PC2[25]
  PIN new_PC2[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 341.400 4.000 342.000 ;
    END
  END new_PC2[26]
  PIN new_PC2[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 344.120 4.000 344.720 ;
    END
  END new_PC2[27]
  PIN new_PC2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 276.120 4.000 276.720 ;
    END
  END new_PC2[2]
  PIN new_PC2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.840 4.000 279.440 ;
    END
  END new_PC2[3]
  PIN new_PC2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 281.560 4.000 282.160 ;
    END
  END new_PC2[4]
  PIN new_PC2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 284.280 4.000 284.880 ;
    END
  END new_PC2[5]
  PIN new_PC2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 287.000 4.000 287.600 ;
    END
  END new_PC2[6]
  PIN new_PC2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.720 4.000 290.320 ;
    END
  END new_PC2[7]
  PIN new_PC2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.440 4.000 293.040 ;
    END
  END new_PC2[8]
  PIN new_PC2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.160 4.000 295.760 ;
    END
  END new_PC2[9]
  PIN pred_idx0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.504000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 631.210 636.000 631.490 640.000 ;
    END
  END pred_idx0[0]
  PIN pred_idx0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.756000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 639.030 636.000 639.310 640.000 ;
    END
  END pred_idx0[1]
  PIN pred_idx0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 646.850 636.000 647.130 640.000 ;
    END
  END pred_idx0[2]
  PIN pred_idx1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.504000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 134.680 2100.000 135.280 ;
    END
  END pred_idx1[0]
  PIN pred_idx1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.756000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 137.400 2100.000 138.000 ;
    END
  END pred_idx1[1]
  PIN pred_idx1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 140.120 2100.000 140.720 ;
    END
  END pred_idx1[2]
  PIN pred_idx2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.504000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.680 4.000 135.280 ;
    END
  END pred_idx2[0]
  PIN pred_idx2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.756000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.400 4.000 138.000 ;
    END
  END pred_idx2[1]
  PIN pred_idx2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.120 4.000 140.720 ;
    END
  END pred_idx2[2]
  PIN pred_val0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.962500 ;
    PORT
      LAYER met2 ;
        RECT 2077.910 636.000 2078.190 640.000 ;
    END
  END pred_val0
  PIN pred_val1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.962500 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 637.880 2100.000 638.480 ;
    END
  END pred_val1
  PIN pred_val2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.962500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 637.880 4.000 638.480 ;
    END
  END pred_val2
  PIN reg1_idx0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.980000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 248.030 636.000 248.310 640.000 ;
    END
  END reg1_idx0[0]
  PIN reg1_idx0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.980000 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met2 ;
        RECT 255.850 636.000 256.130 640.000 ;
    END
  END reg1_idx0[1]
  PIN reg1_idx0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 263.670 636.000 263.950 640.000 ;
    END
  END reg1_idx0[2]
  PIN reg1_idx0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.383000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 271.490 636.000 271.770 640.000 ;
    END
  END reg1_idx0[3]
  PIN reg1_idx0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.293000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 279.310 636.000 279.590 640.000 ;
    END
  END reg1_idx0[4]
  PIN reg1_idx1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 1.400 2100.000 2.000 ;
    END
  END reg1_idx1[0]
  PIN reg1_idx1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.732500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 4.120 2100.000 4.720 ;
    END
  END reg1_idx1[1]
  PIN reg1_idx1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.327000 ;
    ANTENNADIFFAREA 2.173500 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 6.840 2100.000 7.440 ;
    END
  END reg1_idx1[2]
  PIN reg1_idx1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.980000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 9.560 2100.000 10.160 ;
    END
  END reg1_idx1[3]
  PIN reg1_idx1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.980000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 12.280 2100.000 12.880 ;
    END
  END reg1_idx1[4]
  PIN reg1_idx2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.678000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1.400 4.000 2.000 ;
    END
  END reg1_idx2[0]
  PIN reg1_idx2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.130000 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.120 4.000 4.720 ;
    END
  END reg1_idx2[1]
  PIN reg1_idx2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.327000 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END reg1_idx2[2]
  PIN reg1_idx2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.383000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 9.560 4.000 10.160 ;
    END
  END reg1_idx2[3]
  PIN reg1_idx2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.293000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 4.000 12.880 ;
    END
  END reg1_idx2[4]
  PIN reg1_val0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1577.430 636.000 1577.710 640.000 ;
    END
  END reg1_val0[0]
  PIN reg1_val0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1655.630 636.000 1655.910 640.000 ;
    END
  END reg1_val0[10]
  PIN reg1_val0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1663.450 636.000 1663.730 640.000 ;
    END
  END reg1_val0[11]
  PIN reg1_val0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1671.270 636.000 1671.550 640.000 ;
    END
  END reg1_val0[12]
  PIN reg1_val0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1679.090 636.000 1679.370 640.000 ;
    END
  END reg1_val0[13]
  PIN reg1_val0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1686.910 636.000 1687.190 640.000 ;
    END
  END reg1_val0[14]
  PIN reg1_val0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1694.730 636.000 1695.010 640.000 ;
    END
  END reg1_val0[15]
  PIN reg1_val0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1702.550 636.000 1702.830 640.000 ;
    END
  END reg1_val0[16]
  PIN reg1_val0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1710.370 636.000 1710.650 640.000 ;
    END
  END reg1_val0[17]
  PIN reg1_val0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1718.190 636.000 1718.470 640.000 ;
    END
  END reg1_val0[18]
  PIN reg1_val0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1726.010 636.000 1726.290 640.000 ;
    END
  END reg1_val0[19]
  PIN reg1_val0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1585.250 636.000 1585.530 640.000 ;
    END
  END reg1_val0[1]
  PIN reg1_val0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1733.830 636.000 1734.110 640.000 ;
    END
  END reg1_val0[20]
  PIN reg1_val0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1741.650 636.000 1741.930 640.000 ;
    END
  END reg1_val0[21]
  PIN reg1_val0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1749.470 636.000 1749.750 640.000 ;
    END
  END reg1_val0[22]
  PIN reg1_val0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1757.290 636.000 1757.570 640.000 ;
    END
  END reg1_val0[23]
  PIN reg1_val0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1765.110 636.000 1765.390 640.000 ;
    END
  END reg1_val0[24]
  PIN reg1_val0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1772.930 636.000 1773.210 640.000 ;
    END
  END reg1_val0[25]
  PIN reg1_val0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1780.750 636.000 1781.030 640.000 ;
    END
  END reg1_val0[26]
  PIN reg1_val0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1788.570 636.000 1788.850 640.000 ;
    END
  END reg1_val0[27]
  PIN reg1_val0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1796.390 636.000 1796.670 640.000 ;
    END
  END reg1_val0[28]
  PIN reg1_val0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1804.210 636.000 1804.490 640.000 ;
    END
  END reg1_val0[29]
  PIN reg1_val0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1593.070 636.000 1593.350 640.000 ;
    END
  END reg1_val0[2]
  PIN reg1_val0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1812.030 636.000 1812.310 640.000 ;
    END
  END reg1_val0[30]
  PIN reg1_val0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1819.850 636.000 1820.130 640.000 ;
    END
  END reg1_val0[31]
  PIN reg1_val0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1600.890 636.000 1601.170 640.000 ;
    END
  END reg1_val0[3]
  PIN reg1_val0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1608.710 636.000 1608.990 640.000 ;
    END
  END reg1_val0[4]
  PIN reg1_val0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1616.530 636.000 1616.810 640.000 ;
    END
  END reg1_val0[5]
  PIN reg1_val0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1624.350 636.000 1624.630 640.000 ;
    END
  END reg1_val0[6]
  PIN reg1_val0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1632.170 636.000 1632.450 640.000 ;
    END
  END reg1_val0[7]
  PIN reg1_val0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1639.990 636.000 1640.270 640.000 ;
    END
  END reg1_val0[8]
  PIN reg1_val0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1647.810 636.000 1648.090 640.000 ;
    END
  END reg1_val0[9]
  PIN reg1_val1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 463.800 2100.000 464.400 ;
    END
  END reg1_val1[0]
  PIN reg1_val1[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 491.000 2100.000 491.600 ;
    END
  END reg1_val1[10]
  PIN reg1_val1[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 493.720 2100.000 494.320 ;
    END
  END reg1_val1[11]
  PIN reg1_val1[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 496.440 2100.000 497.040 ;
    END
  END reg1_val1[12]
  PIN reg1_val1[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 499.160 2100.000 499.760 ;
    END
  END reg1_val1[13]
  PIN reg1_val1[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 501.880 2100.000 502.480 ;
    END
  END reg1_val1[14]
  PIN reg1_val1[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 504.600 2100.000 505.200 ;
    END
  END reg1_val1[15]
  PIN reg1_val1[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 507.320 2100.000 507.920 ;
    END
  END reg1_val1[16]
  PIN reg1_val1[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 510.040 2100.000 510.640 ;
    END
  END reg1_val1[17]
  PIN reg1_val1[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 512.760 2100.000 513.360 ;
    END
  END reg1_val1[18]
  PIN reg1_val1[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 515.480 2100.000 516.080 ;
    END
  END reg1_val1[19]
  PIN reg1_val1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 466.520 2100.000 467.120 ;
    END
  END reg1_val1[1]
  PIN reg1_val1[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 518.200 2100.000 518.800 ;
    END
  END reg1_val1[20]
  PIN reg1_val1[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 520.920 2100.000 521.520 ;
    END
  END reg1_val1[21]
  PIN reg1_val1[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 523.640 2100.000 524.240 ;
    END
  END reg1_val1[22]
  PIN reg1_val1[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 526.360 2100.000 526.960 ;
    END
  END reg1_val1[23]
  PIN reg1_val1[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 529.080 2100.000 529.680 ;
    END
  END reg1_val1[24]
  PIN reg1_val1[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 531.800 2100.000 532.400 ;
    END
  END reg1_val1[25]
  PIN reg1_val1[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 534.520 2100.000 535.120 ;
    END
  END reg1_val1[26]
  PIN reg1_val1[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 537.240 2100.000 537.840 ;
    END
  END reg1_val1[27]
  PIN reg1_val1[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 539.960 2100.000 540.560 ;
    END
  END reg1_val1[28]
  PIN reg1_val1[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 542.680 2100.000 543.280 ;
    END
  END reg1_val1[29]
  PIN reg1_val1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 469.240 2100.000 469.840 ;
    END
  END reg1_val1[2]
  PIN reg1_val1[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 545.400 2100.000 546.000 ;
    END
  END reg1_val1[30]
  PIN reg1_val1[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 548.120 2100.000 548.720 ;
    END
  END reg1_val1[31]
  PIN reg1_val1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 471.960 2100.000 472.560 ;
    END
  END reg1_val1[3]
  PIN reg1_val1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 474.680 2100.000 475.280 ;
    END
  END reg1_val1[4]
  PIN reg1_val1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 477.400 2100.000 478.000 ;
    END
  END reg1_val1[5]
  PIN reg1_val1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 480.120 2100.000 480.720 ;
    END
  END reg1_val1[6]
  PIN reg1_val1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 482.840 2100.000 483.440 ;
    END
  END reg1_val1[7]
  PIN reg1_val1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 485.560 2100.000 486.160 ;
    END
  END reg1_val1[8]
  PIN reg1_val1[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 488.280 2100.000 488.880 ;
    END
  END reg1_val1[9]
  PIN reg1_val2[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 463.800 4.000 464.400 ;
    END
  END reg1_val2[0]
  PIN reg1_val2[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 491.000 4.000 491.600 ;
    END
  END reg1_val2[10]
  PIN reg1_val2[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 493.720 4.000 494.320 ;
    END
  END reg1_val2[11]
  PIN reg1_val2[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 496.440 4.000 497.040 ;
    END
  END reg1_val2[12]
  PIN reg1_val2[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 499.160 4.000 499.760 ;
    END
  END reg1_val2[13]
  PIN reg1_val2[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 501.880 4.000 502.480 ;
    END
  END reg1_val2[14]
  PIN reg1_val2[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 504.600 4.000 505.200 ;
    END
  END reg1_val2[15]
  PIN reg1_val2[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 507.320 4.000 507.920 ;
    END
  END reg1_val2[16]
  PIN reg1_val2[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 510.040 4.000 510.640 ;
    END
  END reg1_val2[17]
  PIN reg1_val2[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 512.760 4.000 513.360 ;
    END
  END reg1_val2[18]
  PIN reg1_val2[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 515.480 4.000 516.080 ;
    END
  END reg1_val2[19]
  PIN reg1_val2[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 466.520 4.000 467.120 ;
    END
  END reg1_val2[1]
  PIN reg1_val2[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 518.200 4.000 518.800 ;
    END
  END reg1_val2[20]
  PIN reg1_val2[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 520.920 4.000 521.520 ;
    END
  END reg1_val2[21]
  PIN reg1_val2[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 523.640 4.000 524.240 ;
    END
  END reg1_val2[22]
  PIN reg1_val2[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 526.360 4.000 526.960 ;
    END
  END reg1_val2[23]
  PIN reg1_val2[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 529.080 4.000 529.680 ;
    END
  END reg1_val2[24]
  PIN reg1_val2[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 531.800 4.000 532.400 ;
    END
  END reg1_val2[25]
  PIN reg1_val2[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 534.520 4.000 535.120 ;
    END
  END reg1_val2[26]
  PIN reg1_val2[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 537.240 4.000 537.840 ;
    END
  END reg1_val2[27]
  PIN reg1_val2[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 539.960 4.000 540.560 ;
    END
  END reg1_val2[28]
  PIN reg1_val2[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 542.680 4.000 543.280 ;
    END
  END reg1_val2[29]
  PIN reg1_val2[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 469.240 4.000 469.840 ;
    END
  END reg1_val2[2]
  PIN reg1_val2[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 545.400 4.000 546.000 ;
    END
  END reg1_val2[30]
  PIN reg1_val2[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 548.120 4.000 548.720 ;
    END
  END reg1_val2[31]
  PIN reg1_val2[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 471.960 4.000 472.560 ;
    END
  END reg1_val2[3]
  PIN reg1_val2[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 474.680 4.000 475.280 ;
    END
  END reg1_val2[4]
  PIN reg1_val2[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 477.400 4.000 478.000 ;
    END
  END reg1_val2[5]
  PIN reg1_val2[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 480.120 4.000 480.720 ;
    END
  END reg1_val2[6]
  PIN reg1_val2[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 482.840 4.000 483.440 ;
    END
  END reg1_val2[7]
  PIN reg1_val2[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 485.560 4.000 486.160 ;
    END
  END reg1_val2[8]
  PIN reg1_val2[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 488.280 4.000 488.880 ;
    END
  END reg1_val2[9]
  PIN reg2_idx0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.337000 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met2 ;
        RECT 287.130 636.000 287.410 640.000 ;
    END
  END reg2_idx0[0]
  PIN reg2_idx0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 294.950 636.000 295.230 640.000 ;
    END
  END reg2_idx0[1]
  PIN reg2_idx0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.189000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 302.770 636.000 303.050 640.000 ;
    END
  END reg2_idx0[2]
  PIN reg2_idx0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.383000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 310.590 636.000 310.870 640.000 ;
    END
  END reg2_idx0[3]
  PIN reg2_idx0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.293000 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met2 ;
        RECT 318.410 636.000 318.690 640.000 ;
    END
  END reg2_idx0[4]
  PIN reg2_idx1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.842000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 15.000 2100.000 15.600 ;
    END
  END reg2_idx1[0]
  PIN reg2_idx1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.594500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 17.720 2100.000 18.320 ;
    END
  END reg2_idx1[1]
  PIN reg2_idx1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.327000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 20.440 2100.000 21.040 ;
    END
  END reg2_idx1[2]
  PIN reg2_idx1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.980000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 23.160 2100.000 23.760 ;
    END
  END reg2_idx1[3]
  PIN reg2_idx1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.980000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 25.880 2100.000 26.480 ;
    END
  END reg2_idx1[4]
  PIN reg2_idx2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.000 4.000 15.600 ;
    END
  END reg2_idx2[0]
  PIN reg2_idx2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.594500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.720 4.000 18.320 ;
    END
  END reg2_idx2[1]
  PIN reg2_idx2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.041000 ;
    ANTENNADIFFAREA 2.173500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END reg2_idx2[2]
  PIN reg2_idx2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.383000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.160 4.000 23.760 ;
    END
  END reg2_idx2[3]
  PIN reg2_idx2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.293000 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 4.000 26.480 ;
    END
  END reg2_idx2[4]
  PIN reg2_val0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1827.670 636.000 1827.950 640.000 ;
    END
  END reg2_val0[0]
  PIN reg2_val0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1905.870 636.000 1906.150 640.000 ;
    END
  END reg2_val0[10]
  PIN reg2_val0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1913.690 636.000 1913.970 640.000 ;
    END
  END reg2_val0[11]
  PIN reg2_val0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1921.510 636.000 1921.790 640.000 ;
    END
  END reg2_val0[12]
  PIN reg2_val0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1929.330 636.000 1929.610 640.000 ;
    END
  END reg2_val0[13]
  PIN reg2_val0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1937.150 636.000 1937.430 640.000 ;
    END
  END reg2_val0[14]
  PIN reg2_val0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1944.970 636.000 1945.250 640.000 ;
    END
  END reg2_val0[15]
  PIN reg2_val0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1952.790 636.000 1953.070 640.000 ;
    END
  END reg2_val0[16]
  PIN reg2_val0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1960.610 636.000 1960.890 640.000 ;
    END
  END reg2_val0[17]
  PIN reg2_val0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1968.430 636.000 1968.710 640.000 ;
    END
  END reg2_val0[18]
  PIN reg2_val0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1976.250 636.000 1976.530 640.000 ;
    END
  END reg2_val0[19]
  PIN reg2_val0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1835.490 636.000 1835.770 640.000 ;
    END
  END reg2_val0[1]
  PIN reg2_val0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1984.070 636.000 1984.350 640.000 ;
    END
  END reg2_val0[20]
  PIN reg2_val0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1991.890 636.000 1992.170 640.000 ;
    END
  END reg2_val0[21]
  PIN reg2_val0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1999.710 636.000 1999.990 640.000 ;
    END
  END reg2_val0[22]
  PIN reg2_val0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 2007.530 636.000 2007.810 640.000 ;
    END
  END reg2_val0[23]
  PIN reg2_val0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 2015.350 636.000 2015.630 640.000 ;
    END
  END reg2_val0[24]
  PIN reg2_val0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 2023.170 636.000 2023.450 640.000 ;
    END
  END reg2_val0[25]
  PIN reg2_val0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 2030.990 636.000 2031.270 640.000 ;
    END
  END reg2_val0[26]
  PIN reg2_val0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 2038.810 636.000 2039.090 640.000 ;
    END
  END reg2_val0[27]
  PIN reg2_val0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met2 ;
        RECT 2046.630 636.000 2046.910 640.000 ;
    END
  END reg2_val0[28]
  PIN reg2_val0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 2054.450 636.000 2054.730 640.000 ;
    END
  END reg2_val0[29]
  PIN reg2_val0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1843.310 636.000 1843.590 640.000 ;
    END
  END reg2_val0[2]
  PIN reg2_val0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met2 ;
        RECT 2062.270 636.000 2062.550 640.000 ;
    END
  END reg2_val0[30]
  PIN reg2_val0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met2 ;
        RECT 2070.090 636.000 2070.370 640.000 ;
    END
  END reg2_val0[31]
  PIN reg2_val0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1851.130 636.000 1851.410 640.000 ;
    END
  END reg2_val0[3]
  PIN reg2_val0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1858.950 636.000 1859.230 640.000 ;
    END
  END reg2_val0[4]
  PIN reg2_val0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1866.770 636.000 1867.050 640.000 ;
    END
  END reg2_val0[5]
  PIN reg2_val0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1874.590 636.000 1874.870 640.000 ;
    END
  END reg2_val0[6]
  PIN reg2_val0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1882.410 636.000 1882.690 640.000 ;
    END
  END reg2_val0[7]
  PIN reg2_val0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1890.230 636.000 1890.510 640.000 ;
    END
  END reg2_val0[8]
  PIN reg2_val0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1898.050 636.000 1898.330 640.000 ;
    END
  END reg2_val0[9]
  PIN reg2_val1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 550.840 2100.000 551.440 ;
    END
  END reg2_val1[0]
  PIN reg2_val1[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 578.040 2100.000 578.640 ;
    END
  END reg2_val1[10]
  PIN reg2_val1[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 580.760 2100.000 581.360 ;
    END
  END reg2_val1[11]
  PIN reg2_val1[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 583.480 2100.000 584.080 ;
    END
  END reg2_val1[12]
  PIN reg2_val1[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 586.200 2100.000 586.800 ;
    END
  END reg2_val1[13]
  PIN reg2_val1[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 588.920 2100.000 589.520 ;
    END
  END reg2_val1[14]
  PIN reg2_val1[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 591.640 2100.000 592.240 ;
    END
  END reg2_val1[15]
  PIN reg2_val1[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 594.360 2100.000 594.960 ;
    END
  END reg2_val1[16]
  PIN reg2_val1[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 597.080 2100.000 597.680 ;
    END
  END reg2_val1[17]
  PIN reg2_val1[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 599.800 2100.000 600.400 ;
    END
  END reg2_val1[18]
  PIN reg2_val1[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 602.520 2100.000 603.120 ;
    END
  END reg2_val1[19]
  PIN reg2_val1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 553.560 2100.000 554.160 ;
    END
  END reg2_val1[1]
  PIN reg2_val1[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 605.240 2100.000 605.840 ;
    END
  END reg2_val1[20]
  PIN reg2_val1[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 607.960 2100.000 608.560 ;
    END
  END reg2_val1[21]
  PIN reg2_val1[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 610.680 2100.000 611.280 ;
    END
  END reg2_val1[22]
  PIN reg2_val1[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 613.400 2100.000 614.000 ;
    END
  END reg2_val1[23]
  PIN reg2_val1[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 616.120 2100.000 616.720 ;
    END
  END reg2_val1[24]
  PIN reg2_val1[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 618.840 2100.000 619.440 ;
    END
  END reg2_val1[25]
  PIN reg2_val1[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 621.560 2100.000 622.160 ;
    END
  END reg2_val1[26]
  PIN reg2_val1[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 624.280 2100.000 624.880 ;
    END
  END reg2_val1[27]
  PIN reg2_val1[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 627.000 2100.000 627.600 ;
    END
  END reg2_val1[28]
  PIN reg2_val1[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 629.720 2100.000 630.320 ;
    END
  END reg2_val1[29]
  PIN reg2_val1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 556.280 2100.000 556.880 ;
    END
  END reg2_val1[2]
  PIN reg2_val1[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 632.440 2100.000 633.040 ;
    END
  END reg2_val1[30]
  PIN reg2_val1[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 635.160 2100.000 635.760 ;
    END
  END reg2_val1[31]
  PIN reg2_val1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 559.000 2100.000 559.600 ;
    END
  END reg2_val1[3]
  PIN reg2_val1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 561.720 2100.000 562.320 ;
    END
  END reg2_val1[4]
  PIN reg2_val1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 564.440 2100.000 565.040 ;
    END
  END reg2_val1[5]
  PIN reg2_val1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 567.160 2100.000 567.760 ;
    END
  END reg2_val1[6]
  PIN reg2_val1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 569.880 2100.000 570.480 ;
    END
  END reg2_val1[7]
  PIN reg2_val1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 572.600 2100.000 573.200 ;
    END
  END reg2_val1[8]
  PIN reg2_val1[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 575.320 2100.000 575.920 ;
    END
  END reg2_val1[9]
  PIN reg2_val2[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 550.840 4.000 551.440 ;
    END
  END reg2_val2[0]
  PIN reg2_val2[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 578.040 4.000 578.640 ;
    END
  END reg2_val2[10]
  PIN reg2_val2[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 580.760 4.000 581.360 ;
    END
  END reg2_val2[11]
  PIN reg2_val2[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 583.480 4.000 584.080 ;
    END
  END reg2_val2[12]
  PIN reg2_val2[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 586.200 4.000 586.800 ;
    END
  END reg2_val2[13]
  PIN reg2_val2[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 588.920 4.000 589.520 ;
    END
  END reg2_val2[14]
  PIN reg2_val2[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 591.640 4.000 592.240 ;
    END
  END reg2_val2[15]
  PIN reg2_val2[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 594.360 4.000 594.960 ;
    END
  END reg2_val2[16]
  PIN reg2_val2[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 597.080 4.000 597.680 ;
    END
  END reg2_val2[17]
  PIN reg2_val2[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 599.800 4.000 600.400 ;
    END
  END reg2_val2[18]
  PIN reg2_val2[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 602.520 4.000 603.120 ;
    END
  END reg2_val2[19]
  PIN reg2_val2[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 553.560 4.000 554.160 ;
    END
  END reg2_val2[1]
  PIN reg2_val2[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 605.240 4.000 605.840 ;
    END
  END reg2_val2[20]
  PIN reg2_val2[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 607.960 4.000 608.560 ;
    END
  END reg2_val2[21]
  PIN reg2_val2[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 610.680 4.000 611.280 ;
    END
  END reg2_val2[22]
  PIN reg2_val2[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 613.400 4.000 614.000 ;
    END
  END reg2_val2[23]
  PIN reg2_val2[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 616.120 4.000 616.720 ;
    END
  END reg2_val2[24]
  PIN reg2_val2[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 618.840 4.000 619.440 ;
    END
  END reg2_val2[25]
  PIN reg2_val2[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 621.560 4.000 622.160 ;
    END
  END reg2_val2[26]
  PIN reg2_val2[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 624.280 4.000 624.880 ;
    END
  END reg2_val2[27]
  PIN reg2_val2[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 627.000 4.000 627.600 ;
    END
  END reg2_val2[28]
  PIN reg2_val2[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 629.720 4.000 630.320 ;
    END
  END reg2_val2[29]
  PIN reg2_val2[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 556.280 4.000 556.880 ;
    END
  END reg2_val2[2]
  PIN reg2_val2[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 632.440 4.000 633.040 ;
    END
  END reg2_val2[30]
  PIN reg2_val2[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 635.160 4.000 635.760 ;
    END
  END reg2_val2[31]
  PIN reg2_val2[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 559.000 4.000 559.600 ;
    END
  END reg2_val2[3]
  PIN reg2_val2[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 561.720 4.000 562.320 ;
    END
  END reg2_val2[4]
  PIN reg2_val2[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 564.440 4.000 565.040 ;
    END
  END reg2_val2[5]
  PIN reg2_val2[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 567.160 4.000 567.760 ;
    END
  END reg2_val2[6]
  PIN reg2_val2[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 569.880 4.000 570.480 ;
    END
  END reg2_val2[7]
  PIN reg2_val2[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 572.600 4.000 573.200 ;
    END
  END reg2_val2[8]
  PIN reg2_val2[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 575.320 4.000 575.920 ;
    END
  END reg2_val2[9]
  PIN rst_eu
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.862000 ;
    PORT
      LAYER met2 ;
        RECT 21.250 636.000 21.530 640.000 ;
    END
  END rst_eu
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.499500 ;
    PORT
      LAYER met2 ;
        RECT 1982.690 0.000 1982.970 4.000 ;
    END
  END rst_n
  PIN sign_extend0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 951.830 636.000 952.110 640.000 ;
    END
  END sign_extend0
  PIN sign_extend1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 246.200 2100.000 246.800 ;
    END
  END sign_extend1
  PIN sign_extend2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 246.200 4.000 246.800 ;
    END
  END sign_extend2
  PIN take_branch0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.160000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1014.390 636.000 1014.670 640.000 ;
    END
  END take_branch0
  PIN take_branch1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.081500 ;
    PORT
      LAYER met3 ;
        RECT 2096.000 267.960 2100.000 268.560 ;
    END
  END take_branch1
  PIN take_branch2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 267.960 4.000 268.560 ;
    END
  END take_branch2
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 628.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 628.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 628.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 628.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 628.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 628.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 628.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 628.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 628.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 628.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.040 10.640 1558.640 628.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1710.640 10.640 1712.240 628.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1864.240 10.640 1865.840 628.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 2017.840 10.640 2019.440 628.560 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 628.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 628.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 628.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 628.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 628.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 628.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 628.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 628.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 628.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 628.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1633.840 10.640 1635.440 628.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1787.440 10.640 1789.040 628.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 1941.040 10.640 1942.640 628.560 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1964.750 0.000 1965.030 4.000 ;
    END
  END wb_clk_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2094.380 628.405 ;
      LAYER met1 ;
        RECT 5.520 6.160 2094.380 639.840 ;
      LAYER met2 ;
        RECT 12.050 635.720 20.970 639.870 ;
        RECT 21.810 635.720 28.790 639.870 ;
        RECT 29.630 635.720 36.610 639.870 ;
        RECT 37.450 635.720 44.430 639.870 ;
        RECT 45.270 635.720 52.250 639.870 ;
        RECT 53.090 635.720 60.070 639.870 ;
        RECT 60.910 635.720 67.890 639.870 ;
        RECT 68.730 635.720 75.710 639.870 ;
        RECT 76.550 635.720 83.530 639.870 ;
        RECT 84.370 635.720 91.350 639.870 ;
        RECT 92.190 635.720 99.170 639.870 ;
        RECT 100.010 635.720 106.990 639.870 ;
        RECT 107.830 635.720 114.810 639.870 ;
        RECT 115.650 635.720 122.630 639.870 ;
        RECT 123.470 635.720 130.450 639.870 ;
        RECT 131.290 635.720 138.270 639.870 ;
        RECT 139.110 635.720 146.090 639.870 ;
        RECT 146.930 635.720 153.910 639.870 ;
        RECT 154.750 635.720 161.730 639.870 ;
        RECT 162.570 635.720 169.550 639.870 ;
        RECT 170.390 635.720 177.370 639.870 ;
        RECT 178.210 635.720 185.190 639.870 ;
        RECT 186.030 635.720 193.010 639.870 ;
        RECT 193.850 635.720 200.830 639.870 ;
        RECT 201.670 635.720 208.650 639.870 ;
        RECT 209.490 635.720 216.470 639.870 ;
        RECT 217.310 635.720 224.290 639.870 ;
        RECT 225.130 635.720 232.110 639.870 ;
        RECT 232.950 635.720 239.930 639.870 ;
        RECT 240.770 635.720 247.750 639.870 ;
        RECT 248.590 635.720 255.570 639.870 ;
        RECT 256.410 635.720 263.390 639.870 ;
        RECT 264.230 635.720 271.210 639.870 ;
        RECT 272.050 635.720 279.030 639.870 ;
        RECT 279.870 635.720 286.850 639.870 ;
        RECT 287.690 635.720 294.670 639.870 ;
        RECT 295.510 635.720 302.490 639.870 ;
        RECT 303.330 635.720 310.310 639.870 ;
        RECT 311.150 635.720 318.130 639.870 ;
        RECT 318.970 635.720 325.950 639.870 ;
        RECT 326.790 635.720 333.770 639.870 ;
        RECT 334.610 635.720 341.590 639.870 ;
        RECT 342.430 635.720 349.410 639.870 ;
        RECT 350.250 635.720 357.230 639.870 ;
        RECT 358.070 635.720 365.050 639.870 ;
        RECT 365.890 635.720 372.870 639.870 ;
        RECT 373.710 635.720 380.690 639.870 ;
        RECT 381.530 635.720 388.510 639.870 ;
        RECT 389.350 635.720 396.330 639.870 ;
        RECT 397.170 635.720 404.150 639.870 ;
        RECT 404.990 635.720 411.970 639.870 ;
        RECT 412.810 635.720 419.790 639.870 ;
        RECT 420.630 635.720 427.610 639.870 ;
        RECT 428.450 635.720 435.430 639.870 ;
        RECT 436.270 635.720 443.250 639.870 ;
        RECT 444.090 635.720 451.070 639.870 ;
        RECT 451.910 635.720 458.890 639.870 ;
        RECT 459.730 635.720 466.710 639.870 ;
        RECT 467.550 635.720 474.530 639.870 ;
        RECT 475.370 635.720 482.350 639.870 ;
        RECT 483.190 635.720 490.170 639.870 ;
        RECT 491.010 635.720 497.990 639.870 ;
        RECT 498.830 635.720 505.810 639.870 ;
        RECT 506.650 635.720 513.630 639.870 ;
        RECT 514.470 635.720 521.450 639.870 ;
        RECT 522.290 635.720 529.270 639.870 ;
        RECT 530.110 635.720 537.090 639.870 ;
        RECT 537.930 635.720 544.910 639.870 ;
        RECT 545.750 635.720 552.730 639.870 ;
        RECT 553.570 635.720 560.550 639.870 ;
        RECT 561.390 635.720 568.370 639.870 ;
        RECT 569.210 635.720 576.190 639.870 ;
        RECT 577.030 635.720 584.010 639.870 ;
        RECT 584.850 635.720 591.830 639.870 ;
        RECT 592.670 635.720 599.650 639.870 ;
        RECT 600.490 635.720 607.470 639.870 ;
        RECT 608.310 635.720 615.290 639.870 ;
        RECT 616.130 635.720 623.110 639.870 ;
        RECT 623.950 635.720 630.930 639.870 ;
        RECT 631.770 635.720 638.750 639.870 ;
        RECT 639.590 635.720 646.570 639.870 ;
        RECT 647.410 635.720 654.390 639.870 ;
        RECT 655.230 635.720 662.210 639.870 ;
        RECT 663.050 635.720 670.030 639.870 ;
        RECT 670.870 635.720 677.850 639.870 ;
        RECT 678.690 635.720 685.670 639.870 ;
        RECT 686.510 635.720 693.490 639.870 ;
        RECT 694.330 635.720 701.310 639.870 ;
        RECT 702.150 635.720 709.130 639.870 ;
        RECT 709.970 635.720 716.950 639.870 ;
        RECT 717.790 635.720 724.770 639.870 ;
        RECT 725.610 635.720 732.590 639.870 ;
        RECT 733.430 635.720 740.410 639.870 ;
        RECT 741.250 635.720 748.230 639.870 ;
        RECT 749.070 635.720 756.050 639.870 ;
        RECT 756.890 635.720 763.870 639.870 ;
        RECT 764.710 635.720 771.690 639.870 ;
        RECT 772.530 635.720 779.510 639.870 ;
        RECT 780.350 635.720 787.330 639.870 ;
        RECT 788.170 635.720 795.150 639.870 ;
        RECT 795.990 635.720 802.970 639.870 ;
        RECT 803.810 635.720 810.790 639.870 ;
        RECT 811.630 635.720 818.610 639.870 ;
        RECT 819.450 635.720 826.430 639.870 ;
        RECT 827.270 635.720 834.250 639.870 ;
        RECT 835.090 635.720 842.070 639.870 ;
        RECT 842.910 635.720 849.890 639.870 ;
        RECT 850.730 635.720 857.710 639.870 ;
        RECT 858.550 635.720 865.530 639.870 ;
        RECT 866.370 635.720 873.350 639.870 ;
        RECT 874.190 635.720 881.170 639.870 ;
        RECT 882.010 635.720 888.990 639.870 ;
        RECT 889.830 635.720 896.810 639.870 ;
        RECT 897.650 635.720 904.630 639.870 ;
        RECT 905.470 635.720 912.450 639.870 ;
        RECT 913.290 635.720 920.270 639.870 ;
        RECT 921.110 635.720 928.090 639.870 ;
        RECT 928.930 635.720 935.910 639.870 ;
        RECT 936.750 635.720 943.730 639.870 ;
        RECT 944.570 635.720 951.550 639.870 ;
        RECT 952.390 635.720 959.370 639.870 ;
        RECT 960.210 635.720 967.190 639.870 ;
        RECT 968.030 635.720 975.010 639.870 ;
        RECT 975.850 635.720 982.830 639.870 ;
        RECT 983.670 635.720 990.650 639.870 ;
        RECT 991.490 635.720 998.470 639.870 ;
        RECT 999.310 635.720 1006.290 639.870 ;
        RECT 1007.130 635.720 1014.110 639.870 ;
        RECT 1014.950 635.720 1021.930 639.870 ;
        RECT 1022.770 635.720 1029.750 639.870 ;
        RECT 1030.590 635.720 1037.570 639.870 ;
        RECT 1038.410 635.720 1045.390 639.870 ;
        RECT 1046.230 635.720 1053.210 639.870 ;
        RECT 1054.050 635.720 1061.030 639.870 ;
        RECT 1061.870 635.720 1068.850 639.870 ;
        RECT 1069.690 635.720 1076.670 639.870 ;
        RECT 1077.510 635.720 1084.490 639.870 ;
        RECT 1085.330 635.720 1092.310 639.870 ;
        RECT 1093.150 635.720 1100.130 639.870 ;
        RECT 1100.970 635.720 1107.950 639.870 ;
        RECT 1108.790 635.720 1115.770 639.870 ;
        RECT 1116.610 635.720 1123.590 639.870 ;
        RECT 1124.430 635.720 1131.410 639.870 ;
        RECT 1132.250 635.720 1139.230 639.870 ;
        RECT 1140.070 635.720 1147.050 639.870 ;
        RECT 1147.890 635.720 1154.870 639.870 ;
        RECT 1155.710 635.720 1162.690 639.870 ;
        RECT 1163.530 635.720 1170.510 639.870 ;
        RECT 1171.350 635.720 1178.330 639.870 ;
        RECT 1179.170 635.720 1186.150 639.870 ;
        RECT 1186.990 635.720 1193.970 639.870 ;
        RECT 1194.810 635.720 1201.790 639.870 ;
        RECT 1202.630 635.720 1209.610 639.870 ;
        RECT 1210.450 635.720 1217.430 639.870 ;
        RECT 1218.270 635.720 1225.250 639.870 ;
        RECT 1226.090 635.720 1233.070 639.870 ;
        RECT 1233.910 635.720 1240.890 639.870 ;
        RECT 1241.730 635.720 1248.710 639.870 ;
        RECT 1249.550 635.720 1256.530 639.870 ;
        RECT 1257.370 635.720 1264.350 639.870 ;
        RECT 1265.190 635.720 1272.170 639.870 ;
        RECT 1273.010 635.720 1279.990 639.870 ;
        RECT 1280.830 635.720 1287.810 639.870 ;
        RECT 1288.650 635.720 1295.630 639.870 ;
        RECT 1296.470 635.720 1303.450 639.870 ;
        RECT 1304.290 635.720 1311.270 639.870 ;
        RECT 1312.110 635.720 1319.090 639.870 ;
        RECT 1319.930 635.720 1326.910 639.870 ;
        RECT 1327.750 635.720 1334.730 639.870 ;
        RECT 1335.570 635.720 1342.550 639.870 ;
        RECT 1343.390 635.720 1350.370 639.870 ;
        RECT 1351.210 635.720 1358.190 639.870 ;
        RECT 1359.030 635.720 1366.010 639.870 ;
        RECT 1366.850 635.720 1373.830 639.870 ;
        RECT 1374.670 635.720 1381.650 639.870 ;
        RECT 1382.490 635.720 1389.470 639.870 ;
        RECT 1390.310 635.720 1397.290 639.870 ;
        RECT 1398.130 635.720 1405.110 639.870 ;
        RECT 1405.950 635.720 1412.930 639.870 ;
        RECT 1413.770 635.720 1420.750 639.870 ;
        RECT 1421.590 635.720 1428.570 639.870 ;
        RECT 1429.410 635.720 1436.390 639.870 ;
        RECT 1437.230 635.720 1444.210 639.870 ;
        RECT 1445.050 635.720 1452.030 639.870 ;
        RECT 1452.870 635.720 1459.850 639.870 ;
        RECT 1460.690 635.720 1467.670 639.870 ;
        RECT 1468.510 635.720 1475.490 639.870 ;
        RECT 1476.330 635.720 1483.310 639.870 ;
        RECT 1484.150 635.720 1491.130 639.870 ;
        RECT 1491.970 635.720 1498.950 639.870 ;
        RECT 1499.790 635.720 1506.770 639.870 ;
        RECT 1507.610 635.720 1514.590 639.870 ;
        RECT 1515.430 635.720 1522.410 639.870 ;
        RECT 1523.250 635.720 1530.230 639.870 ;
        RECT 1531.070 635.720 1538.050 639.870 ;
        RECT 1538.890 635.720 1545.870 639.870 ;
        RECT 1546.710 635.720 1553.690 639.870 ;
        RECT 1554.530 635.720 1561.510 639.870 ;
        RECT 1562.350 635.720 1569.330 639.870 ;
        RECT 1570.170 635.720 1577.150 639.870 ;
        RECT 1577.990 635.720 1584.970 639.870 ;
        RECT 1585.810 635.720 1592.790 639.870 ;
        RECT 1593.630 635.720 1600.610 639.870 ;
        RECT 1601.450 635.720 1608.430 639.870 ;
        RECT 1609.270 635.720 1616.250 639.870 ;
        RECT 1617.090 635.720 1624.070 639.870 ;
        RECT 1624.910 635.720 1631.890 639.870 ;
        RECT 1632.730 635.720 1639.710 639.870 ;
        RECT 1640.550 635.720 1647.530 639.870 ;
        RECT 1648.370 635.720 1655.350 639.870 ;
        RECT 1656.190 635.720 1663.170 639.870 ;
        RECT 1664.010 635.720 1670.990 639.870 ;
        RECT 1671.830 635.720 1678.810 639.870 ;
        RECT 1679.650 635.720 1686.630 639.870 ;
        RECT 1687.470 635.720 1694.450 639.870 ;
        RECT 1695.290 635.720 1702.270 639.870 ;
        RECT 1703.110 635.720 1710.090 639.870 ;
        RECT 1710.930 635.720 1717.910 639.870 ;
        RECT 1718.750 635.720 1725.730 639.870 ;
        RECT 1726.570 635.720 1733.550 639.870 ;
        RECT 1734.390 635.720 1741.370 639.870 ;
        RECT 1742.210 635.720 1749.190 639.870 ;
        RECT 1750.030 635.720 1757.010 639.870 ;
        RECT 1757.850 635.720 1764.830 639.870 ;
        RECT 1765.670 635.720 1772.650 639.870 ;
        RECT 1773.490 635.720 1780.470 639.870 ;
        RECT 1781.310 635.720 1788.290 639.870 ;
        RECT 1789.130 635.720 1796.110 639.870 ;
        RECT 1796.950 635.720 1803.930 639.870 ;
        RECT 1804.770 635.720 1811.750 639.870 ;
        RECT 1812.590 635.720 1819.570 639.870 ;
        RECT 1820.410 635.720 1827.390 639.870 ;
        RECT 1828.230 635.720 1835.210 639.870 ;
        RECT 1836.050 635.720 1843.030 639.870 ;
        RECT 1843.870 635.720 1850.850 639.870 ;
        RECT 1851.690 635.720 1858.670 639.870 ;
        RECT 1859.510 635.720 1866.490 639.870 ;
        RECT 1867.330 635.720 1874.310 639.870 ;
        RECT 1875.150 635.720 1882.130 639.870 ;
        RECT 1882.970 635.720 1889.950 639.870 ;
        RECT 1890.790 635.720 1897.770 639.870 ;
        RECT 1898.610 635.720 1905.590 639.870 ;
        RECT 1906.430 635.720 1913.410 639.870 ;
        RECT 1914.250 635.720 1921.230 639.870 ;
        RECT 1922.070 635.720 1929.050 639.870 ;
        RECT 1929.890 635.720 1936.870 639.870 ;
        RECT 1937.710 635.720 1944.690 639.870 ;
        RECT 1945.530 635.720 1952.510 639.870 ;
        RECT 1953.350 635.720 1960.330 639.870 ;
        RECT 1961.170 635.720 1968.150 639.870 ;
        RECT 1968.990 635.720 1975.970 639.870 ;
        RECT 1976.810 635.720 1983.790 639.870 ;
        RECT 1984.630 635.720 1991.610 639.870 ;
        RECT 1992.450 635.720 1999.430 639.870 ;
        RECT 2000.270 635.720 2007.250 639.870 ;
        RECT 2008.090 635.720 2015.070 639.870 ;
        RECT 2015.910 635.720 2022.890 639.870 ;
        RECT 2023.730 635.720 2030.710 639.870 ;
        RECT 2031.550 635.720 2038.530 639.870 ;
        RECT 2039.370 635.720 2046.350 639.870 ;
        RECT 2047.190 635.720 2054.170 639.870 ;
        RECT 2055.010 635.720 2061.990 639.870 ;
        RECT 2062.830 635.720 2069.810 639.870 ;
        RECT 2070.650 635.720 2077.630 639.870 ;
        RECT 2078.470 635.720 2091.990 639.870 ;
        RECT 12.050 4.280 2091.990 635.720 ;
        RECT 12.050 1.515 26.950 4.280 ;
        RECT 27.790 1.515 44.890 4.280 ;
        RECT 45.730 1.515 62.830 4.280 ;
        RECT 63.670 1.515 80.770 4.280 ;
        RECT 81.610 1.515 98.710 4.280 ;
        RECT 99.550 1.515 116.650 4.280 ;
        RECT 117.490 1.515 134.590 4.280 ;
        RECT 135.430 1.515 152.530 4.280 ;
        RECT 153.370 1.515 170.470 4.280 ;
        RECT 171.310 1.515 188.410 4.280 ;
        RECT 189.250 1.515 206.350 4.280 ;
        RECT 207.190 1.515 224.290 4.280 ;
        RECT 225.130 1.515 242.230 4.280 ;
        RECT 243.070 1.515 260.170 4.280 ;
        RECT 261.010 1.515 278.110 4.280 ;
        RECT 278.950 1.515 296.050 4.280 ;
        RECT 296.890 1.515 313.990 4.280 ;
        RECT 314.830 1.515 331.930 4.280 ;
        RECT 332.770 1.515 349.870 4.280 ;
        RECT 350.710 1.515 367.810 4.280 ;
        RECT 368.650 1.515 385.750 4.280 ;
        RECT 386.590 1.515 403.690 4.280 ;
        RECT 404.530 1.515 421.630 4.280 ;
        RECT 422.470 1.515 439.570 4.280 ;
        RECT 440.410 1.515 457.510 4.280 ;
        RECT 458.350 1.515 475.450 4.280 ;
        RECT 476.290 1.515 493.390 4.280 ;
        RECT 494.230 1.515 511.330 4.280 ;
        RECT 512.170 1.515 529.270 4.280 ;
        RECT 530.110 1.515 547.210 4.280 ;
        RECT 548.050 1.515 565.150 4.280 ;
        RECT 565.990 1.515 583.090 4.280 ;
        RECT 583.930 1.515 601.030 4.280 ;
        RECT 601.870 1.515 618.970 4.280 ;
        RECT 619.810 1.515 636.910 4.280 ;
        RECT 637.750 1.515 654.850 4.280 ;
        RECT 655.690 1.515 672.790 4.280 ;
        RECT 673.630 1.515 690.730 4.280 ;
        RECT 691.570 1.515 708.670 4.280 ;
        RECT 709.510 1.515 726.610 4.280 ;
        RECT 727.450 1.515 744.550 4.280 ;
        RECT 745.390 1.515 762.490 4.280 ;
        RECT 763.330 1.515 780.430 4.280 ;
        RECT 781.270 1.515 798.370 4.280 ;
        RECT 799.210 1.515 816.310 4.280 ;
        RECT 817.150 1.515 834.250 4.280 ;
        RECT 835.090 1.515 852.190 4.280 ;
        RECT 853.030 1.515 870.130 4.280 ;
        RECT 870.970 1.515 888.070 4.280 ;
        RECT 888.910 1.515 906.010 4.280 ;
        RECT 906.850 1.515 923.950 4.280 ;
        RECT 924.790 1.515 941.890 4.280 ;
        RECT 942.730 1.515 959.830 4.280 ;
        RECT 960.670 1.515 977.770 4.280 ;
        RECT 978.610 1.515 995.710 4.280 ;
        RECT 996.550 1.515 1013.650 4.280 ;
        RECT 1014.490 1.515 1031.590 4.280 ;
        RECT 1032.430 1.515 1049.530 4.280 ;
        RECT 1050.370 1.515 1067.470 4.280 ;
        RECT 1068.310 1.515 1085.410 4.280 ;
        RECT 1086.250 1.515 1103.350 4.280 ;
        RECT 1104.190 1.515 1121.290 4.280 ;
        RECT 1122.130 1.515 1139.230 4.280 ;
        RECT 1140.070 1.515 1157.170 4.280 ;
        RECT 1158.010 1.515 1175.110 4.280 ;
        RECT 1175.950 1.515 1193.050 4.280 ;
        RECT 1193.890 1.515 1210.990 4.280 ;
        RECT 1211.830 1.515 1228.930 4.280 ;
        RECT 1229.770 1.515 1246.870 4.280 ;
        RECT 1247.710 1.515 1264.810 4.280 ;
        RECT 1265.650 1.515 1282.750 4.280 ;
        RECT 1283.590 1.515 1300.690 4.280 ;
        RECT 1301.530 1.515 1318.630 4.280 ;
        RECT 1319.470 1.515 1336.570 4.280 ;
        RECT 1337.410 1.515 1354.510 4.280 ;
        RECT 1355.350 1.515 1372.450 4.280 ;
        RECT 1373.290 1.515 1390.390 4.280 ;
        RECT 1391.230 1.515 1408.330 4.280 ;
        RECT 1409.170 1.515 1426.270 4.280 ;
        RECT 1427.110 1.515 1444.210 4.280 ;
        RECT 1445.050 1.515 1462.150 4.280 ;
        RECT 1462.990 1.515 1480.090 4.280 ;
        RECT 1480.930 1.515 1498.030 4.280 ;
        RECT 1498.870 1.515 1515.970 4.280 ;
        RECT 1516.810 1.515 1533.910 4.280 ;
        RECT 1534.750 1.515 1551.850 4.280 ;
        RECT 1552.690 1.515 1569.790 4.280 ;
        RECT 1570.630 1.515 1587.730 4.280 ;
        RECT 1588.570 1.515 1605.670 4.280 ;
        RECT 1606.510 1.515 1623.610 4.280 ;
        RECT 1624.450 1.515 1641.550 4.280 ;
        RECT 1642.390 1.515 1659.490 4.280 ;
        RECT 1660.330 1.515 1677.430 4.280 ;
        RECT 1678.270 1.515 1695.370 4.280 ;
        RECT 1696.210 1.515 1713.310 4.280 ;
        RECT 1714.150 1.515 1731.250 4.280 ;
        RECT 1732.090 1.515 1749.190 4.280 ;
        RECT 1750.030 1.515 1767.130 4.280 ;
        RECT 1767.970 1.515 1785.070 4.280 ;
        RECT 1785.910 1.515 1803.010 4.280 ;
        RECT 1803.850 1.515 1820.950 4.280 ;
        RECT 1821.790 1.515 1838.890 4.280 ;
        RECT 1839.730 1.515 1856.830 4.280 ;
        RECT 1857.670 1.515 1874.770 4.280 ;
        RECT 1875.610 1.515 1892.710 4.280 ;
        RECT 1893.550 1.515 1910.650 4.280 ;
        RECT 1911.490 1.515 1928.590 4.280 ;
        RECT 1929.430 1.515 1946.530 4.280 ;
        RECT 1947.370 1.515 1964.470 4.280 ;
        RECT 1965.310 1.515 1982.410 4.280 ;
        RECT 1983.250 1.515 2000.350 4.280 ;
        RECT 2001.190 1.515 2018.290 4.280 ;
        RECT 2019.130 1.515 2036.230 4.280 ;
        RECT 2037.070 1.515 2054.170 4.280 ;
        RECT 2055.010 1.515 2072.110 4.280 ;
        RECT 2072.950 1.515 2091.990 4.280 ;
      LAYER met3 ;
        RECT 4.400 637.480 2095.600 638.345 ;
        RECT 4.000 636.160 2096.000 637.480 ;
        RECT 4.400 634.760 2095.600 636.160 ;
        RECT 4.000 633.440 2096.000 634.760 ;
        RECT 4.400 632.040 2095.600 633.440 ;
        RECT 4.000 630.720 2096.000 632.040 ;
        RECT 4.400 629.320 2095.600 630.720 ;
        RECT 4.000 628.000 2096.000 629.320 ;
        RECT 4.400 626.600 2095.600 628.000 ;
        RECT 4.000 625.280 2096.000 626.600 ;
        RECT 4.400 623.880 2095.600 625.280 ;
        RECT 4.000 622.560 2096.000 623.880 ;
        RECT 4.400 621.160 2095.600 622.560 ;
        RECT 4.000 619.840 2096.000 621.160 ;
        RECT 4.400 618.440 2095.600 619.840 ;
        RECT 4.000 617.120 2096.000 618.440 ;
        RECT 4.400 615.720 2095.600 617.120 ;
        RECT 4.000 614.400 2096.000 615.720 ;
        RECT 4.400 613.000 2095.600 614.400 ;
        RECT 4.000 611.680 2096.000 613.000 ;
        RECT 4.400 610.280 2095.600 611.680 ;
        RECT 4.000 608.960 2096.000 610.280 ;
        RECT 4.400 607.560 2095.600 608.960 ;
        RECT 4.000 606.240 2096.000 607.560 ;
        RECT 4.400 604.840 2095.600 606.240 ;
        RECT 4.000 603.520 2096.000 604.840 ;
        RECT 4.400 602.120 2095.600 603.520 ;
        RECT 4.000 600.800 2096.000 602.120 ;
        RECT 4.400 599.400 2095.600 600.800 ;
        RECT 4.000 598.080 2096.000 599.400 ;
        RECT 4.400 596.680 2095.600 598.080 ;
        RECT 4.000 595.360 2096.000 596.680 ;
        RECT 4.400 593.960 2095.600 595.360 ;
        RECT 4.000 592.640 2096.000 593.960 ;
        RECT 4.400 591.240 2095.600 592.640 ;
        RECT 4.000 589.920 2096.000 591.240 ;
        RECT 4.400 588.520 2095.600 589.920 ;
        RECT 4.000 587.200 2096.000 588.520 ;
        RECT 4.400 585.800 2095.600 587.200 ;
        RECT 4.000 584.480 2096.000 585.800 ;
        RECT 4.400 583.080 2095.600 584.480 ;
        RECT 4.000 581.760 2096.000 583.080 ;
        RECT 4.400 580.360 2095.600 581.760 ;
        RECT 4.000 579.040 2096.000 580.360 ;
        RECT 4.400 577.640 2095.600 579.040 ;
        RECT 4.000 576.320 2096.000 577.640 ;
        RECT 4.400 574.920 2095.600 576.320 ;
        RECT 4.000 573.600 2096.000 574.920 ;
        RECT 4.400 572.200 2095.600 573.600 ;
        RECT 4.000 570.880 2096.000 572.200 ;
        RECT 4.400 569.480 2095.600 570.880 ;
        RECT 4.000 568.160 2096.000 569.480 ;
        RECT 4.400 566.760 2095.600 568.160 ;
        RECT 4.000 565.440 2096.000 566.760 ;
        RECT 4.400 564.040 2095.600 565.440 ;
        RECT 4.000 562.720 2096.000 564.040 ;
        RECT 4.400 561.320 2095.600 562.720 ;
        RECT 4.000 560.000 2096.000 561.320 ;
        RECT 4.400 558.600 2095.600 560.000 ;
        RECT 4.000 557.280 2096.000 558.600 ;
        RECT 4.400 555.880 2095.600 557.280 ;
        RECT 4.000 554.560 2096.000 555.880 ;
        RECT 4.400 553.160 2095.600 554.560 ;
        RECT 4.000 551.840 2096.000 553.160 ;
        RECT 4.400 550.440 2095.600 551.840 ;
        RECT 4.000 549.120 2096.000 550.440 ;
        RECT 4.400 547.720 2095.600 549.120 ;
        RECT 4.000 546.400 2096.000 547.720 ;
        RECT 4.400 545.000 2095.600 546.400 ;
        RECT 4.000 543.680 2096.000 545.000 ;
        RECT 4.400 542.280 2095.600 543.680 ;
        RECT 4.000 540.960 2096.000 542.280 ;
        RECT 4.400 539.560 2095.600 540.960 ;
        RECT 4.000 538.240 2096.000 539.560 ;
        RECT 4.400 536.840 2095.600 538.240 ;
        RECT 4.000 535.520 2096.000 536.840 ;
        RECT 4.400 534.120 2095.600 535.520 ;
        RECT 4.000 532.800 2096.000 534.120 ;
        RECT 4.400 531.400 2095.600 532.800 ;
        RECT 4.000 530.080 2096.000 531.400 ;
        RECT 4.400 528.680 2095.600 530.080 ;
        RECT 4.000 527.360 2096.000 528.680 ;
        RECT 4.400 525.960 2095.600 527.360 ;
        RECT 4.000 524.640 2096.000 525.960 ;
        RECT 4.400 523.240 2095.600 524.640 ;
        RECT 4.000 521.920 2096.000 523.240 ;
        RECT 4.400 520.520 2095.600 521.920 ;
        RECT 4.000 519.200 2096.000 520.520 ;
        RECT 4.400 517.800 2095.600 519.200 ;
        RECT 4.000 516.480 2096.000 517.800 ;
        RECT 4.400 515.080 2095.600 516.480 ;
        RECT 4.000 513.760 2096.000 515.080 ;
        RECT 4.400 512.360 2095.600 513.760 ;
        RECT 4.000 511.040 2096.000 512.360 ;
        RECT 4.400 509.640 2095.600 511.040 ;
        RECT 4.000 508.320 2096.000 509.640 ;
        RECT 4.400 506.920 2095.600 508.320 ;
        RECT 4.000 505.600 2096.000 506.920 ;
        RECT 4.400 504.200 2095.600 505.600 ;
        RECT 4.000 502.880 2096.000 504.200 ;
        RECT 4.400 501.480 2095.600 502.880 ;
        RECT 4.000 500.160 2096.000 501.480 ;
        RECT 4.400 498.760 2095.600 500.160 ;
        RECT 4.000 497.440 2096.000 498.760 ;
        RECT 4.400 496.040 2095.600 497.440 ;
        RECT 4.000 494.720 2096.000 496.040 ;
        RECT 4.400 493.320 2095.600 494.720 ;
        RECT 4.000 492.000 2096.000 493.320 ;
        RECT 4.400 490.600 2095.600 492.000 ;
        RECT 4.000 489.280 2096.000 490.600 ;
        RECT 4.400 487.880 2095.600 489.280 ;
        RECT 4.000 486.560 2096.000 487.880 ;
        RECT 4.400 485.160 2095.600 486.560 ;
        RECT 4.000 483.840 2096.000 485.160 ;
        RECT 4.400 482.440 2095.600 483.840 ;
        RECT 4.000 481.120 2096.000 482.440 ;
        RECT 4.400 479.720 2095.600 481.120 ;
        RECT 4.000 478.400 2096.000 479.720 ;
        RECT 4.400 477.000 2095.600 478.400 ;
        RECT 4.000 475.680 2096.000 477.000 ;
        RECT 4.400 474.280 2095.600 475.680 ;
        RECT 4.000 472.960 2096.000 474.280 ;
        RECT 4.400 471.560 2095.600 472.960 ;
        RECT 4.000 470.240 2096.000 471.560 ;
        RECT 4.400 468.840 2095.600 470.240 ;
        RECT 4.000 467.520 2096.000 468.840 ;
        RECT 4.400 466.120 2095.600 467.520 ;
        RECT 4.000 464.800 2096.000 466.120 ;
        RECT 4.400 463.400 2095.600 464.800 ;
        RECT 4.000 462.080 2096.000 463.400 ;
        RECT 4.400 460.680 2095.600 462.080 ;
        RECT 4.000 459.360 2096.000 460.680 ;
        RECT 4.400 457.960 2095.600 459.360 ;
        RECT 4.000 456.640 2096.000 457.960 ;
        RECT 4.400 455.240 2095.600 456.640 ;
        RECT 4.000 453.920 2096.000 455.240 ;
        RECT 4.400 452.520 2095.600 453.920 ;
        RECT 4.000 451.200 2096.000 452.520 ;
        RECT 4.400 449.800 2095.600 451.200 ;
        RECT 4.000 448.480 2096.000 449.800 ;
        RECT 4.400 447.080 2095.600 448.480 ;
        RECT 4.000 445.760 2096.000 447.080 ;
        RECT 4.400 444.360 2095.600 445.760 ;
        RECT 4.000 443.040 2096.000 444.360 ;
        RECT 4.400 441.640 2095.600 443.040 ;
        RECT 4.000 440.320 2096.000 441.640 ;
        RECT 4.400 438.920 2095.600 440.320 ;
        RECT 4.000 437.600 2096.000 438.920 ;
        RECT 4.400 436.200 2095.600 437.600 ;
        RECT 4.000 434.880 2096.000 436.200 ;
        RECT 4.400 433.480 2095.600 434.880 ;
        RECT 4.000 432.160 2096.000 433.480 ;
        RECT 4.400 430.760 2095.600 432.160 ;
        RECT 4.000 429.440 2096.000 430.760 ;
        RECT 4.400 428.040 2095.600 429.440 ;
        RECT 4.000 426.720 2096.000 428.040 ;
        RECT 4.400 425.320 2095.600 426.720 ;
        RECT 4.000 424.000 2096.000 425.320 ;
        RECT 4.400 422.600 2095.600 424.000 ;
        RECT 4.000 421.280 2096.000 422.600 ;
        RECT 4.400 419.880 2095.600 421.280 ;
        RECT 4.000 418.560 2096.000 419.880 ;
        RECT 4.400 417.160 2095.600 418.560 ;
        RECT 4.000 415.840 2096.000 417.160 ;
        RECT 4.400 414.440 2095.600 415.840 ;
        RECT 4.000 413.120 2096.000 414.440 ;
        RECT 4.400 411.720 2095.600 413.120 ;
        RECT 4.000 410.400 2096.000 411.720 ;
        RECT 4.400 409.000 2095.600 410.400 ;
        RECT 4.000 407.680 2096.000 409.000 ;
        RECT 4.400 406.280 2095.600 407.680 ;
        RECT 4.000 404.960 2096.000 406.280 ;
        RECT 4.400 403.560 2095.600 404.960 ;
        RECT 4.000 402.240 2096.000 403.560 ;
        RECT 4.400 400.840 2095.600 402.240 ;
        RECT 4.000 399.520 2096.000 400.840 ;
        RECT 4.400 398.120 2095.600 399.520 ;
        RECT 4.000 396.800 2096.000 398.120 ;
        RECT 4.400 395.400 2095.600 396.800 ;
        RECT 4.000 394.080 2096.000 395.400 ;
        RECT 4.400 392.680 2095.600 394.080 ;
        RECT 4.000 391.360 2096.000 392.680 ;
        RECT 4.400 389.960 2095.600 391.360 ;
        RECT 4.000 388.640 2096.000 389.960 ;
        RECT 4.400 387.240 2095.600 388.640 ;
        RECT 4.000 385.920 2096.000 387.240 ;
        RECT 4.400 384.520 2095.600 385.920 ;
        RECT 4.000 383.200 2096.000 384.520 ;
        RECT 4.400 381.800 2095.600 383.200 ;
        RECT 4.000 380.480 2096.000 381.800 ;
        RECT 4.400 379.080 2095.600 380.480 ;
        RECT 4.000 377.760 2096.000 379.080 ;
        RECT 4.400 376.360 2095.600 377.760 ;
        RECT 4.000 375.040 2096.000 376.360 ;
        RECT 4.400 373.640 2095.600 375.040 ;
        RECT 4.000 372.320 2096.000 373.640 ;
        RECT 4.400 370.920 2095.600 372.320 ;
        RECT 4.000 369.600 2096.000 370.920 ;
        RECT 4.400 368.200 2095.600 369.600 ;
        RECT 4.000 366.880 2096.000 368.200 ;
        RECT 4.400 365.480 2095.600 366.880 ;
        RECT 4.000 364.160 2096.000 365.480 ;
        RECT 4.400 362.760 2095.600 364.160 ;
        RECT 4.000 361.440 2096.000 362.760 ;
        RECT 4.400 360.040 2095.600 361.440 ;
        RECT 4.000 358.720 2096.000 360.040 ;
        RECT 4.400 357.320 2095.600 358.720 ;
        RECT 4.000 356.000 2096.000 357.320 ;
        RECT 4.400 354.600 2095.600 356.000 ;
        RECT 4.000 353.280 2096.000 354.600 ;
        RECT 4.400 351.880 2095.600 353.280 ;
        RECT 4.000 350.560 2096.000 351.880 ;
        RECT 4.400 349.160 2095.600 350.560 ;
        RECT 4.000 347.840 2096.000 349.160 ;
        RECT 4.400 346.440 2095.600 347.840 ;
        RECT 4.000 345.120 2096.000 346.440 ;
        RECT 4.400 343.720 2095.600 345.120 ;
        RECT 4.000 342.400 2096.000 343.720 ;
        RECT 4.400 341.000 2095.600 342.400 ;
        RECT 4.000 339.680 2096.000 341.000 ;
        RECT 4.400 338.280 2095.600 339.680 ;
        RECT 4.000 336.960 2096.000 338.280 ;
        RECT 4.400 335.560 2095.600 336.960 ;
        RECT 4.000 334.240 2096.000 335.560 ;
        RECT 4.400 332.840 2095.600 334.240 ;
        RECT 4.000 331.520 2096.000 332.840 ;
        RECT 4.400 330.120 2095.600 331.520 ;
        RECT 4.000 328.800 2096.000 330.120 ;
        RECT 4.400 327.400 2095.600 328.800 ;
        RECT 4.000 326.080 2096.000 327.400 ;
        RECT 4.400 324.680 2095.600 326.080 ;
        RECT 4.000 323.360 2096.000 324.680 ;
        RECT 4.400 321.960 2095.600 323.360 ;
        RECT 4.000 320.640 2096.000 321.960 ;
        RECT 4.400 319.240 2095.600 320.640 ;
        RECT 4.000 317.920 2096.000 319.240 ;
        RECT 4.400 316.520 2095.600 317.920 ;
        RECT 4.000 315.200 2096.000 316.520 ;
        RECT 4.400 313.800 2095.600 315.200 ;
        RECT 4.000 312.480 2096.000 313.800 ;
        RECT 4.400 311.080 2095.600 312.480 ;
        RECT 4.000 309.760 2096.000 311.080 ;
        RECT 4.400 308.360 2095.600 309.760 ;
        RECT 4.000 307.040 2096.000 308.360 ;
        RECT 4.400 305.640 2095.600 307.040 ;
        RECT 4.000 304.320 2096.000 305.640 ;
        RECT 4.400 302.920 2095.600 304.320 ;
        RECT 4.000 301.600 2096.000 302.920 ;
        RECT 4.400 300.200 2095.600 301.600 ;
        RECT 4.000 298.880 2096.000 300.200 ;
        RECT 4.400 297.480 2095.600 298.880 ;
        RECT 4.000 296.160 2096.000 297.480 ;
        RECT 4.400 294.760 2095.600 296.160 ;
        RECT 4.000 293.440 2096.000 294.760 ;
        RECT 4.400 292.040 2095.600 293.440 ;
        RECT 4.000 290.720 2096.000 292.040 ;
        RECT 4.400 289.320 2095.600 290.720 ;
        RECT 4.000 288.000 2096.000 289.320 ;
        RECT 4.400 286.600 2095.600 288.000 ;
        RECT 4.000 285.280 2096.000 286.600 ;
        RECT 4.400 283.880 2095.600 285.280 ;
        RECT 4.000 282.560 2096.000 283.880 ;
        RECT 4.400 281.160 2095.600 282.560 ;
        RECT 4.000 279.840 2096.000 281.160 ;
        RECT 4.400 278.440 2095.600 279.840 ;
        RECT 4.000 277.120 2096.000 278.440 ;
        RECT 4.400 275.720 2095.600 277.120 ;
        RECT 4.000 274.400 2096.000 275.720 ;
        RECT 4.400 273.000 2095.600 274.400 ;
        RECT 4.000 271.680 2096.000 273.000 ;
        RECT 4.400 270.280 2095.600 271.680 ;
        RECT 4.000 268.960 2096.000 270.280 ;
        RECT 4.400 267.560 2095.600 268.960 ;
        RECT 4.000 266.240 2096.000 267.560 ;
        RECT 4.400 264.840 2095.600 266.240 ;
        RECT 4.000 263.520 2096.000 264.840 ;
        RECT 4.400 262.120 2095.600 263.520 ;
        RECT 4.000 260.800 2096.000 262.120 ;
        RECT 4.400 259.400 2095.600 260.800 ;
        RECT 4.000 258.080 2096.000 259.400 ;
        RECT 4.400 256.680 2095.600 258.080 ;
        RECT 4.000 255.360 2096.000 256.680 ;
        RECT 4.400 253.960 2095.600 255.360 ;
        RECT 4.000 252.640 2096.000 253.960 ;
        RECT 4.400 251.240 2095.600 252.640 ;
        RECT 4.000 249.920 2096.000 251.240 ;
        RECT 4.400 248.520 2095.600 249.920 ;
        RECT 4.000 247.200 2096.000 248.520 ;
        RECT 4.400 245.800 2095.600 247.200 ;
        RECT 4.000 244.480 2096.000 245.800 ;
        RECT 4.400 243.080 2095.600 244.480 ;
        RECT 4.000 241.760 2096.000 243.080 ;
        RECT 4.400 240.360 2095.600 241.760 ;
        RECT 4.000 239.040 2096.000 240.360 ;
        RECT 4.400 237.640 2095.600 239.040 ;
        RECT 4.000 236.320 2096.000 237.640 ;
        RECT 4.400 234.920 2095.600 236.320 ;
        RECT 4.000 233.600 2096.000 234.920 ;
        RECT 4.400 232.200 2095.600 233.600 ;
        RECT 4.000 230.880 2096.000 232.200 ;
        RECT 4.400 229.480 2095.600 230.880 ;
        RECT 4.000 228.160 2096.000 229.480 ;
        RECT 4.400 226.760 2095.600 228.160 ;
        RECT 4.000 225.440 2096.000 226.760 ;
        RECT 4.400 224.040 2095.600 225.440 ;
        RECT 4.000 222.720 2096.000 224.040 ;
        RECT 4.400 221.320 2095.600 222.720 ;
        RECT 4.000 220.000 2096.000 221.320 ;
        RECT 4.400 218.600 2095.600 220.000 ;
        RECT 4.000 217.280 2096.000 218.600 ;
        RECT 4.400 215.880 2095.600 217.280 ;
        RECT 4.000 214.560 2096.000 215.880 ;
        RECT 4.400 213.160 2095.600 214.560 ;
        RECT 4.000 211.840 2096.000 213.160 ;
        RECT 4.400 210.440 2095.600 211.840 ;
        RECT 4.000 209.120 2096.000 210.440 ;
        RECT 4.400 207.720 2095.600 209.120 ;
        RECT 4.000 206.400 2096.000 207.720 ;
        RECT 4.400 205.000 2095.600 206.400 ;
        RECT 4.000 203.680 2096.000 205.000 ;
        RECT 4.400 202.280 2095.600 203.680 ;
        RECT 4.000 200.960 2096.000 202.280 ;
        RECT 4.400 199.560 2095.600 200.960 ;
        RECT 4.000 198.240 2096.000 199.560 ;
        RECT 4.400 196.840 2095.600 198.240 ;
        RECT 4.000 195.520 2096.000 196.840 ;
        RECT 4.400 194.120 2095.600 195.520 ;
        RECT 4.000 192.800 2096.000 194.120 ;
        RECT 4.400 191.400 2095.600 192.800 ;
        RECT 4.000 190.080 2096.000 191.400 ;
        RECT 4.400 188.680 2095.600 190.080 ;
        RECT 4.000 187.360 2096.000 188.680 ;
        RECT 4.400 185.960 2095.600 187.360 ;
        RECT 4.000 184.640 2096.000 185.960 ;
        RECT 4.400 183.240 2095.600 184.640 ;
        RECT 4.000 181.920 2096.000 183.240 ;
        RECT 4.400 180.520 2095.600 181.920 ;
        RECT 4.000 179.200 2096.000 180.520 ;
        RECT 4.400 177.800 2095.600 179.200 ;
        RECT 4.000 176.480 2096.000 177.800 ;
        RECT 4.400 175.080 2095.600 176.480 ;
        RECT 4.000 173.760 2096.000 175.080 ;
        RECT 4.400 172.360 2095.600 173.760 ;
        RECT 4.000 171.040 2096.000 172.360 ;
        RECT 4.400 169.640 2095.600 171.040 ;
        RECT 4.000 168.320 2096.000 169.640 ;
        RECT 4.400 166.920 2095.600 168.320 ;
        RECT 4.000 165.600 2096.000 166.920 ;
        RECT 4.400 164.200 2095.600 165.600 ;
        RECT 4.000 162.880 2096.000 164.200 ;
        RECT 4.400 161.480 2095.600 162.880 ;
        RECT 4.000 160.160 2096.000 161.480 ;
        RECT 4.400 158.760 2095.600 160.160 ;
        RECT 4.000 157.440 2096.000 158.760 ;
        RECT 4.400 156.040 2095.600 157.440 ;
        RECT 4.000 154.720 2096.000 156.040 ;
        RECT 4.400 153.320 2095.600 154.720 ;
        RECT 4.000 152.000 2096.000 153.320 ;
        RECT 4.400 150.600 2095.600 152.000 ;
        RECT 4.000 149.280 2096.000 150.600 ;
        RECT 4.400 147.880 2095.600 149.280 ;
        RECT 4.000 146.560 2096.000 147.880 ;
        RECT 4.400 145.160 2095.600 146.560 ;
        RECT 4.000 143.840 2096.000 145.160 ;
        RECT 4.400 142.440 2095.600 143.840 ;
        RECT 4.000 141.120 2096.000 142.440 ;
        RECT 4.400 139.720 2095.600 141.120 ;
        RECT 4.000 138.400 2096.000 139.720 ;
        RECT 4.400 137.000 2095.600 138.400 ;
        RECT 4.000 135.680 2096.000 137.000 ;
        RECT 4.400 134.280 2095.600 135.680 ;
        RECT 4.000 132.960 2096.000 134.280 ;
        RECT 4.400 131.560 2095.600 132.960 ;
        RECT 4.000 130.240 2096.000 131.560 ;
        RECT 4.400 128.840 2095.600 130.240 ;
        RECT 4.000 127.520 2096.000 128.840 ;
        RECT 4.400 126.120 2095.600 127.520 ;
        RECT 4.000 124.800 2096.000 126.120 ;
        RECT 4.400 123.400 2095.600 124.800 ;
        RECT 4.000 122.080 2096.000 123.400 ;
        RECT 4.400 120.680 2095.600 122.080 ;
        RECT 4.000 119.360 2096.000 120.680 ;
        RECT 4.400 117.960 2095.600 119.360 ;
        RECT 4.000 116.640 2096.000 117.960 ;
        RECT 4.400 115.240 2095.600 116.640 ;
        RECT 4.000 113.920 2096.000 115.240 ;
        RECT 4.400 112.520 2095.600 113.920 ;
        RECT 4.000 111.200 2096.000 112.520 ;
        RECT 4.400 109.800 2095.600 111.200 ;
        RECT 4.000 108.480 2096.000 109.800 ;
        RECT 4.400 107.080 2095.600 108.480 ;
        RECT 4.000 105.760 2096.000 107.080 ;
        RECT 4.400 104.360 2095.600 105.760 ;
        RECT 4.000 103.040 2096.000 104.360 ;
        RECT 4.400 101.640 2095.600 103.040 ;
        RECT 4.000 100.320 2096.000 101.640 ;
        RECT 4.400 98.920 2095.600 100.320 ;
        RECT 4.000 97.600 2096.000 98.920 ;
        RECT 4.400 96.200 2095.600 97.600 ;
        RECT 4.000 94.880 2096.000 96.200 ;
        RECT 4.400 93.480 2095.600 94.880 ;
        RECT 4.000 92.160 2096.000 93.480 ;
        RECT 4.400 90.760 2095.600 92.160 ;
        RECT 4.000 89.440 2096.000 90.760 ;
        RECT 4.400 88.040 2095.600 89.440 ;
        RECT 4.000 86.720 2096.000 88.040 ;
        RECT 4.400 85.320 2095.600 86.720 ;
        RECT 4.000 84.000 2096.000 85.320 ;
        RECT 4.400 82.600 2095.600 84.000 ;
        RECT 4.000 81.280 2096.000 82.600 ;
        RECT 4.400 79.880 2095.600 81.280 ;
        RECT 4.000 78.560 2096.000 79.880 ;
        RECT 4.400 77.160 2095.600 78.560 ;
        RECT 4.000 75.840 2096.000 77.160 ;
        RECT 4.400 74.440 2095.600 75.840 ;
        RECT 4.000 73.120 2096.000 74.440 ;
        RECT 4.400 71.720 2095.600 73.120 ;
        RECT 4.000 70.400 2096.000 71.720 ;
        RECT 4.400 69.000 2095.600 70.400 ;
        RECT 4.000 67.680 2096.000 69.000 ;
        RECT 4.400 66.280 2095.600 67.680 ;
        RECT 4.000 64.960 2096.000 66.280 ;
        RECT 4.400 63.560 2095.600 64.960 ;
        RECT 4.000 62.240 2096.000 63.560 ;
        RECT 4.400 60.840 2095.600 62.240 ;
        RECT 4.000 59.520 2096.000 60.840 ;
        RECT 4.400 58.120 2095.600 59.520 ;
        RECT 4.000 56.800 2096.000 58.120 ;
        RECT 4.400 55.400 2095.600 56.800 ;
        RECT 4.000 54.080 2096.000 55.400 ;
        RECT 4.400 52.680 2095.600 54.080 ;
        RECT 4.000 51.360 2096.000 52.680 ;
        RECT 4.400 49.960 2095.600 51.360 ;
        RECT 4.000 48.640 2096.000 49.960 ;
        RECT 4.400 47.240 2095.600 48.640 ;
        RECT 4.000 45.920 2096.000 47.240 ;
        RECT 4.400 44.520 2095.600 45.920 ;
        RECT 4.000 43.200 2096.000 44.520 ;
        RECT 4.400 41.800 2095.600 43.200 ;
        RECT 4.000 40.480 2096.000 41.800 ;
        RECT 4.400 39.080 2095.600 40.480 ;
        RECT 4.000 37.760 2096.000 39.080 ;
        RECT 4.400 36.360 2095.600 37.760 ;
        RECT 4.000 35.040 2096.000 36.360 ;
        RECT 4.400 33.640 2095.600 35.040 ;
        RECT 4.000 32.320 2096.000 33.640 ;
        RECT 4.400 30.920 2095.600 32.320 ;
        RECT 4.000 29.600 2096.000 30.920 ;
        RECT 4.400 28.200 2095.600 29.600 ;
        RECT 4.000 26.880 2096.000 28.200 ;
        RECT 4.400 25.480 2095.600 26.880 ;
        RECT 4.000 24.160 2096.000 25.480 ;
        RECT 4.400 22.760 2095.600 24.160 ;
        RECT 4.000 21.440 2096.000 22.760 ;
        RECT 4.400 20.040 2095.600 21.440 ;
        RECT 4.000 18.720 2096.000 20.040 ;
        RECT 4.400 17.320 2095.600 18.720 ;
        RECT 4.000 16.000 2096.000 17.320 ;
        RECT 4.400 14.600 2095.600 16.000 ;
        RECT 4.000 13.280 2096.000 14.600 ;
        RECT 4.400 11.880 2095.600 13.280 ;
        RECT 4.000 10.560 2096.000 11.880 ;
        RECT 4.400 9.160 2095.600 10.560 ;
        RECT 4.000 7.840 2096.000 9.160 ;
        RECT 4.400 6.440 2095.600 7.840 ;
        RECT 4.000 5.120 2096.000 6.440 ;
        RECT 4.400 3.720 2095.600 5.120 ;
        RECT 4.000 2.400 2096.000 3.720 ;
        RECT 4.400 1.535 2095.600 2.400 ;
      LAYER met4 ;
        RECT 350.815 628.960 2083.505 638.345 ;
        RECT 350.815 10.240 404.640 628.960 ;
        RECT 407.040 10.240 481.440 628.960 ;
        RECT 483.840 10.240 558.240 628.960 ;
        RECT 560.640 10.240 635.040 628.960 ;
        RECT 637.440 10.240 711.840 628.960 ;
        RECT 714.240 10.240 788.640 628.960 ;
        RECT 791.040 10.240 865.440 628.960 ;
        RECT 867.840 10.240 942.240 628.960 ;
        RECT 944.640 10.240 1019.040 628.960 ;
        RECT 1021.440 10.240 1095.840 628.960 ;
        RECT 1098.240 10.240 1172.640 628.960 ;
        RECT 1175.040 10.240 1249.440 628.960 ;
        RECT 1251.840 10.240 1326.240 628.960 ;
        RECT 1328.640 10.240 1403.040 628.960 ;
        RECT 1405.440 10.240 1479.840 628.960 ;
        RECT 1482.240 10.240 1556.640 628.960 ;
        RECT 1559.040 10.240 1633.440 628.960 ;
        RECT 1635.840 10.240 1710.240 628.960 ;
        RECT 1712.640 10.240 1787.040 628.960 ;
        RECT 1789.440 10.240 1863.840 628.960 ;
        RECT 1866.240 10.240 1940.640 628.960 ;
        RECT 1943.040 10.240 2017.440 628.960 ;
        RECT 2019.840 10.240 2083.505 628.960 ;
        RECT 350.815 1.535 2083.505 10.240 ;
  END
END vliw
END LIBRARY

