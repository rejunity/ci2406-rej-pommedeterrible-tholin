* NGSPICE file created from wrapped_6502.ext - technology: sky130B

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_4 abstract view
.subckt sky130_fd_sc_hd__and2b_4 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_4 abstract view
.subckt sky130_fd_sc_hd__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_4 abstract view
.subckt sky130_fd_sc_hd__nor4b_4 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

.subckt wrapped_6502 custom_settings[0] custom_settings[1] io_in[0] io_in[10] io_in[11]
+ io_in[12] io_in[13] io_in[14] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19]
+ io_in[1] io_in[20] io_in[21] io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[27]
+ io_in[28] io_in[29] io_in[2] io_in[30] io_in[31] io_in[32] io_in[33] io_in[34] io_in[35]
+ io_in[3] io_in[4] io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb io_out[0]
+ io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15] io_out[16] io_out[17]
+ io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22] io_out[23] io_out[24]
+ io_out[25] io_out[26] io_out[27] io_out[28] io_out[29] io_out[2] io_out[30] io_out[31]
+ io_out[32] io_out[33] io_out[34] io_out[35] io_out[3] io_out[4] io_out[5] io_out[6]
+ io_out[7] io_out[8] io_out[9] rst_n vccd1 vssd1 wb_clk_i
X_2106_ _2226_/CLK hold6/X vssd1 vssd1 vccd1 vccd1 hold5/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2037_ _1273_/X _2036_/Y _2043_/B vssd1 vssd1 vccd1 vccd1 _2037_/X sky130_fd_sc_hd__a21o_1
XTAP_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1534__A _1548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout75_A _1871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1445__B2 _2117_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1270_ _1728_/B _1945_/A vssd1 vssd1 vccd1 vccd1 _2001_/A sky130_fd_sc_hd__nand2_4
XFILLER_0_3_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1436__A1 _1025_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1606_ _1606_/A _1606_/B vssd1 vssd1 vccd1 vccd1 _1607_/B sky130_fd_sc_hd__and2_1
X_1468_ _1468_/A vssd1 vssd1 vccd1 vccd1 _1468_/Y sky130_fd_sc_hd__inv_2
X_1537_ _2116_/Q _1538_/B vssd1 vssd1 vccd1 vccd1 _1539_/A sky130_fd_sc_hd__nand2_1
X_1399_ _1830_/B _1415_/A3 _1340_/B _1830_/C vssd1 vssd1 vccd1 vccd1 _1417_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_49_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1427__B2 _2161_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold181 _1710_/X vssd1 vssd1 vccd1 vccd1 _2115_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold192 _1699_/X vssd1 vssd1 vccd1 vccd1 _2108_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold170 _2010_/X vssd1 vssd1 vccd1 vccd1 _2191_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1203__S _1994_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1253_ _1728_/B _1253_/B vssd1 vssd1 vccd1 vccd1 _2015_/A sky130_fd_sc_hd__nand2_2
X_1322_ _1486_/D _1365_/A _1340_/B _1907_/S vssd1 vssd1 vccd1 vccd1 _1414_/B sky130_fd_sc_hd__a22o_1
X_1184_ hold59/A _1499_/B _1182_/X _1882_/A vssd1 vssd1 vccd1 vccd1 _1186_/A sky130_fd_sc_hd__o211ai_2
XFILLER_0_27_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1896__A1 _1871_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1820__B2 _2053_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1940_ hold7/X _1920_/Y _1939_/X vssd1 vssd1 vccd1 vccd1 hold8/A sky130_fd_sc_hd__a21o_1
X_1871_ _1871_/A _1871_/B vssd1 vssd1 vccd1 vccd1 _2159_/D sky130_fd_sc_hd__and2_1
XFILLER_0_56_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1811__A1 _2053_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1305_ _1306_/A _1306_/B vssd1 vssd1 vccd1 vccd1 _2001_/C sky130_fd_sc_hd__and2_2
XANTENNA__1878__A1 _1864_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1236_ _1114_/B _1821_/B _1821_/A _1236_/D vssd1 vssd1 vccd1 vccd1 _1245_/C sky130_fd_sc_hd__and4b_2
XFILLER_0_19_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1167_ hold15/A hold63/A _1499_/B vssd1 vssd1 vccd1 vccd1 _1167_/X sky130_fd_sc_hd__mux2_1
X_1098_ _1236_/D _1114_/B _1821_/B _1821_/A vssd1 vssd1 vccd1 vccd1 _1121_/B sky130_fd_sc_hd__or4bb_4
XFILLER_0_19_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1717__A _1922_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2070_ hold39/X _1519_/X _2075_/S vssd1 vssd1 vccd1 vccd1 hold40/A sky130_fd_sc_hd__mux2_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1088__A2 _1922_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1923_ _1923_/A _1923_/B vssd1 vssd1 vccd1 vccd1 _1923_/Y sky130_fd_sc_hd__nand2_1
X_1785_ _1785_/A _1785_/B _1785_/C _1785_/D vssd1 vssd1 vccd1 vccd1 _1785_/Y sky130_fd_sc_hd__nand4_1
XFILLER_0_31_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1854_ hold186/X _1181_/X _1862_/S vssd1 vssd1 vccd1 vccd1 _1854_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_12_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2199_ _1233_/A _2199_/D vssd1 vssd1 vccd1 vccd1 _2199_/Q sky130_fd_sc_hd__dfxtp_1
X_1219_ hold200/X _1828_/B _1150_/S _1788_/A _1218_/X vssd1 vssd1 vccd1 vccd1 _1219_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_47_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold30 hold30/A vssd1 vssd1 vccd1 vccd1 hold30/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 hold41/A vssd1 vssd1 vccd1 vccd1 hold41/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold63 hold63/A vssd1 vssd1 vccd1 vccd1 hold63/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1272__A _1728_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold52 hold52/A vssd1 vssd1 vccd1 vccd1 hold52/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 hold74/A vssd1 vssd1 vccd1 vccd1 hold74/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold96 hold96/A vssd1 vssd1 vccd1 vccd1 hold96/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 hold85/A vssd1 vssd1 vccd1 vccd1 hold85/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1570_ _1570_/A _1570_/B vssd1 vssd1 vccd1 vccd1 _1571_/B sky130_fd_sc_hd__nand2_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2053_ hold73/X _2054_/A2 _1995_/B _2053_/B2 vssd1 vssd1 vccd1 vccd1 hold74/A sky130_fd_sc_hd__a22o_1
X_2122_ _2164_/CLK _2122_/D vssd1 vssd1 vccd1 vccd1 _2122_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1906_ _1028_/Y hold194/X _1912_/A vssd1 vssd1 vccd1 vccd1 _1906_/X sky130_fd_sc_hd__mux2_1
X_1768_ _2053_/B2 _1772_/A _1767_/Y _1820_/A2 _1763_/A vssd1 vssd1 vccd1 vccd1 _1768_/X
+ sky130_fd_sc_hd__a32o_1
X_1837_ _1863_/A _1837_/B vssd1 vssd1 vccd1 vccd1 _2137_/D sky130_fd_sc_hd__and2_1
XFILLER_0_12_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1699_ _1239_/B _1698_/X _1920_/A vssd1 vssd1 vccd1 vccd1 _1699_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_12_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput31 _1438_/X vssd1 vssd1 vccd1 vccd1 io_out[23] sky130_fd_sc_hd__buf_12
Xoutput20 _1219_/X vssd1 vssd1 vccd1 vccd1 io_out[13] sky130_fd_sc_hd__buf_12
Xoutput42 _1190_/X vssd1 vssd1 vccd1 vccd1 io_out[5] sky130_fd_sc_hd__buf_12
XFILLER_0_73_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1876__S _1912_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1622_ _1622_/A _1622_/B vssd1 vssd1 vccd1 vccd1 _1622_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_26_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1553_ _2049_/A input5/X vssd1 vssd1 vccd1 vccd1 _2093_/D sky130_fd_sc_hd__and2_1
X_1484_ _1116_/C _1119_/A _1716_/B _2108_/Q vssd1 vssd1 vccd1 vccd1 _1488_/A sky130_fd_sc_hd__o31a_1
XTAP_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2105_ _2225_/CLK hold20/X vssd1 vssd1 vccd1 vccd1 hold19/A sky130_fd_sc_hd__dfxtp_1
X_2036_ _2036_/A _2036_/B vssd1 vssd1 vccd1 vccd1 _2036_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_64_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1678__C1 _1448_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1381__A1 _1826_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1536_ hold41/X _1535_/X _1550_/S vssd1 vssd1 vccd1 vccd1 hold42/A sky130_fd_sc_hd__mux2_1
X_1605_ _1606_/A _1606_/B vssd1 vssd1 vccd1 vccd1 _1691_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_10_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1467_ _1467_/A _1467_/B _1920_/B _1467_/D vssd1 vssd1 vccd1 vccd1 _1468_/A sky130_fd_sc_hd__or4_4
XFILLER_0_38_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1398_ _1487_/A _1365_/A _1403_/A2 _1129_/B _1418_/B vssd1 vssd1 vccd1 vccd1 _1413_/C
+ sky130_fd_sc_hd__a221o_1
X_2019_ _2019_/A _2019_/B vssd1 vssd1 vccd1 vccd1 _2019_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_37_307 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_362 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1545__A _2108_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold193 _2116_/Q vssd1 vssd1 vccd1 vccd1 hold193/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold171 _2114_/Q vssd1 vssd1 vccd1 vccd1 hold171/X sky130_fd_sc_hd__buf_1
Xhold160 _2117_/Q vssd1 vssd1 vccd1 vccd1 _1545_/B sky130_fd_sc_hd__buf_2
Xhold182 _2147_/Q vssd1 vssd1 vccd1 vccd1 hold182/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1252_ _1728_/B _1253_/B vssd1 vssd1 vccd1 vccd1 _1980_/A sky130_fd_sc_hd__and2_2
Xclkbuf_4_12_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _2219_/CLK sky130_fd_sc_hd__clkbuf_8
X_1321_ _1716_/A _1403_/A2 _1320_/Y _1415_/A3 vssd1 vssd1 vccd1 vccd1 _1410_/B sky130_fd_sc_hd__a22o_1
X_1183_ _1174_/B _1174_/C hold75/A vssd1 vssd1 vccd1 vccd1 _1183_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_19_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1519_ _1518_/X _1542_/A vssd1 vssd1 vccd1 vccd1 _1519_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold232_A _2165_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1870_ _1871_/A _1870_/B vssd1 vssd1 vccd1 vccd1 _2158_/D sky130_fd_sc_hd__and2_1
XFILLER_0_56_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1304_ _1980_/B _2001_/A _2015_/D vssd1 vssd1 vccd1 vccd1 _1304_/X sky130_fd_sc_hd__o21a_1
X_1235_ _1921_/A _2003_/A vssd1 vssd1 vccd1 vccd1 _1735_/A sky130_fd_sc_hd__nor2_1
X_1166_ _1757_/A _1149_/Y _1165_/X vssd1 vssd1 vccd1 vccd1 _1166_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_19_73 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1263__A0 _1868_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1097_ _1236_/D _1114_/B _1821_/B _1821_/A vssd1 vssd1 vccd1 vccd1 _1097_/X sky130_fd_sc_hd__and4bb_1
XFILLER_0_19_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1999_ hold214/X _2001_/A _1996_/Y _1997_/B _2188_/Q vssd1 vssd1 vccd1 vccd1 _1999_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_42_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1717__B _1717_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1922_ _1994_/A _1922_/B vssd1 vssd1 vccd1 vccd1 _1922_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_8_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1784_ _1784_/A _1808_/B vssd1 vssd1 vccd1 vccd1 _1785_/D sky130_fd_sc_hd__nand2_1
XFILLER_0_24_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1853_ _1863_/A _1853_/B vssd1 vssd1 vccd1 vccd1 _2145_/D sky130_fd_sc_hd__and2_1
XFILLER_0_12_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2198_ _2201_/CLK _2198_/D vssd1 vssd1 vccd1 vccd1 _2198_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1484__B1 _2108_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1149_ _1467_/A _1149_/B _1149_/C _1827_/B vssd1 vssd1 vccd1 vccd1 _1149_/Y sky130_fd_sc_hd__nor4_4
X_1218_ _1130_/B _1866_/B _1207_/X hold218/X vssd1 vssd1 vccd1 vccd1 _1218_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1787__A1 _2053_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold20 hold20/A vssd1 vssd1 vccd1 vccd1 hold20/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 hold75/A vssd1 vssd1 vccd1 vccd1 hold75/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 hold31/A vssd1 vssd1 vccd1 vccd1 hold31/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 hold42/A vssd1 vssd1 vccd1 vccd1 hold42/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 hold53/A vssd1 vssd1 vccd1 vccd1 hold53/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 hold97/A vssd1 vssd1 vccd1 vccd1 hold97/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 hold64/A vssd1 vssd1 vccd1 vccd1 hold64/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold86 hold86/A vssd1 vssd1 vccd1 vccd1 hold86/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1699__S _1920_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1447__B _2164_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2052_ hold87/X _2054_/A2 _1995_/A _1296_/B vssd1 vssd1 vccd1 vccd1 hold88/A sky130_fd_sc_hd__a22o_1
X_2121_ _2164_/CLK _2121_/D vssd1 vssd1 vccd1 vccd1 _2121_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1905_ _1912_/A _1028_/A hold188/X _1921_/B _1881_/X vssd1 vssd1 vccd1 vccd1 _1908_/S
+ sky130_fd_sc_hd__o41a_1
XFILLER_0_29_298 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1769__A1 _2117_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1698_ _1690_/X _1695_/X _1696_/Y _1697_/X vssd1 vssd1 vccd1 vccd1 _1698_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_32_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1836_ hold218/X _1219_/X _1862_/S vssd1 vssd1 vccd1 vccd1 _1836_/X sky130_fd_sc_hd__mux2_1
X_1767_ _1767_/A _1767_/B _1767_/C _1767_/D vssd1 vssd1 vccd1 vccd1 _1767_/Y sky130_fd_sc_hd__nand4_1
XFILLER_0_4_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1548__A _1548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1283__A _1728_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput32 _1440_/X vssd1 vssd1 vccd1 vccd1 io_out[24] sky130_fd_sc_hd__buf_12
XFILLER_0_31_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput21 _1217_/X vssd1 vssd1 vccd1 vccd1 io_out[14] sky130_fd_sc_hd__buf_12
Xoutput43 _1181_/X vssd1 vssd1 vccd1 vccd1 io_out[6] sky130_fd_sc_hd__buf_12
X_1552_ _2000_/A input4/X vssd1 vssd1 vccd1 vccd1 _2092_/D sky130_fd_sc_hd__and2_1
X_1621_ _2113_/Q _1460_/A _1620_/X vssd1 vssd1 vccd1 vccd1 _1622_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__1620__B1 _1796_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2104_ _2226_/CLK hold32/X vssd1 vssd1 vccd1 vccd1 hold31/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__1921__A _1921_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1483_ _2192_/Q _2160_/Q _1482_/Y _2186_/Q vssd1 vssd1 vccd1 vccd1 _1483_/X sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_4_10_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2035_ _2057_/A _2035_/B vssd1 vssd1 vccd1 vccd1 _2199_/D sky130_fd_sc_hd__and2_1
XFILLER_0_43_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1914__B2 _1912_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1819_ _1819_/A _1819_/B vssd1 vssd1 vccd1 vccd1 _1819_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1905__A1 _1912_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1535_ _1548_/A _1808_/A _1542_/A _1534_/Y vssd1 vssd1 vccd1 vccd1 _1535_/X sky130_fd_sc_hd__o211a_1
X_1604_ _1650_/B _1603_/B _1602_/X _1603_/Y vssd1 vssd1 vccd1 vccd1 _1606_/B sky130_fd_sc_hd__a211o_1
XFILLER_0_10_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1466_ _1032_/Y _1448_/B _1378_/C _1458_/A vssd1 vssd1 vccd1 vccd1 _1467_/D sky130_fd_sc_hd__a211o_1
X_1397_ _1075_/C _2054_/A2 _1960_/B _1317_/Y vssd1 vssd1 vccd1 vccd1 _1418_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_54_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2018_ _2015_/C _1984_/C _1955_/B _2015_/Y _2017_/X vssd1 vssd1 vccd1 vccd1 _2019_/B
+ sky130_fd_sc_hd__a311o_1
XFILLER_0_49_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold161 _2182_/Q vssd1 vssd1 vccd1 vccd1 _1982_/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1545__B _1545_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold194 _2113_/Q vssd1 vssd1 vccd1 vccd1 hold194/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold172 _1709_/X vssd1 vssd1 vccd1 vccd1 _2114_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold150 _1987_/X vssd1 vssd1 vccd1 vccd1 _2184_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold183 _2148_/Q vssd1 vssd1 vccd1 vccd1 hold183/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1320_ _1345_/A _1320_/B vssd1 vssd1 vccd1 vccd1 _1320_/Y sky130_fd_sc_hd__nor2_1
X_1251_ _1866_/B _2169_/Q _2166_/Q vssd1 vssd1 vccd1 vccd1 _1253_/B sky130_fd_sc_hd__mux2_1
X_1182_ _1174_/B _1174_/C hold49/A vssd1 vssd1 vccd1 vccd1 _1182_/X sky130_fd_sc_hd__a21o_1
XANTENNA__2067__B1 _2003_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1518_ _1517_/A _1515_/X _1516_/Y _1517_/Y vssd1 vssd1 vccd1 vccd1 _1518_/X sky130_fd_sc_hd__o31a_1
XFILLER_0_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1449_ _1450_/A _1829_/B vssd1 vssd1 vccd1 vccd1 _1650_/A sky130_fd_sc_hd__and2_1
XANTENNA__1365__B _1826_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2058__B1 _2003_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold225_A _1784_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_300 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1303_ _2015_/D vssd1 vssd1 vccd1 vccd1 _1303_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_10_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1096_ _1094_/X _1095_/X _1499_/A vssd1 vssd1 vccd1 vccd1 _1096_/X sky130_fd_sc_hd__mux2_1
X_1234_ input2/X _1233_/Y _1232_/X _1231_/Y vssd1 vssd1 vccd1 vccd1 _1234_/Y sky130_fd_sc_hd__a211oi_2
X_1165_ hold180/X _1149_/B _1162_/X _1467_/A _1164_/X vssd1 vssd1 vccd1 vccd1 _1165_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_19_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1998_ _1996_/Y _1997_/X _2000_/A vssd1 vssd1 vccd1 vccd1 _2187_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_42_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_15_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1921_ _1921_/A _1921_/B vssd1 vssd1 vccd1 vccd1 _2031_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_29_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1852_ hold190/X _1190_/X _1862_/S vssd1 vssd1 vccd1 vccd1 _1853_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_52_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1783_ _2111_/Q _1135_/A _1776_/X _2136_/Q _1717_/B vssd1 vssd1 vccd1 vccd1 _1785_/C
+ sky130_fd_sc_hd__a221oi_2
XFILLER_0_24_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2197_ _2219_/CLK _2197_/D vssd1 vssd1 vccd1 vccd1 _2197_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1148_ _1467_/A _1096_/X _1149_/B _1545_/B _1147_/X vssd1 vssd1 vccd1 vccd1 _1148_/X
+ sky130_fd_sc_hd__a221o_1
X_1217_ hold194/X _1828_/B _1150_/S _1794_/A _1216_/X vssd1 vssd1 vccd1 vccd1 _1217_/X
+ sky130_fd_sc_hd__a221o_2
X_1079_ _1377_/A _1080_/B _1144_/B _1345_/A vssd1 vssd1 vccd1 vccd1 _1079_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_62_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold54 hold54/A vssd1 vssd1 vccd1 vccd1 hold54/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 hold32/A vssd1 vssd1 vccd1 vccd1 hold32/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 hold65/A vssd1 vssd1 vccd1 vccd1 hold65/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 hold43/A vssd1 vssd1 vccd1 vccd1 hold43/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 hold21/A vssd1 vssd1 vccd1 vccd1 hold21/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 hold76/A vssd1 vssd1 vccd1 vccd1 hold76/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold10 hold10/A vssd1 vssd1 vccd1 vccd1 hold10/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 hold87/A vssd1 vssd1 vccd1 vccd1 hold87/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold98 hold98/A vssd1 vssd1 vccd1 vccd1 hold98/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1728__B _1728_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2120_ _2164_/CLK _2120_/D vssd1 vssd1 vccd1 vccd1 _2120_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2051_ _1912_/A _2031_/A _2050_/Y _2057_/A vssd1 vssd1 vccd1 vccd1 _2206_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_16_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1919__A _1920_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1904_ hold167/X _1900_/X _1903_/X _2057_/A vssd1 vssd1 vccd1 vccd1 _1904_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_32_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1835_ _1863_/A _1835_/B vssd1 vssd1 vccd1 vccd1 _2136_/D sky130_fd_sc_hd__and2_1
XFILLER_0_25_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1926__C1 _1871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1697_ _1697_/A _1697_/B _1697_/C _1697_/D vssd1 vssd1 vccd1 vccd1 _1697_/X sky130_fd_sc_hd__and4_1
X_1766_ _1767_/B _1767_/C _1767_/D _1767_/A vssd1 vssd1 vccd1 vccd1 _1772_/A sky130_fd_sc_hd__a31o_1
XFILLER_0_4_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1209__A1 _1545_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput33 _1443_/X vssd1 vssd1 vccd1 vccd1 io_out[25] sky130_fd_sc_hd__buf_12
Xoutput22 _1215_/X vssd1 vssd1 vccd1 vccd1 io_out[15] sky130_fd_sc_hd__buf_12
XFILLER_0_9_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput44 _1173_/X vssd1 vssd1 vccd1 vccd1 io_out[7] sky130_fd_sc_hd__buf_12
XFILLER_0_73_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1551_ _2000_/A input3/X vssd1 vssd1 vccd1 vccd1 _2091_/D sky130_fd_sc_hd__and2_1
X_1482_ _2192_/Q _2189_/Q vssd1 vssd1 vccd1 vccd1 _1482_/Y sky130_fd_sc_hd__nor2_1
X_1620_ _2138_/Q _1776_/A _1796_/A _1469_/X vssd1 vssd1 vccd1 vccd1 _1620_/X sky130_fd_sc_hd__a22o_1
X_2103_ _2223_/CLK hold16/X vssd1 vssd1 vccd1 vccd1 hold15/A sky130_fd_sc_hd__dfxtp_1
XTAP_169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2034_ hold184/X _2043_/B _2031_/X _1273_/X vssd1 vssd1 vccd1 vccd1 _2035_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_9_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1818_ _1871_/B _1808_/B _1806_/B hold116/X _1817_/X vssd1 vssd1 vccd1 vccd1 _1819_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_4_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1749_ _1749_/A _1749_/B _1749_/C _1749_/D vssd1 vssd1 vccd1 vccd1 _1749_/Y sky130_fd_sc_hd__nand4_1
XFILLER_0_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1534_ _1548_/A _1534_/B vssd1 vssd1 vccd1 vccd1 _1534_/Y sky130_fd_sc_hd__nand2_1
X_1603_ _1651_/A _1603_/B vssd1 vssd1 vccd1 vccd1 _1603_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_38_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1465_ _1486_/A _1465_/B vssd1 vssd1 vccd1 vccd1 _1920_/B sky130_fd_sc_hd__or2_4
XFILLER_0_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2017_ _2001_/A _1984_/B _1996_/C _2008_/Y vssd1 vssd1 vccd1 vccd1 _2017_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_49_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1396_ _1413_/B _1396_/B vssd1 vssd1 vccd1 vccd1 _1408_/C sky130_fd_sc_hd__or2_1
XFILLER_0_70_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold162 _1983_/X vssd1 vssd1 vccd1 vccd1 _2182_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2003__A _2003_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold151 hold243/X vssd1 vssd1 vccd1 vccd1 _1029_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold140 _1727_/X vssd1 vssd1 vccd1 vccd1 _2119_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold173 _2190_/Q vssd1 vssd1 vccd1 vccd1 _2006_/A sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold184 _2199_/Q vssd1 vssd1 vccd1 vccd1 hold184/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1899__B2 _1912_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout73_A _1918_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold195 _2150_/Q vssd1 vssd1 vccd1 vccd1 hold195/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1339__B1 _1826_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1250_ _1297_/A vssd1 vssd1 vccd1 vccd1 _1336_/A sky130_fd_sc_hd__inv_2
X_1181_ _1745_/A _1149_/Y _1180_/X vssd1 vssd1 vccd1 vccd1 _1181_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_54_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1517_ _1517_/A _1866_/B vssd1 vssd1 vccd1 vccd1 _1517_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_49_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1448_ _1459_/C _1448_/B vssd1 vssd1 vccd1 vccd1 _1829_/B sky130_fd_sc_hd__or2_4
XFILLER_0_4_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1379_ _1331_/X _1776_/A vssd1 vssd1 vccd1 vccd1 _1379_/X sky130_fd_sc_hd__and2b_1
XANTENNA__1805__A1 _2053_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1837__A _1863_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1302_ _1355_/B _2043_/A vssd1 vssd1 vccd1 vccd1 _2015_/D sky130_fd_sc_hd__or2_2
X_1233_ _1233_/A input1/X vssd1 vssd1 vccd1 vccd1 _1233_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_19_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1095_ hold17/X hold21/X _1499_/B vssd1 vssd1 vccd1 vccd1 _1095_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_35_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1164_ hold183/X _1149_/C _1827_/B _1808_/A vssd1 vssd1 vccd1 vccd1 _1164_/X sky130_fd_sc_hd__a22o_1
X_1997_ _1997_/A _1997_/B vssd1 vssd1 vccd1 vccd1 _1997_/X sky130_fd_sc_hd__and2_1
XFILLER_0_42_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1920_ _1920_/A _1920_/B vssd1 vssd1 vccd1 vccd1 _1920_/Y sky130_fd_sc_hd__nand2_4
X_1851_ _1863_/A _1851_/B vssd1 vssd1 vccd1 vccd1 _2144_/D sky130_fd_sc_hd__and2_1
XFILLER_0_8_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1782_ hold98/X _1806_/B vssd1 vssd1 vccd1 vccd1 _1785_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_24_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_87 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2196_ _2206_/CLK _2196_/D vssd1 vssd1 vccd1 vccd1 _2196_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1216_ _1130_/B _1796_/A _1207_/X hold209/X vssd1 vssd1 vccd1 vccd1 _1216_/X sky130_fd_sc_hd__a22o_1
X_1147_ hold195/X _1149_/C _1827_/B _1871_/B vssd1 vssd1 vccd1 vccd1 _1147_/X sky130_fd_sc_hd__a22o_1
X_1078_ _1377_/A _1080_/B vssd1 vssd1 vccd1 vccd1 _1826_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_35_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold11 hold11/A vssd1 vssd1 vccd1 vccd1 hold11/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold22 hold22/A vssd1 vssd1 vccd1 vccd1 hold22/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold55 hold55/A vssd1 vssd1 vccd1 vccd1 hold55/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 hold33/A vssd1 vssd1 vccd1 vccd1 hold33/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 hold44/A vssd1 vssd1 vccd1 vccd1 hold44/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 hold66/A vssd1 vssd1 vccd1 vccd1 hold66/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 hold77/A vssd1 vssd1 vccd1 vccd1 hold77/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 hold88/A vssd1 vssd1 vccd1 vccd1 hold88/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 hold99/A vssd1 vssd1 vccd1 vccd1 hold99/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1935__B1 _2003_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2050_ _2036_/A _2015_/D _2031_/A vssd1 vssd1 vccd1 vccd1 _2050_/Y sky130_fd_sc_hd__o21ai_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1466__A2 _1448_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1218__A2 _1866_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1919__B _1920_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1903_ _1903_/A _1903_/B _1900_/X vssd1 vssd1 vccd1 vccd1 _1903_/X sky130_fd_sc_hd__or3b_1
XFILLER_0_40_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1765_ _2116_/Q _1765_/B vssd1 vssd1 vccd1 vccd1 _1767_/D sky130_fd_sc_hd__nand2_1
X_1834_ hold227/X _1221_/X _1862_/S vssd1 vssd1 vccd1 vccd1 _1835_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_4_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1146__S _1994_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1696_ _1697_/A _1697_/C _1697_/D _1697_/B vssd1 vssd1 vccd1 vccd1 _1696_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_0_4_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2179_ _2219_/CLK _2179_/D vssd1 vssd1 vccd1 vccd1 _2179_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput34 _1446_/X vssd1 vssd1 vccd1 vccd1 io_out[26] sky130_fd_sc_hd__buf_12
XANTENNA_hold200_A _2112_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1845__A _1863_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput23 _1213_/X vssd1 vssd1 vccd1 vccd1 io_out[16] sky130_fd_sc_hd__buf_12
XFILLER_0_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput45 _1166_/X vssd1 vssd1 vccd1 vccd1 io_out[8] sky130_fd_sc_hd__buf_12
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1458__C _1826_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1620__A2 _1776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1550_ hold21/X _1549_/X _1550_/S vssd1 vssd1 vccd1 vccd1 hold22/A sky130_fd_sc_hd__mux2_1
X_1481_ _1030_/Y _2190_/Q _2160_/Q _1480_/Y vssd1 vssd1 vccd1 vccd1 _1481_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_4_9_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _2206_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_34_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2102_ _2225_/CLK hold70/X vssd1 vssd1 vccd1 vccd1 hold69/A sky130_fd_sc_hd__dfxtp_1
X_2033_ _2049_/A _2033_/B vssd1 vssd1 vccd1 vccd1 _2198_/D sky130_fd_sc_hd__and2_1
XTAP_159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1817_ _2117_/Q _1135_/A _1776_/X _2142_/Q _1717_/B vssd1 vssd1 vccd1 vccd1 _1817_/X
+ sky130_fd_sc_hd__a221o_1
X_1748_ _1749_/B _1749_/C _1749_/D _1749_/A vssd1 vssd1 vccd1 vccd1 _1755_/A sky130_fd_sc_hd__a31o_1
XFILLER_0_25_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1679_ _1628_/A _1661_/X _1676_/Y vssd1 vssd1 vccd1 vccd1 _1705_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_63_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1469__B _1826_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1602_ _1650_/B _1606_/A _1650_/A vssd1 vssd1 vccd1 vccd1 _1602_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_22_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1533_ _2115_/Q _1533_/B vssd1 vssd1 vccd1 vccd1 _1534_/B sky130_fd_sc_hd__xor2_1
X_1464_ _2193_/Q _1829_/B _1462_/Y vssd1 vssd1 vccd1 vccd1 _1669_/A sky130_fd_sc_hd__a21o_2
XFILLER_0_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1395_ _1057_/A _1085_/A _1340_/B _1415_/A3 _1907_/S vssd1 vssd1 vccd1 vccd1 _1396_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2016_ _2015_/A _1995_/A _2008_/B _1948_/B _1996_/A vssd1 vssd1 vccd1 vccd1 _2016_/X
+ sky130_fd_sc_hd__o311a_1
XANTENNA__1817__C1 _1717_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1596__B2 _1868_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1379__B _1776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold152 hold245/X vssd1 vssd1 vccd1 vccd1 _1923_/A sky130_fd_sc_hd__buf_1
Xhold174 _2007_/X vssd1 vssd1 vccd1 vccd1 _2190_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold185 _2204_/Q vssd1 vssd1 vccd1 vccd1 _1873_/B sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold163 _2175_/Q vssd1 vssd1 vccd1 vccd1 _2055_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold130 _1750_/X vssd1 vssd1 vccd1 vccd1 _2122_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold141 _2124_/Q vssd1 vssd1 vccd1 vccd1 _1757_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold196 _2205_/Q vssd1 vssd1 vccd1 vccd1 hold196/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1511__A1 _1548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1180_ _2113_/Q _1149_/B _1177_/X _1467_/A _1179_/X vssd1 vssd1 vccd1 vccd1 _1180_/X
+ sky130_fd_sc_hd__a221o_1
X_1516_ _1515_/B _1515_/C _1515_/A vssd1 vssd1 vccd1 vccd1 _1516_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_40_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1447_ _1997_/A _2164_/Q vssd1 vssd1 vccd1 vccd1 _1447_/X sky130_fd_sc_hd__and2_1
XFILLER_0_49_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1378_ _1421_/A _1723_/A _1378_/C _1830_/C vssd1 vssd1 vccd1 vccd1 _1378_/X sky130_fd_sc_hd__or4_1
XFILLER_0_4_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1750__A1 _2053_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1853__A _1863_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1301_ _1355_/C _1995_/B vssd1 vssd1 vccd1 vccd1 _2043_/A sky130_fd_sc_hd__or2_1
X_1232_ input2/X input1/X _1233_/A vssd1 vssd1 vccd1 vccd1 _1232_/X sky130_fd_sc_hd__and3b_2
XFILLER_0_19_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1163_ hold222/X _2096_/Q _1994_/A vssd1 vssd1 vccd1 vccd1 _1808_/A sky130_fd_sc_hd__mux2_4
X_1094_ hold5/X hold45/X _1499_/B vssd1 vssd1 vccd1 vccd1 _1094_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1248__A0 _1796_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1702__S _1920_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1799__A1 _2053_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1996_ _1996_/A _1997_/B _1996_/C vssd1 vssd1 vccd1 vccd1 _1996_/Y sky130_fd_sc_hd__nor3_1
XFILLER_0_51_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_11_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _2201_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_73_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1781_ _2053_/B2 _1785_/A _1780_/Y _1820_/A2 _1775_/A vssd1 vssd1 vccd1 vccd1 _1781_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_29_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1850_ hold201/X _1197_/X _1862_/S vssd1 vssd1 vccd1 vccd1 _1851_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_21_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1146_ hold226/X hold108/X _1994_/A vssd1 vssd1 vccd1 vccd1 _1871_/B sky130_fd_sc_hd__mux2_4
X_2195_ _2208_/CLK _2195_/D vssd1 vssd1 vccd1 vccd1 _2195_/Q sky130_fd_sc_hd__dfxtp_1
X_1215_ hold171/X _1828_/B _1150_/S _1800_/A _1214_/X vssd1 vssd1 vccd1 vccd1 _1215_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_47_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1641__B1 _1864_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1077_ _1345_/A _1144_/B vssd1 vssd1 vccd1 vccd1 _1830_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_70_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1979_ hold79/X _2028_/B _1978_/X _2000_/A vssd1 vssd1 vccd1 vccd1 hold80/A sky130_fd_sc_hd__o211a_1
XFILLER_0_43_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold56 hold56/A vssd1 vssd1 vccd1 vccd1 hold56/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 hold45/A vssd1 vssd1 vccd1 vccd1 hold45/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 hold34/A vssd1 vssd1 vccd1 vccd1 hold34/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 hold23/A vssd1 vssd1 vccd1 vccd1 hold23/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold12 hold12/A vssd1 vssd1 vccd1 vccd1 hold12/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold78 hold78/A vssd1 vssd1 vccd1 vccd1 hold78/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 hold67/A vssd1 vssd1 vccd1 vccd1 hold67/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold89 hold89/A vssd1 vssd1 vccd1 vccd1 hold89/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1935__A1 _1920_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1699__A0 _1239_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1902_ _1901_/X _1866_/B _1907_/S vssd1 vssd1 vccd1 vccd1 _1903_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_29_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1764_ _2149_/Q _1776_/B _1717_/B vssd1 vssd1 vccd1 vccd1 _1767_/C sky130_fd_sc_hd__a21oi_1
XFILLER_0_25_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1833_ _1863_/A _1833_/B vssd1 vssd1 vccd1 vccd1 _2135_/D sky130_fd_sc_hd__and2_1
XFILLER_0_4_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1695_ _1692_/Y _1694_/Y _2188_/Q _1448_/B vssd1 vssd1 vccd1 vccd1 _1695_/X sky130_fd_sc_hd__o211a_1
X_2178_ _2219_/CLK _2178_/D vssd1 vssd1 vccd1 vccd1 _2178_/Q sky130_fd_sc_hd__dfxtp_1
X_1129_ _1776_/A _1129_/B _1229_/B _1827_/A vssd1 vssd1 vccd1 vccd1 _1130_/C sky130_fd_sc_hd__or4_1
XFILLER_0_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput35 _1234_/Y vssd1 vssd1 vccd1 vccd1 io_out[27] sky130_fd_sc_hd__buf_1
XFILLER_0_43_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput24 _1211_/X vssd1 vssd1 vccd1 vccd1 io_out[17] sky130_fd_sc_hd__buf_12
Xoutput46 _1159_/X vssd1 vssd1 vccd1 vccd1 io_out[9] sky130_fd_sc_hd__buf_12
XANTENNA__1861__A _1863_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1480_ _2189_/Q _2185_/Q _1030_/Y vssd1 vssd1 vccd1 vccd1 _1480_/Y sky130_fd_sc_hd__o21ai_1
XTAP_149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2101_ _2225_/CLK hold60/X vssd1 vssd1 vccd1 vccd1 hold59/A sky130_fd_sc_hd__dfxtp_1
X_2032_ _1912_/B _1923_/B _1984_/C _2031_/X vssd1 vssd1 vccd1 vccd1 _2033_/B sky130_fd_sc_hd__a22o_1
XANTENNA__1710__S _1920_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1678_ _1662_/X _1663_/Y _1677_/X _1448_/B _2188_/Q vssd1 vssd1 vccd1 vccd1 _1680_/B
+ sky130_fd_sc_hd__o2111a_1
X_1816_ hold118/X _1820_/A2 _1819_/A _1815_/Y vssd1 vssd1 vccd1 vccd1 _1816_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_32_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1747_ _2113_/Q _1765_/B vssd1 vssd1 vccd1 vccd1 _1749_/D sky130_fd_sc_hd__nand2_1
XFILLER_0_25_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1532_ _1533_/B _2115_/Q vssd1 vssd1 vccd1 vccd1 _1540_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_54_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1601_ _1697_/A _1584_/X _1600_/X vssd1 vssd1 vccd1 vccd1 _1606_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1463_ _2193_/Q _1829_/B _1462_/Y vssd1 vssd1 vccd1 vccd1 _1632_/A sky130_fd_sc_hd__a21oi_4
X_1394_ _1279_/Y _1360_/C _1346_/B _1403_/A2 vssd1 vssd1 vccd1 vccd1 _1413_/B sky130_fd_sc_hd__a22o_1
X_2015_ _2015_/A _2015_/B _2015_/C _2015_/D vssd1 vssd1 vccd1 vccd1 _2015_/Y sky130_fd_sc_hd__nor4_1
XFILLER_0_72_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1596__A2 _1826_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold131 _2183_/Q vssd1 vssd1 vccd1 vccd1 _1239_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold153 _2185_/Q vssd1 vssd1 vccd1 vccd1 hold153/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold120 _2177_/Q vssd1 vssd1 vccd1 vccd1 hold120/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold175 _2110_/Q vssd1 vssd1 vccd1 vccd1 hold175/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold197 _2048_/X vssd1 vssd1 vccd1 vccd1 _2049_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold164 _2055_/X vssd1 vssd1 vccd1 vccd1 hold164/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1826__D _1826_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold142 _1762_/X vssd1 vssd1 vccd1 vccd1 _2124_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold186 _2146_/Q vssd1 vssd1 vccd1 vccd1 hold186/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1511__A2 _1784_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1983__C1 _1871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1515_ _1515_/A _1515_/B _1515_/C vssd1 vssd1 vccd1 vccd1 _1515_/X sky130_fd_sc_hd__and3_1
XFILLER_0_2_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1446_ _1096_/X _1228_/Y _1445_/X vssd1 vssd1 vccd1 vccd1 _1446_/X sky130_fd_sc_hd__a21o_1
X_1377_ _1377_/A _1377_/B vssd1 vssd1 vccd1 vccd1 _1830_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_4_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1170__S _1994_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout70 _2078_/Q vssd1 vssd1 vccd1 vccd1 _1114_/B sky130_fd_sc_hd__buf_4
X_1162_ _1160_/X _1161_/X _1499_/A vssd1 vssd1 vccd1 vccd1 _1162_/X sky130_fd_sc_hd__mux2_1
X_1300_ _1282_/X _1300_/B _1300_/C _1300_/D vssd1 vssd1 vccd1 vccd1 _1311_/A sky130_fd_sc_hd__and4b_1
X_1231_ _1895_/B _1228_/B _1230_/X _2057_/A vssd1 vssd1 vccd1 vccd1 _1231_/Y sky130_fd_sc_hd__o31ai_4
XFILLER_0_19_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1093_ _1174_/B _1174_/C vssd1 vssd1 vccd1 vccd1 _1499_/B sky130_fd_sc_hd__nand2_8
XFILLER_0_47_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1995_ _1995_/A _1995_/B vssd1 vssd1 vccd1 vccd1 _1996_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_51_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1429_ _1193_/X _1228_/Y _1427_/X _1428_/X vssd1 vssd1 vccd1 vccd1 _1429_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_23_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold223_A _1808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1780_ _1780_/A _1780_/B _1780_/C _1780_/D vssd1 vssd1 vccd1 vccd1 _1780_/Y sky130_fd_sc_hd__nand4_1
XFILLER_0_21_12 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1713__S _1920_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2194_ _2206_/CLK hold84/X vssd1 vssd1 vccd1 vccd1 hold83/A sky130_fd_sc_hd__dfxtp_1
X_1145_ _1487_/B _1229_/D vssd1 vssd1 vccd1 vccd1 _1827_/B sky130_fd_sc_hd__or2_4
X_1214_ _1130_/B _1868_/B _1207_/X hold207/X vssd1 vssd1 vccd1 vccd1 _1214_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1076_ _1821_/A _1236_/D _1114_/B _1821_/B vssd1 vssd1 vccd1 vccd1 _1144_/B sky130_fd_sc_hd__nand4_2
XFILLER_0_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1978_ _1978_/A _1978_/B _1977_/X vssd1 vssd1 vccd1 vccd1 _1978_/X sky130_fd_sc_hd__or3b_1
Xhold46 hold46/A vssd1 vssd1 vccd1 vccd1 hold46/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold13 hold13/A vssd1 vssd1 vccd1 vccd1 hold13/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 hold24/A vssd1 vssd1 vccd1 vccd1 hold24/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold68 hold68/A vssd1 vssd1 vccd1 vccd1 hold68/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 hold35/A vssd1 vssd1 vccd1 vccd1 hold35/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold57 hold57/A vssd1 vssd1 vccd1 vccd1 hold57/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 hold79/A vssd1 vssd1 vccd1 vccd1 hold79/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1859__A _1863_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1901_ _1029_/Y _2112_/Q _1901_/S vssd1 vssd1 vccd1 vccd1 _1901_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1832_ hold230/X _1224_/X _1862_/S vssd1 vssd1 vccd1 vccd1 _1832_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_52_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1694_ _1694_/A _1694_/B vssd1 vssd1 vccd1 vccd1 _1694_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_40_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1763_ _1763_/A _1763_/B vssd1 vssd1 vccd1 vccd1 _1767_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_57_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2177_ _2219_/CLK _2177_/D vssd1 vssd1 vccd1 vccd1 _2177_/Q sky130_fd_sc_hd__dfxtp_1
X_1128_ _1128_/A _1487_/A vssd1 vssd1 vccd1 vccd1 _1827_/A sky130_fd_sc_hd__or2_1
X_1059_ _2082_/Q _2081_/Q vssd1 vssd1 vccd1 vccd1 _1127_/A sky130_fd_sc_hd__or2_1
XFILLER_0_28_280 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput25 _1209_/X vssd1 vssd1 vccd1 vccd1 io_out[18] sky130_fd_sc_hd__buf_12
Xoutput36 _2164_/Q vssd1 vssd1 vccd1 vccd1 io_out[2] sky130_fd_sc_hd__buf_12
XFILLER_0_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2100_ _2226_/CLK hold56/X vssd1 vssd1 vccd1 vccd1 hold55/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__1541__A0 _1156_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2031_ _2031_/A _2031_/B vssd1 vssd1 vccd1 vccd1 _2031_/X sky130_fd_sc_hd__and2_1
XFILLER_0_43_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1815_ _1814_/A _1814_/B _2053_/B2 vssd1 vssd1 vccd1 vccd1 _1815_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_0_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1677_ _1662_/A _1662_/B _1676_/Y _1628_/A vssd1 vssd1 vccd1 vccd1 _1677_/X sky130_fd_sc_hd__a211o_1
X_1746_ _2146_/Q _1776_/B _1717_/B vssd1 vssd1 vccd1 vccd1 _1749_/C sky130_fd_sc_hd__a21oi_1
XFILLER_0_4_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1531_ _2108_/Q _1546_/S _1538_/B vssd1 vssd1 vccd1 vccd1 _1533_/B sky130_fd_sc_hd__o21ba_1
X_1600_ _1597_/Y _1598_/X _1599_/X _1654_/A vssd1 vssd1 vccd1 vccd1 _1600_/X sky130_fd_sc_hd__o211a_1
X_1462_ _1922_/B _1462_/B _1829_/B vssd1 vssd1 vccd1 vccd1 _1462_/Y sky130_fd_sc_hd__nor3_2
XFILLER_0_1_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1393_ _1393_/A _1393_/B vssd1 vssd1 vccd1 vccd1 _1401_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_38_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2014_ hold143/X _1923_/B _2013_/X _2003_/A vssd1 vssd1 vccd1 vccd1 _2193_/D sky130_fd_sc_hd__a211o_1
XANTENNA__1817__A1 _2117_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold110 _2130_/Q vssd1 vssd1 vccd1 vccd1 _1794_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold132 _1985_/X vssd1 vssd1 vccd1 vccd1 _2183_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold121 _1959_/X vssd1 vssd1 vccd1 vccd1 _2177_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold154 _2203_/Q vssd1 vssd1 vccd1 vccd1 _1873_/C sky130_fd_sc_hd__dlygate4sd3_1
Xhold143 _2193_/Q vssd1 vssd1 vccd1 vccd1 hold143/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold165 _2056_/Y vssd1 vssd1 vccd1 vccd1 _2057_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold198 _2082_/Q vssd1 vssd1 vccd1 vccd1 _1057_/A sky130_fd_sc_hd__buf_1
X_1729_ _1132_/Y _1732_/B _1728_/B _1035_/Y vssd1 vssd1 vccd1 vccd1 _1729_/X sky130_fd_sc_hd__a211o_1
Xhold187 _1854_/X vssd1 vssd1 vccd1 vccd1 _1855_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold176 _2143_/Q vssd1 vssd1 vccd1 vccd1 hold176/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1541__S _1548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1514_ _2112_/Q _1514_/B vssd1 vssd1 vccd1 vccd1 _1515_/C sky130_fd_sc_hd__or2_1
XFILLER_0_57_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1445_ _2134_/Q _1227_/B _1422_/Y _2117_/Q _1444_/X vssd1 vssd1 vccd1 vccd1 _1445_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_2_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1376_ _1378_/C _2054_/A2 _1282_/X _1360_/C vssd1 vssd1 vccd1 vccd1 _1420_/C sky130_fd_sc_hd__a22o_1
XFILLER_0_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout60 _1243_/Y vssd1 vssd1 vccd1 vccd1 _1820_/A2 sky130_fd_sc_hd__buf_4
Xfanout71 _2077_/Q vssd1 vssd1 vccd1 vccd1 _1821_/B sky130_fd_sc_hd__buf_4
X_1092_ _1174_/B _1174_/C vssd1 vssd1 vccd1 vccd1 _1882_/B sky130_fd_sc_hd__and2_2
X_1161_ hold25/A hold41/A _1499_/B vssd1 vssd1 vccd1 vccd1 _1161_/X sky130_fd_sc_hd__mux2_1
X_1230_ _1238_/A _1238_/B _1229_/X _2183_/Q vssd1 vssd1 vccd1 vccd1 _1230_/X sky130_fd_sc_hd__o31a_1
XFILLER_0_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1994_ _1994_/A _1994_/B vssd1 vssd1 vccd1 vccd1 _1997_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_47_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1428_ hold98/A _1227_/B _1422_/Y _2111_/Q vssd1 vssd1 vccd1 vccd1 _1428_/X sky130_fd_sc_hd__a22o_1
X_1359_ _1288_/Y _1360_/C _1320_/Y _1403_/A2 _1358_/X vssd1 vssd1 vccd1 vccd1 _1413_/A
+ sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_4_2_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1864__B _1864_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1880__A _2057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1883__C1 _1912_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1790__A _1866_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1213_ hold180/X _1828_/B _1150_/S _1806_/A _1212_/X vssd1 vssd1 vccd1 vccd1 _1213_/X
+ sky130_fd_sc_hd__a221o_1
X_2193_ _2208_/CLK _2193_/D vssd1 vssd1 vccd1 vccd1 _2193_/Q sky130_fd_sc_hd__dfxtp_1
X_1075_ _1825_/A _1128_/A _1075_/C _1922_/B vssd1 vssd1 vccd1 vccd1 wire51/A sky130_fd_sc_hd__nor4_1
X_1144_ _1377_/A _1144_/B vssd1 vssd1 vccd1 vccd1 _1229_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_62_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1977_ _2015_/B _1355_/B _2005_/A _1972_/X vssd1 vssd1 vccd1 vccd1 _1977_/X sky130_fd_sc_hd__o31a_1
XANTENNA__2051__C1 _2057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1641__A2 _1776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1157__B2 _1156_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold14 hold14/A vssd1 vssd1 vccd1 vccd1 hold14/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 hold47/A vssd1 vssd1 vccd1 vccd1 hold47/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold69 hold69/A vssd1 vssd1 vccd1 vccd1 hold69/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 hold36/A vssd1 vssd1 vccd1 vccd1 hold36/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 hold25/A vssd1 vssd1 vccd1 vccd1 hold25/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 hold58/A vssd1 vssd1 vccd1 vccd1 hold58/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1935__A3 _1920_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1148__B2 _1545_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1900_ _1029_/A _2199_/Q _1901_/S _1899_/X vssd1 vssd1 vccd1 vccd1 _1900_/X sky130_fd_sc_hd__o31a_1
XFILLER_0_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1831_ _1830_/X _1831_/B vssd1 vssd1 vccd1 vccd1 _1862_/S sky130_fd_sc_hd__and2b_4
XFILLER_0_29_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output15_A _1231_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1693_ _1693_/A _1693_/B _1693_/C vssd1 vssd1 vccd1 vccd1 _1694_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_40_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1762_ _2053_/B2 _1760_/Y _1767_/A _1820_/A2 _1757_/A vssd1 vssd1 vccd1 vccd1 _1762_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_57_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2176_ _2209_/CLK _2176_/D vssd1 vssd1 vccd1 vccd1 _2176_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1058_ _1089_/B _1225_/B vssd1 vssd1 vccd1 vccd1 _1467_/A sky130_fd_sc_hd__nand2_4
X_1127_ _1127_/A _1144_/B vssd1 vssd1 vccd1 vccd1 _1487_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_28_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput37 _2163_/Q vssd1 vssd1 vccd1 vccd1 io_out[31] sky130_fd_sc_hd__buf_12
Xoutput26 _1426_/X vssd1 vssd1 vccd1 vccd1 io_out[19] sky130_fd_sc_hd__buf_12
Xoutput15 _1231_/Y vssd1 vssd1 vccd1 vccd1 io_oeb sky130_fd_sc_hd__buf_12
XFILLER_0_11_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2030_ _2036_/A _2030_/B vssd1 vssd1 vccd1 vccd1 _2031_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_43_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1814_ _1814_/A _1814_/B vssd1 vssd1 vccd1 vccd1 _1819_/A sky130_fd_sc_hd__or2_1
X_1745_ _1745_/A _1763_/B vssd1 vssd1 vccd1 vccd1 _1749_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_68_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1676_ _1680_/A _1676_/B vssd1 vssd1 vccd1 vccd1 _1676_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_40_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2159_ _2214_/CLK _2159_/D vssd1 vssd1 vccd1 vccd1 _2159_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1530_ _2188_/Q _2108_/Q _2151_/Q vssd1 vssd1 vccd1 vccd1 _1538_/B sky130_fd_sc_hd__and3_1
X_1461_ _2126_/Q _1826_/D _1460_/Y _1871_/B vssd1 vssd1 vccd1 vccd1 _1492_/A sky130_fd_sc_hd__a22o_1
X_1392_ _1392_/A _1392_/B vssd1 vssd1 vccd1 vccd1 _2079_/D sky130_fd_sc_hd__or2_1
XFILLER_0_1_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1762__A1 _2053_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2013_ _1995_/A _1355_/C _1996_/A _2028_/B vssd1 vssd1 vccd1 vccd1 _2013_/X sky130_fd_sc_hd__o31a_1
XANTENNA__1817__A2 _1135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_7_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold144 _2198_/Q vssd1 vssd1 vccd1 vccd1 _1912_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold122 _2196_/Q vssd1 vssd1 vccd1 vccd1 _1450_/A sky130_fd_sc_hd__buf_1
Xhold100 _2127_/Q vssd1 vssd1 vccd1 vccd1 _1775_/A sky130_fd_sc_hd__buf_1
Xhold111 _1799_/X vssd1 vssd1 vccd1 vccd1 _2130_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1728_ _1732_/A _1728_/B vssd1 vssd1 vccd1 vccd1 _1728_/Y sky130_fd_sc_hd__nand2_1
Xhold133 _2121_/Q vssd1 vssd1 vccd1 vccd1 hold133/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold177 _2111_/Q vssd1 vssd1 vccd1 vccd1 hold177/X sky130_fd_sc_hd__buf_1
X_1659_ _1639_/X _1659_/B vssd1 vssd1 vccd1 vccd1 _1663_/B sky130_fd_sc_hd__nand2b_1
Xhold188 _2201_/Q vssd1 vssd1 vccd1 vccd1 hold188/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold155 _2044_/X vssd1 vssd1 vccd1 vccd1 _2045_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold166 _2206_/Q vssd1 vssd1 vccd1 vccd1 _1912_/A sky130_fd_sc_hd__clkbuf_4
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold199 _1225_/B vssd1 vssd1 vccd1 vccd1 _1456_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_8_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _2210_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_63_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1744__A1 _1922_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1496__C _1922_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1513_ _2112_/Q _1514_/B vssd1 vssd1 vccd1 vccd1 _1515_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_49_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1444_ _2126_/Q _1441_/B _1423_/X _2162_/Q vssd1 vssd1 vccd1 vccd1 _1444_/X sky130_fd_sc_hd__a22o_1
X_1375_ _1375_/A _1402_/B _1402_/C vssd1 vssd1 vccd1 vccd1 _2078_/D sky130_fd_sc_hd__or3_1
XFILLER_0_4_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout72 _1243_/B vssd1 vssd1 vccd1 vccd1 _2003_/A sky130_fd_sc_hd__clkbuf_8
Xfanout50 _2031_/A vssd1 vssd1 vccd1 vccd1 _2028_/B sky130_fd_sc_hd__buf_4
Xfanout61 _1365_/A vssd1 vssd1 vccd1 vccd1 _1415_/A3 sky130_fd_sc_hd__buf_4
XFILLER_0_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1160_ hold31/A hold23/A _1499_/B vssd1 vssd1 vccd1 vccd1 _1160_/X sky130_fd_sc_hd__mux2_1
X_1091_ _2182_/Q _1467_/B wire51/X _1090_/X vssd1 vssd1 vccd1 vccd1 _1174_/C sky130_fd_sc_hd__a211o_4
XFILLER_0_55_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1993_ _2049_/A _1993_/B vssd1 vssd1 vccd1 vccd1 _2186_/D sky130_fd_sc_hd__and2_1
XFILLER_0_27_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1427_ _2120_/Q _1441_/B _1423_/X _2161_/Q vssd1 vssd1 vccd1 vccd1 _1427_/X sky130_fd_sc_hd__a22o_1
X_1358_ _1903_/B _1723_/B _1415_/A3 vssd1 vssd1 vccd1 vccd1 _1358_/X sky130_fd_sc_hd__o21a_1
X_1289_ _1306_/A _1306_/B vssd1 vssd1 vccd1 vccd1 _1984_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_38_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2192_ _2201_/CLK _2192_/D vssd1 vssd1 vccd1 vccd1 _2192_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1212_ _1130_/B _1808_/A _1207_/X hold211/X vssd1 vssd1 vccd1 vccd1 _1212_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_20_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1143_ _1143_/A _1345_/A vssd1 vssd1 vccd1 vccd1 _1487_/B sky130_fd_sc_hd__nor2_1
X_1074_ _1344_/A _1080_/B vssd1 vssd1 vccd1 vccd1 _1921_/B sky130_fd_sc_hd__or2_4
XFILLER_0_1_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1976_ _1980_/A _1306_/A _2015_/C _1984_/C _1923_/B vssd1 vssd1 vccd1 vccd1 _1978_/B
+ sky130_fd_sc_hd__a41o_1
XFILLER_0_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold48 hold48/A vssd1 vssd1 vccd1 vccd1 hold48/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 hold26/A vssd1 vssd1 vccd1 vccd1 hold26/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold15 hold15/A vssd1 vssd1 vccd1 vccd1 hold15/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 hold37/A vssd1 vssd1 vccd1 vccd1 hold37/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 hold59/A vssd1 vssd1 vccd1 vccd1 hold59/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1830_ _1921_/A _1830_/B _1830_/C _1920_/B vssd1 vssd1 vccd1 vccd1 _1830_/X sky130_fd_sc_hd__or4_1
X_1761_ _1760_/B _1760_/C _1760_/D _1760_/A vssd1 vssd1 vccd1 vccd1 _1767_/A sky130_fd_sc_hd__a31o_1
X_1692_ _1693_/B _1692_/B vssd1 vssd1 vccd1 vccd1 _1692_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_73_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_10_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _1233_/A sky130_fd_sc_hd__clkbuf_8
X_2175_ _1233_/A _2175_/D vssd1 vssd1 vccd1 vccd1 _2175_/Q sky130_fd_sc_hd__dfxtp_1
X_1126_ _1126_/A _1335_/B vssd1 vssd1 vccd1 vccd1 _1229_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_73_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1057_ _1057_/A _2081_/Q _1345_/B vssd1 vssd1 vccd1 vccd1 _1225_/B sky130_fd_sc_hd__or3_4
XANTENNA__1187__S _1994_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1959_ hold120/X _2028_/B _1978_/A _1958_/X _2000_/A vssd1 vssd1 vccd1 vccd1 _1959_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA__1783__C1 _1717_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput38 _2165_/Q vssd1 vssd1 vccd1 vccd1 io_out[32] sky130_fd_sc_hd__buf_12
Xoutput27 _2161_/Q vssd1 vssd1 vccd1 vccd1 io_out[1] sky130_fd_sc_hd__buf_12
XFILLER_0_3_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput16 _2160_/Q vssd1 vssd1 vccd1 vccd1 io_out[0] sky130_fd_sc_hd__buf_12
XFILLER_0_11_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2047__A _2057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1796__A _1796_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1813_ _1156_/X _1808_/B _1806_/B hold118/X _1812_/X vssd1 vssd1 vccd1 vccd1 _1814_/B
+ sky130_fd_sc_hd__a221oi_2
X_1744_ _1922_/B _1765_/B _1724_/C vssd1 vssd1 vccd1 vccd1 _1763_/B sky130_fd_sc_hd__o21bai_4
XFILLER_0_25_241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1675_ _1674_/B _1674_/C _1674_/A vssd1 vssd1 vccd1 vccd1 _1676_/B sky130_fd_sc_hd__a21oi_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2158_ _2182_/CLK _2158_/D vssd1 vssd1 vccd1 vccd1 _2158_/Q sky130_fd_sc_hd__dfxtp_1
X_2089_ _2225_/CLK hold68/X vssd1 vssd1 vccd1 vccd1 hold67/A sky130_fd_sc_hd__dfxtp_1
X_1109_ _2082_/Q _1085_/A _1079_/X vssd1 vssd1 vccd1 vccd1 _1110_/D sky130_fd_sc_hd__a21bo_1
XFILLER_0_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1460_ _1460_/A _1825_/C _1460_/C _1460_/D vssd1 vssd1 vccd1 vccd1 _1460_/Y sky130_fd_sc_hd__nor4_4
X_1391_ _1391_/A _1391_/B _1401_/A _1391_/D vssd1 vssd1 vccd1 vccd1 _1392_/B sky130_fd_sc_hd__or4_1
XFILLER_0_1_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2012_ _2049_/A _2012_/B vssd1 vssd1 vccd1 vccd1 _2192_/D sky130_fd_sc_hd__and2_1
XFILLER_0_72_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold156 hold244/X vssd1 vssd1 vccd1 vccd1 _1874_/B sky130_fd_sc_hd__buf_1
Xhold145 _2186_/Q vssd1 vssd1 vccd1 vccd1 hold145/X sky130_fd_sc_hd__dlygate4sd3_1
X_1658_ _1639_/B _1639_/C _1639_/A vssd1 vssd1 vccd1 vccd1 _1659_/B sky130_fd_sc_hd__a21o_1
Xhold123 _2027_/X vssd1 vssd1 vccd1 vccd1 _2196_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold167 _2163_/Q vssd1 vssd1 vccd1 vccd1 hold167/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold112 _2132_/Q vssd1 vssd1 vccd1 vccd1 _1806_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold101 _1781_/X vssd1 vssd1 vccd1 vccd1 _2127_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1727_ _1735_/A _1734_/A _1726_/X _1820_/A2 hold139/X vssd1 vssd1 vccd1 vccd1 _1727_/X
+ sky130_fd_sc_hd__a32o_1
Xhold134 _1743_/X vssd1 vssd1 vccd1 vccd1 _2121_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold189 _2039_/X vssd1 vssd1 vccd1 vccd1 _2040_/B sky130_fd_sc_hd__dlygate4sd3_1
X_1589_ _1586_/Y _1587_/X _1588_/X _1654_/A vssd1 vssd1 vccd1 vccd1 _1589_/X sky130_fd_sc_hd__o211a_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold178 _2149_/Q vssd1 vssd1 vccd1 vccd1 hold178/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1512_ hold9/X _1511_/X _1550_/S vssd1 vssd1 vccd1 vccd1 hold10/A sky130_fd_sc_hd__mux2_1
XFILLER_0_35_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1374_ _1299_/A _1393_/A _1373_/Y vssd1 vssd1 vccd1 vccd1 _1402_/C sky130_fd_sc_hd__o21ai_1
X_1443_ _1155_/Y _1228_/Y _1422_/Y _2116_/Q _1442_/X vssd1 vssd1 vccd1 vccd1 _1443_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_58_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout62 _1296_/B vssd1 vssd1 vccd1 vccd1 _1365_/A sky130_fd_sc_hd__clkbuf_4
Xfanout73 _1918_/A vssd1 vssd1 vccd1 vccd1 _1863_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_36 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output38_A _2165_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1090_ _2178_/Q _1922_/B vssd1 vssd1 vccd1 vccd1 _1090_/X sky130_fd_sc_hd__and2_1
XFILLER_0_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1992_ hold145/X _2043_/B _1990_/Y _1991_/X vssd1 vssd1 vccd1 vccd1 _1992_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_51_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1288_ _1300_/B vssd1 vssd1 vccd1 vccd1 _1288_/Y sky130_fd_sc_hd__inv_2
X_1426_ _1202_/Y _1228_/Y _1424_/X _1425_/X vssd1 vssd1 vccd1 vccd1 _1426_/X sky130_fd_sc_hd__a211o_1
X_1357_ _1417_/B _1412_/B vssd1 vssd1 vccd1 vccd1 _1408_/B sky130_fd_sc_hd__or2_1
XFILLER_0_65_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1644__B2 _1864_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1129__A _1776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2191_ _2206_/CLK _2191_/D vssd1 vssd1 vccd1 vccd1 _2191_/Q sky130_fd_sc_hd__dfxtp_1
X_1211_ hold193/X _1828_/B _1150_/S hold118/X _1210_/X vssd1 vssd1 vccd1 vccd1 _1211_/X
+ sky130_fd_sc_hd__a221o_1
X_1142_ _1828_/B _1459_/C _1895_/B vssd1 vssd1 vccd1 vccd1 _1149_/C sky130_fd_sc_hd__or3_4
X_1073_ _1344_/A _1080_/B vssd1 vssd1 vccd1 vccd1 _1881_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_1_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1975_ hold61/X _1923_/B _1974_/Y _2003_/A vssd1 vssd1 vccd1 vccd1 hold62/A sky130_fd_sc_hd__a211o_1
XANTENNA__2051__A1 _1912_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1039__A _1039_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold27 hold27/A vssd1 vssd1 vccd1 vccd1 hold27/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold16 hold16/A vssd1 vssd1 vccd1 vccd1 hold16/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold38 hold38/A vssd1 vssd1 vccd1 vccd1 hold38/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1409_ _1409_/A _1409_/B _1402_/X vssd1 vssd1 vccd1 vccd1 _2080_/D sky130_fd_sc_hd__or3b_1
Xhold49 hold49/A vssd1 vssd1 vccd1 vccd1 hold49/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1502__A _1548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1691_ _1691_/A _1708_/B _1691_/C vssd1 vssd1 vccd1 vccd1 _1692_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_44_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1760_ _1760_/A _1760_/B _1760_/C _1760_/D vssd1 vssd1 vccd1 vccd1 _1760_/Y sky130_fd_sc_hd__nand4_1
XFILLER_0_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2174_ _2214_/CLK hold8/X vssd1 vssd1 vccd1 vccd1 hold7/A sky130_fd_sc_hd__dfxtp_1
X_1125_ _1345_/A _1377_/B vssd1 vssd1 vccd1 vccd1 _1129_/B sky130_fd_sc_hd__nor2_1
X_1056_ _2081_/Q _1345_/B vssd1 vssd1 vccd1 vccd1 _1085_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_28_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput39 _2162_/Q vssd1 vssd1 vccd1 vccd1 io_out[33] sky130_fd_sc_hd__buf_12
X_1958_ _1255_/Y _2001_/C _1957_/X _1955_/X vssd1 vssd1 vccd1 vccd1 _1958_/X sky130_fd_sc_hd__a31o_1
X_1889_ _2115_/Q _2116_/Q _2114_/Q _2113_/Q vssd1 vssd1 vccd1 vccd1 _1889_/X sky130_fd_sc_hd__or4_1
Xoutput28 _1429_/X vssd1 vssd1 vccd1 vccd1 io_out[20] sky130_fd_sc_hd__buf_12
XFILLER_0_43_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput17 _1150_/X vssd1 vssd1 vccd1 vccd1 io_out[10] sky130_fd_sc_hd__buf_12
XFILLER_0_11_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1674_ _1674_/A _1674_/B _1674_/C vssd1 vssd1 vccd1 vccd1 _1680_/A sky130_fd_sc_hd__and3_1
X_1812_ _2116_/Q _1135_/A _1776_/X _2141_/Q _1717_/B vssd1 vssd1 vccd1 vccd1 _1812_/X
+ sky130_fd_sc_hd__a221o_1
X_1743_ _2053_/B2 _1749_/A _1742_/Y _1820_/A2 hold133/X vssd1 vssd1 vccd1 vccd1 _1743_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_25_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2226_ _2226_/CLK hold18/X vssd1 vssd1 vccd1 vccd1 hold17/A sky130_fd_sc_hd__dfxtp_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2157_ _2172_/CLK _2157_/D vssd1 vssd1 vccd1 vccd1 _2157_/Q sky130_fd_sc_hd__dfxtp_1
X_2088_ _2226_/CLK hold42/X vssd1 vssd1 vccd1 vccd1 hold41/A sky130_fd_sc_hd__dfxtp_1
X_1039_ _1039_/A vssd1 vssd1 vccd1 vccd1 _1039_/Y sky130_fd_sc_hd__inv_2
X_1108_ _1377_/A _1320_/B vssd1 vssd1 vccd1 vccd1 _1486_/D sky130_fd_sc_hd__nor2_2
XFILLER_0_48_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1220__A2 _1865_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1836__S _1862_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1390_ _1390_/A _1390_/B _1390_/C _1404_/A vssd1 vssd1 vccd1 vccd1 _1391_/D sky130_fd_sc_hd__or4_1
XFILLER_0_22_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2011_ hold203/X _2043_/B _2001_/X _1995_/A vssd1 vssd1 vccd1 vccd1 _2012_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_72_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold102 _2093_/Q vssd1 vssd1 vccd1 vccd1 hold102/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold124 _2178_/Q vssd1 vssd1 vccd1 vccd1 _1965_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold157 _2197_/Q vssd1 vssd1 vccd1 vccd1 _2028_/A sky130_fd_sc_hd__dlygate4sd3_1
X_1657_ _1701_/A _1656_/B _1653_/Y vssd1 vssd1 vccd1 vccd1 _1663_/A sky130_fd_sc_hd__a21o_1
Xhold146 _1992_/X vssd1 vssd1 vccd1 vccd1 _1993_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 _1904_/X vssd1 vssd1 vccd1 vccd1 _2163_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1588_ _1632_/A _1592_/S _1584_/X vssd1 vssd1 vccd1 vccd1 _1588_/X sky130_fd_sc_hd__a21o_1
Xhold113 _1811_/X vssd1 vssd1 vccd1 vccd1 _2132_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1726_ _1726_/A _1726_/B _1726_/C vssd1 vssd1 vccd1 vccd1 _1726_/X sky130_fd_sc_hd__or3_1
Xhold135 _2120_/Q vssd1 vssd1 vccd1 vccd1 _1732_/A sky130_fd_sc_hd__buf_1
Xhold179 _1860_/X vssd1 vssd1 vccd1 vccd1 _1861_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2209_ _2209_/CLK hold82/X vssd1 vssd1 vccd1 vccd1 hold81/A sky130_fd_sc_hd__dfxtp_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1729__B1 _1728_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_11_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1511_ _1548_/A _1784_/A _1542_/A _1510_/Y vssd1 vssd1 vccd1 vccd1 _1511_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_50_384 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1442_ _2133_/Q _1227_/B _1423_/X _2165_/Q _1441_/X vssd1 vssd1 vccd1 vccd1 _1442_/X
+ sky130_fd_sc_hd__a221o_1
X_1373_ _1062_/Y _1373_/A2 _1405_/B _1417_/C _1411_/B vssd1 vssd1 vccd1 vccd1 _1373_/Y
+ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_73_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1709_ _1708_/X _1707_/Y hold171/X _1921_/A vssd1 vssd1 vccd1 vccd1 _1709_/X sky130_fd_sc_hd__a2bb2o_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout74 _1871_/A vssd1 vssd1 vccd1 vccd1 _2000_/A sky130_fd_sc_hd__buf_4
Xfanout63 _2053_/B2 vssd1 vssd1 vccd1 vccd1 _1296_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_0_36_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout52 _1284_/A vssd1 vssd1 vccd1 vccd1 _1728_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_24_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1991_ _1980_/A _1995_/A _2001_/C _1955_/B vssd1 vssd1 vccd1 vccd1 _1991_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1425_ _2119_/Q _1441_/B _1422_/Y _2110_/Q vssd1 vssd1 vccd1 vccd1 _1425_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_2_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1287_ _2008_/A _1287_/B _1947_/A vssd1 vssd1 vccd1 vccd1 _1300_/B sky130_fd_sc_hd__or3_1
X_1356_ _1486_/A _1373_/A2 _1355_/X vssd1 vssd1 vccd1 vccd1 _1412_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_65_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1644__A2 _1826_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1801__C1 _1717_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1235__A _1921_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1332__B2 _1135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1332__A1 _1776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1844__S _1862_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2190_ _2219_/CLK _2190_/D vssd1 vssd1 vccd1 vccd1 _2190_/Q sky130_fd_sc_hd__dfxtp_1
X_1141_ _1377_/A _1141_/B vssd1 vssd1 vccd1 vccd1 _1141_/X sky130_fd_sc_hd__or2_2
X_1210_ _1130_/B _1156_/X _1207_/X hold206/X vssd1 vssd1 vccd1 vccd1 _1210_/X sky130_fd_sc_hd__a22o_1
X_1072_ _1114_/B _1821_/B _1821_/A _1236_/D vssd1 vssd1 vccd1 vccd1 _1080_/B sky130_fd_sc_hd__or4bb_4
XFILLER_0_1_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1974_ _1972_/X _1973_/X _2043_/B vssd1 vssd1 vccd1 vccd1 _1974_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_47_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold17 hold17/A vssd1 vssd1 vccd1 vccd1 hold17/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold28 hold28/A vssd1 vssd1 vccd1 vccd1 hold28/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold39 hold39/A vssd1 vssd1 vccd1 vccd1 hold39/X sky130_fd_sc_hd__dlygate4sd3_1
X_1408_ _1408_/A _1408_/B _1408_/C _1408_/D vssd1 vssd1 vccd1 vccd1 _1409_/B sky130_fd_sc_hd__or4_1
XANTENNA__1502__B _1864_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1339_ _1960_/B _1313_/Y _1826_/D _1373_/A2 vssd1 vssd1 vccd1 vccd1 _1390_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_46_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold214_A _2164_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1690_ _1697_/D _1690_/B vssd1 vssd1 vccd1 vccd1 _1690_/X sky130_fd_sc_hd__and2_1
XFILLER_0_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2173_ _2182_/CLK hold54/X vssd1 vssd1 vccd1 vccd1 hold53/A sky130_fd_sc_hd__dfxtp_1
X_1124_ _1344_/A _1320_/B vssd1 vssd1 vccd1 vccd1 _1716_/B sky130_fd_sc_hd__nor2_2
X_1055_ _1236_/D _1114_/B _1821_/B _1821_/A vssd1 vssd1 vccd1 vccd1 _1345_/B sky130_fd_sc_hd__or4b_2
X_1957_ _1973_/A _2030_/B _2001_/A _1285_/B vssd1 vssd1 vccd1 vccd1 _1957_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_28_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1535__A1 _1548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput29 _1432_/X vssd1 vssd1 vccd1 vccd1 io_out[21] sky130_fd_sc_hd__buf_12
X_1888_ _2112_/Q _2111_/Q _2110_/Q _2117_/Q vssd1 vssd1 vccd1 vccd1 _1888_/X sky130_fd_sc_hd__or4_1
XFILLER_0_43_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput18 _1224_/X vssd1 vssd1 vccd1 vccd1 io_out[11] sky130_fd_sc_hd__buf_12
XANTENNA__1513__A _2112_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1811_ _2053_/B2 _1809_/Y _1814_/A _1820_/A2 _1806_/A vssd1 vssd1 vccd1 vccd1 _1811_/X
+ sky130_fd_sc_hd__a32o_1
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1673_ _1651_/A _1491_/B _1673_/S vssd1 vssd1 vccd1 vccd1 _1674_/C sky130_fd_sc_hd__mux2_1
X_1742_ _1742_/A _1742_/B _1742_/C _1742_/D vssd1 vssd1 vccd1 vccd1 _1742_/Y sky130_fd_sc_hd__nand4_1
XFILLER_0_25_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2225_ _2225_/CLK hold48/X vssd1 vssd1 vccd1 vccd1 hold47/A sky130_fd_sc_hd__dfxtp_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1038_ _2000_/A vssd1 vssd1 vccd1 vccd1 _1243_/B sky130_fd_sc_hd__inv_2
X_2156_ _2182_/CLK _2156_/D vssd1 vssd1 vccd1 vccd1 _2156_/Q sky130_fd_sc_hd__dfxtp_1
X_2087_ _2223_/CLK hold52/X vssd1 vssd1 vccd1 vccd1 hold51/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1107_ _1821_/A _1821_/B _1114_/B _1236_/D vssd1 vssd1 vccd1 vccd1 _1320_/B sky130_fd_sc_hd__or4bb_2
XFILLER_0_8_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1756__A1 _2053_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1243__A _1994_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2010_ _1923_/B _2008_/Y _2009_/X _2000_/A vssd1 vssd1 vccd1 vccd1 _2010_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_38_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1852__S _1862_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1725_ _1726_/A _1726_/B _1726_/C vssd1 vssd1 vccd1 vccd1 _1734_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__1738__A1 _1025_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold103 _1930_/X vssd1 vssd1 vccd1 vccd1 _2169_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold158 _2029_/X vssd1 vssd1 vccd1 vccd1 _2197_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold169 _2191_/Q vssd1 vssd1 vccd1 vccd1 _2009_/A sky130_fd_sc_hd__buf_1
Xhold114 _2187_/Q vssd1 vssd1 vccd1 vccd1 _1997_/A sky130_fd_sc_hd__buf_1
X_1656_ _1653_/Y _1656_/B vssd1 vssd1 vccd1 vccd1 _1701_/B sky130_fd_sc_hd__nand2b_1
Xhold147 _2161_/Q vssd1 vssd1 vccd1 vccd1 hold147/X sky130_fd_sc_hd__dlygate4sd3_1
X_1587_ _1476_/C _1584_/X _1592_/S _1475_/Y vssd1 vssd1 vccd1 vccd1 _1587_/X sky130_fd_sc_hd__a31o_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold125 _2126_/Q vssd1 vssd1 vccd1 vccd1 hold125/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold136 _1736_/X vssd1 vssd1 vccd1 vccd1 _2120_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2208_ _2208_/CLK hold74/X vssd1 vssd1 vccd1 vccd1 hold73/A sky130_fd_sc_hd__dfxtp_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2139_ _2142_/CLK _2139_/D vssd1 vssd1 vccd1 vccd1 _2139_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1901__A1 _2112_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1510_ _1515_/A _1509_/Y _1548_/A vssd1 vssd1 vccd1 vccd1 _1510_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_50_396 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1441_ _2125_/Q _1441_/B vssd1 vssd1 vccd1 vccd1 _1441_/X sky130_fd_sc_hd__and2_1
XFILLER_0_65_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1372_ _1487_/B _1373_/A2 _1960_/B _1360_/X vssd1 vssd1 vccd1 vccd1 _1411_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_73_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1708_ _1921_/A _1708_/B vssd1 vssd1 vccd1 vccd1 _1708_/X sky130_fd_sc_hd__or2_1
X_1639_ _1639_/A _1639_/B _1639_/C vssd1 vssd1 vccd1 vccd1 _1639_/X sky130_fd_sc_hd__and3_1
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout75 _1871_/A vssd1 vssd1 vccd1 vccd1 _2049_/A sky130_fd_sc_hd__clkbuf_4
Xfanout64 _1735_/A vssd1 vssd1 vccd1 vccd1 _2053_/B2 sky130_fd_sc_hd__buf_4
Xfanout53 _1716_/B vssd1 vssd1 vccd1 vccd1 _1776_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_32_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1990_ _2043_/B _2005_/A vssd1 vssd1 vccd1 vccd1 _1990_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_42_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_7_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _2225_/CLK sky130_fd_sc_hd__clkbuf_8
X_1355_ _2036_/A _1355_/B _1355_/C _1393_/A vssd1 vssd1 vccd1 vccd1 _1355_/X sky130_fd_sc_hd__or4_1
X_1424_ _2127_/Q _1227_/B _1423_/X _2160_/Q vssd1 vssd1 vccd1 vccd1 _1424_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_23_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1286_ _2008_/A _1947_/A vssd1 vssd1 vccd1 vccd1 _1286_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__1629__B1 _1784_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1235__B _2003_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1071_ _1821_/A _1236_/D vssd1 vssd1 vccd1 vccd1 _1071_/Y sky130_fd_sc_hd__nand2_1
X_1140_ _1377_/A _1141_/B vssd1 vssd1 vccd1 vccd1 _1895_/B sky130_fd_sc_hd__nor2_8
XFILLER_0_1_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1860__S _1862_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1973_ _1973_/A _1973_/B _2030_/B vssd1 vssd1 vccd1 vccd1 _1973_/X sky130_fd_sc_hd__or3_1
XFILLER_0_28_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1795__C1 _1717_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold29 hold29/A vssd1 vssd1 vccd1 vccd1 hold29/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold18 hold18/A vssd1 vssd1 vccd1 vccd1 hold18/X sky130_fd_sc_hd__dlygate4sd3_1
X_1338_ _1338_/A _1344_/A vssd1 vssd1 vccd1 vccd1 _1826_/D sky130_fd_sc_hd__nor2_8
X_1407_ _1407_/A _1407_/B _1407_/C _1407_/D vssd1 vssd1 vccd1 vccd1 _1408_/D sky130_fd_sc_hd__or4_1
X_1269_ _1728_/B _1945_/A vssd1 vssd1 vccd1 vccd1 _1355_/C sky130_fd_sc_hd__and2_2
XFILLER_0_36_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1777__C1 _1717_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2172_ _2172_/CLK hold28/X vssd1 vssd1 vccd1 vccd1 hold27/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1054_ _1421_/A _1548_/A _1054_/C vssd1 vssd1 vccd1 vccd1 _1089_/B sky130_fd_sc_hd__and3b_2
X_1123_ _1123_/A _1828_/A _1123_/C vssd1 vssd1 vccd1 vccd1 _1130_/B sky130_fd_sc_hd__or3_4
X_1956_ _1980_/B _1995_/A vssd1 vssd1 vccd1 vccd1 _2030_/B sky130_fd_sc_hd__nand2_1
X_1887_ _2206_/Q _1907_/S _1141_/X vssd1 vssd1 vccd1 vccd1 _1887_/X sky130_fd_sc_hd__o21a_1
XANTENNA__1783__A2 _1135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1535__A2 _1808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput19 _1221_/X vssd1 vssd1 vccd1 vccd1 io_out[12] sky130_fd_sc_hd__buf_12
XFILLER_0_3_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1471__A1 _2117_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1810_ _1809_/B _1809_/C _1809_/D _1809_/A vssd1 vssd1 vccd1 vccd1 _1814_/A sky130_fd_sc_hd__a31o_1
X_1741_ _1742_/B _1742_/C _1742_/D _1742_/A vssd1 vssd1 vccd1 vccd1 _1749_/A sky130_fd_sc_hd__a31o_1
XFILLER_0_25_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1672_ _1491_/B _1674_/A _1491_/A vssd1 vssd1 vccd1 vccd1 _1674_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_7_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2155_ _2172_/CLK _2155_/D vssd1 vssd1 vccd1 vccd1 _2155_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2224_ _2226_/CLK hold26/X vssd1 vssd1 vccd1 vccd1 hold25/A sky130_fd_sc_hd__dfxtp_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1106_ _1106_/A _1344_/A vssd1 vssd1 vccd1 vccd1 _1455_/B sky130_fd_sc_hd__nor2_2
X_2086_ _2225_/CLK hold44/X vssd1 vssd1 vccd1 vccd1 hold43/A sky130_fd_sc_hd__dfxtp_1
X_1037_ _2081_/Q vssd1 vssd1 vccd1 vccd1 _1245_/B sky130_fd_sc_hd__inv_2
XFILLER_0_8_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1939_ _1994_/A _2098_/Q _1920_/B _2003_/A vssd1 vssd1 vccd1 vccd1 _1939_/X sky130_fd_sc_hd__a31o_1
XANTENNA__1495__S _1920_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1444__B2 _2162_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1904__C1 _2057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1380__B1 _1448_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold115 _1447_/X vssd1 vssd1 vccd1 vccd1 _2151_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold104 _2129_/Q vssd1 vssd1 vccd1 vccd1 _1788_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold126 _1773_/X vssd1 vssd1 vccd1 vccd1 _2126_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1724_ _1724_/A _1724_/B _1724_/C _1724_/D vssd1 vssd1 vccd1 vccd1 _1726_/C sky130_fd_sc_hd__or4_1
XFILLER_0_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold159 _2195_/Q vssd1 vssd1 vccd1 vccd1 hold159/X sky130_fd_sc_hd__dlygate4sd3_1
X_1655_ _1650_/A _1653_/B _1653_/A vssd1 vssd1 vccd1 vccd1 _1656_/B sky130_fd_sc_hd__o21ai_1
Xhold148 _1892_/X vssd1 vssd1 vccd1 vccd1 _2161_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1586_ _1584_/X _1592_/S _1669_/A vssd1 vssd1 vccd1 vccd1 _1586_/Y sky130_fd_sc_hd__a21oi_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold137 _2123_/Q vssd1 vssd1 vccd1 vccd1 _1751_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2069_ hold57/X _1511_/X _2075_/S vssd1 vssd1 vccd1 vccd1 hold58/A sky130_fd_sc_hd__mux2_1
X_2207_ _2208_/CLK hold88/X vssd1 vssd1 vccd1 vccd1 hold87/A sky130_fd_sc_hd__dfxtp_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2138_ _2150_/CLK _2138_/D vssd1 vssd1 vccd1 vccd1 _2138_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1362__A0 _2162_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1440_ _2132_/Q _1227_/B _1228_/Y _1162_/X _1439_/X vssd1 vssd1 vccd1 vccd1 _1440_/X
+ sky130_fd_sc_hd__a221o_1
X_1371_ _1421_/A _1373_/A2 _1465_/B _1296_/B vssd1 vssd1 vccd1 vccd1 _1417_/C sky130_fd_sc_hd__a22o_1
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1707_ _1707_/A _1707_/B vssd1 vssd1 vccd1 vccd1 _1707_/Y sky130_fd_sc_hd__nor2_1
X_1638_ _1491_/B _1651_/A _1638_/S vssd1 vssd1 vccd1 vccd1 _1639_/C sky130_fd_sc_hd__mux2_1
XFILLER_0_41_364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1569_ _1570_/A _1570_/B vssd1 vssd1 vccd1 vccd1 _1697_/B sky130_fd_sc_hd__or2_1
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1802__A _1868_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1249__A _1728_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout76 _2057_/A vssd1 vssd1 vccd1 vccd1 _1871_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_36_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout65 _1127_/A vssd1 vssd1 vccd1 vccd1 _1344_/A sky130_fd_sc_hd__buf_8
Xfanout54 _1455_/B vssd1 vssd1 vccd1 vccd1 _1717_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_24_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1583__B1 _1808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1858__S _1862_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1285_ _2015_/C _1285_/B vssd1 vssd1 vccd1 vccd1 _1947_/A sky130_fd_sc_hd__nand2_1
XANTENNA__1877__A1 _1239_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1354_ _1469_/A _1296_/B _1373_/A2 _1895_/B vssd1 vssd1 vccd1 vccd1 _1417_/B sky130_fd_sc_hd__a22o_1
X_1423_ _2205_/Q _1421_/A _1455_/B vssd1 vssd1 vccd1 vccd1 _1423_/X sky130_fd_sc_hd__a21o_2
XFILLER_0_46_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1087__A2 _1922_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1070_ _1825_/A _1128_/A _1075_/C vssd1 vssd1 vccd1 vccd1 _1467_/B sky130_fd_sc_hd__or3_4
XANTENNA_output36_A _2164_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1972_ _2015_/B _1995_/A _2001_/A _1972_/D vssd1 vssd1 vccd1 vccd1 _1972_/X sky130_fd_sc_hd__or4_1
XFILLER_0_28_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold19 hold19/A vssd1 vssd1 vccd1 vccd1 hold19/X sky130_fd_sc_hd__dlygate4sd3_1
X_1268_ _1871_/B hold7/X _2166_/Q vssd1 vssd1 vccd1 vccd1 _1945_/A sky130_fd_sc_hd__mux2_4
X_1337_ _1373_/A2 _1465_/B _1336_/X vssd1 vssd1 vccd1 vccd1 _1419_/A sky130_fd_sc_hd__a21bo_1
X_1406_ _1406_/A _1411_/C _1406_/C vssd1 vssd1 vccd1 vccd1 _1407_/D sky130_fd_sc_hd__or3_1
X_1199_ _1174_/B _1174_/C hold65/A vssd1 vssd1 vccd1 vccd1 _1199_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_52_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1527__A _1548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2171_ _2182_/CLK hold97/X vssd1 vssd1 vccd1 vccd1 _2171_/Q sky130_fd_sc_hd__dfxtp_1
X_1122_ _1462_/B _1723_/B vssd1 vssd1 vccd1 vccd1 _1123_/C sky130_fd_sc_hd__or2_1
XFILLER_0_20_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1053_ _1548_/A _1054_/C vssd1 vssd1 vccd1 vccd1 _1459_/A sky130_fd_sc_hd__nand2_1
X_1955_ _2043_/B _1955_/B _1955_/C _1955_/D vssd1 vssd1 vccd1 vccd1 _1955_/X sky130_fd_sc_hd__or4_1
XFILLER_0_43_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1886_ _1907_/S _1784_/A _1885_/X vssd1 vssd1 vccd1 vccd1 _1886_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_31_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1223__A2 _1864_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1257__A _1728_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1931__B1 _2003_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1695__C1 _1448_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1671_ _1697_/A _1595_/X _1668_/X _1670_/X vssd1 vssd1 vccd1 vccd1 _1674_/A sky130_fd_sc_hd__a22o_1
XANTENNA__1214__A2 _1868_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1740_ _2112_/Q _1765_/B vssd1 vssd1 vccd1 vccd1 _1742_/D sky130_fd_sc_hd__nand2_1
XFILLER_0_25_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2085_ _2225_/CLK hold76/X vssd1 vssd1 vccd1 vccd1 hold75/A sky130_fd_sc_hd__dfxtp_1
X_2154_ _2201_/CLK _2154_/D vssd1 vssd1 vccd1 vccd1 _2154_/Q sky130_fd_sc_hd__dfxtp_1
X_2223_ _2223_/CLK hold12/X vssd1 vssd1 vccd1 vccd1 hold11/A sky130_fd_sc_hd__dfxtp_1
X_1105_ _1441_/B _1486_/B _1907_/S vssd1 vssd1 vccd1 vccd1 _1829_/A sky130_fd_sc_hd__or3_1
XFILLER_0_48_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1036_ _1040_/B vssd1 vssd1 vccd1 vccd1 _1245_/A sky130_fd_sc_hd__inv_2
XFILLER_0_8_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1938_ hold53/X _1920_/Y _1937_/X vssd1 vssd1 vccd1 vccd1 hold54/A sky130_fd_sc_hd__a21o_1
X_1869_ _1871_/A _1869_/B vssd1 vssd1 vccd1 vccd1 _2157_/D sky130_fd_sc_hd__and2_1
XFILLER_0_31_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1654_ _1654_/A _1654_/B _1654_/C vssd1 vssd1 vccd1 vccd1 _1701_/A sky130_fd_sc_hd__and3_1
Xhold149 _2184_/Q vssd1 vssd1 vccd1 vccd1 _1033_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold116 _2134_/Q vssd1 vssd1 vccd1 vccd1 hold116/X sky130_fd_sc_hd__dlygate4sd3_1
X_1723_ _1723_/A _1723_/B _1723_/C vssd1 vssd1 vccd1 vccd1 _1724_/D sky130_fd_sc_hd__or3_1
Xhold105 _1793_/X vssd1 vssd1 vccd1 vccd1 _2129_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 _1756_/X vssd1 vssd1 vccd1 vccd1 _2123_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold127 _2125_/Q vssd1 vssd1 vccd1 vccd1 _1763_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2206_ _2206_/CLK _2206_/D vssd1 vssd1 vccd1 vccd1 _2206_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1585_ _2124_/Q _1826_/D _1460_/Y _1808_/A vssd1 vssd1 vccd1 vccd1 _1592_/S sky130_fd_sc_hd__a22o_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2068_ hold37/X _1503_/X _2075_/S vssd1 vssd1 vccd1 vccd1 hold38/A sky130_fd_sc_hd__mux2_1
X_2137_ _2150_/CLK _2137_/D vssd1 vssd1 vccd1 vccd1 _2137_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1270__A _1728_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1362__A1 _2160_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1370_ _1459_/B _1296_/B _1373_/A2 _1455_/B vssd1 vssd1 vccd1 vccd1 _1405_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_58_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1706_ _1921_/A hold194/X _1677_/X _1705_/Y vssd1 vssd1 vccd1 vccd1 _2113_/D sky130_fd_sc_hd__a22o_1
X_1637_ _1491_/B _1639_/A _1491_/A vssd1 vssd1 vccd1 vccd1 _1639_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_41_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1568_ _2107_/Q hold108/X _1994_/A vssd1 vssd1 vccd1 vccd1 _1568_/X sky130_fd_sc_hd__mux2_1
X_1499_ _1499_/A _1499_/B _1542_/A vssd1 vssd1 vccd1 vccd1 _1500_/B sky130_fd_sc_hd__and3_1
XFILLER_0_39_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout55 _1881_/A vssd1 vssd1 vccd1 vccd1 _1922_/B sky130_fd_sc_hd__buf_6
XFILLER_0_64_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout77 _1918_/A vssd1 vssd1 vccd1 vccd1 _2057_/A sky130_fd_sc_hd__buf_4
XFILLER_0_32_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout66 _1084_/A vssd1 vssd1 vccd1 vccd1 _1345_/A sky130_fd_sc_hd__buf_6
XFILLER_0_17_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1265__A _1728_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1886__A2 _1784_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1271__A0 _1156_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1422_ _2205_/Q _1141_/X _1421_/X vssd1 vssd1 vccd1 vccd1 _1422_/Y sky130_fd_sc_hd__a21boi_4
XANTENNA__1574__B2 _1156_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1284_ _1284_/A _1980_/B vssd1 vssd1 vccd1 vccd1 _1285_/B sky130_fd_sc_hd__nand2_2
XANTENNA__1629__A2 _1776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1353_ _1420_/B _1412_/A vssd1 vssd1 vccd1 vccd1 _1408_/A sky130_fd_sc_hd__or2_1
XANTENNA__1326__A1 _1717_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1801__A2 _1135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1971_ _1360_/B _1980_/B _1995_/B vssd1 vssd1 vccd1 vccd1 _1972_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_43_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1405_ _1405_/A _1405_/B _1405_/C _1414_/D vssd1 vssd1 vccd1 vccd1 _1406_/C sky130_fd_sc_hd__or4_1
XFILLER_0_11_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1198_ _1174_/B _1174_/C hold35/A vssd1 vssd1 vccd1 vccd1 _1198_/X sky130_fd_sc_hd__a21o_1
X_1267_ _1980_/B _2015_/C vssd1 vssd1 vccd1 vccd1 _1355_/B sky130_fd_sc_hd__or2_1
Xinput1 custom_settings[0] vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__buf_1
X_1336_ _1336_/A _1336_/B _1393_/A vssd1 vssd1 vccd1 vccd1 _1336_/X sky130_fd_sc_hd__or3_1
XFILLER_0_46_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1527__B _1868_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1808__A _1808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1718__A _1922_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2170_ _2172_/CLK hold2/X vssd1 vssd1 vccd1 vccd1 hold1/A sky130_fd_sc_hd__dfxtp_1
X_1052_ _1106_/A _1338_/A _1041_/Y vssd1 vssd1 vccd1 vccd1 _1054_/C sky130_fd_sc_hd__a21o_1
X_1121_ _1345_/A _1121_/B vssd1 vssd1 vccd1 vccd1 _1723_/B sky130_fd_sc_hd__nor2_1
X_1954_ _1996_/A _1954_/B vssd1 vssd1 vccd1 vccd1 _1955_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_7_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1885_ _1907_/S _2111_/Q _2206_/Q vssd1 vssd1 vccd1 vccd1 _1885_/X sky130_fd_sc_hd__and3b_1
XFILLER_0_43_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1768__A1 _2053_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1319_ _1061_/Y _1296_/B _2054_/A2 _1487_/A _1418_/A vssd1 vssd1 vccd1 vccd1 _1407_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1931__A1 _1920_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1720__B _1728_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1670_ _1622_/Y _1669_/Y _1654_/A vssd1 vssd1 vccd1 vccd1 _1670_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_7_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2222_ _2225_/CLK hold34/X vssd1 vssd1 vccd1 vccd1 hold33/A sky130_fd_sc_hd__dfxtp_1
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2153_ _2214_/CLK _2153_/D vssd1 vssd1 vccd1 vccd1 _2153_/Q sky130_fd_sc_hd__dfxtp_1
X_2084_ _2226_/CLK hold10/X vssd1 vssd1 vccd1 vccd1 hold9/A sky130_fd_sc_hd__dfxtp_1
X_1104_ _1104_/A _1131_/C vssd1 vssd1 vccd1 vccd1 _1907_/S sky130_fd_sc_hd__and2_4
X_1035_ _2144_/Q vssd1 vssd1 vccd1 vccd1 _1035_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_17_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1937_ _1920_/A _2097_/Q _1920_/B _1243_/B vssd1 vssd1 vccd1 vccd1 _1937_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_8_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1868_ _2049_/A _1868_/B vssd1 vssd1 vccd1 vccd1 _2156_/D sky130_fd_sc_hd__and2_1
X_1799_ _2053_/B2 _1797_/Y _1804_/A _1820_/A2 _1794_/A vssd1 vssd1 vccd1 vccd1 _1799_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_58_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1653_ _1653_/A _1653_/B vssd1 vssd1 vccd1 vccd1 _1653_/Y sky130_fd_sc_hd__nor2_1
X_1584_ _2115_/Q _1460_/A _1468_/A _1162_/X _1583_/X vssd1 vssd1 vccd1 vccd1 _1584_/X
+ sky130_fd_sc_hd__a221o_1
Xhold117 _1820_/X vssd1 vssd1 vccd1 vccd1 _2134_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold106 _2131_/Q vssd1 vssd1 vccd1 vccd1 _1800_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1722_ _1104_/A _1245_/C _1826_/D _1062_/Y _1903_/B vssd1 vssd1 vccd1 vccd1 _1723_/C
+ sky130_fd_sc_hd__a2111o_1
Xhold139 _2119_/Q vssd1 vssd1 vccd1 vccd1 hold139/X sky130_fd_sc_hd__buf_1
Xhold128 _1768_/X vssd1 vssd1 vccd1 vccd1 _2125_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2205_ _2206_/CLK _2205_/D vssd1 vssd1 vccd1 vccd1 _2205_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2067_ _1499_/A _1882_/B _1498_/B _2003_/A vssd1 vssd1 vccd1 vccd1 _2075_/S sky130_fd_sc_hd__a31o_4
XFILLER_0_48_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2136_ _2150_/CLK _2136_/D vssd1 vssd1 vccd1 vccd1 _2136_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1362__A2 _2165_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout78_A _1920_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1705_ _1921_/A _1705_/B vssd1 vssd1 vccd1 vccd1 _1705_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_45_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1567_ hold5/X _1549_/X _1567_/S vssd1 vssd1 vccd1 vccd1 hold6/A sky130_fd_sc_hd__mux2_1
X_1636_ _1611_/Y _1635_/X _1654_/A vssd1 vssd1 vccd1 vccd1 _1639_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_41_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1498_ _1918_/A _1498_/B vssd1 vssd1 vccd1 vccd1 _1542_/A sky130_fd_sc_hd__and2_2
XANTENNA__1090__B _1922_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2119_ _2164_/CLK _2119_/D vssd1 vssd1 vccd1 vccd1 _2119_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout78 _1920_/A vssd1 vssd1 vccd1 vccd1 _1994_/A sky130_fd_sc_hd__buf_6
Xfanout56 _1403_/A2 vssd1 vssd1 vccd1 vccd1 _1340_/B sky130_fd_sc_hd__buf_4
Xfanout67 _1041_/Y vssd1 vssd1 vccd1 vccd1 _1377_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_44_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1583__A2 _1776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1574__A2 _1826_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1421_ _1421_/A _1895_/B vssd1 vssd1 vccd1 vccd1 _1421_/X sky130_fd_sc_hd__or2_1
X_1283_ _1728_/B _1980_/B vssd1 vssd1 vccd1 vccd1 _1960_/B sky130_fd_sc_hd__and2_2
X_1352_ _1517_/A _1373_/A2 _1303_/Y _1313_/Y vssd1 vssd1 vccd1 vccd1 _1412_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_61_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1619_ _1882_/A _1175_/X _1176_/X _1468_/A vssd1 vssd1 vccd1 vccd1 _1622_/A sky130_fd_sc_hd__o211ai_4
XFILLER_0_1_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1789__C1 _1717_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1970_ _2028_/B _1964_/A _1968_/X _1969_/X vssd1 vssd1 vccd1 vccd1 _2179_/D sky130_fd_sc_hd__a31o_1
XFILLER_0_70_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1795__A2 _1135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1335_ _1377_/A _1335_/B vssd1 vssd1 vccd1 vccd1 _1465_/B sky130_fd_sc_hd__nor2_1
X_1404_ _1404_/A _1404_/B vssd1 vssd1 vccd1 vccd1 _1411_/C sky130_fd_sc_hd__or2_1
Xinput2 custom_settings[1] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__buf_1
X_1266_ _1728_/B _1266_/B vssd1 vssd1 vccd1 vccd1 _2015_/C sky130_fd_sc_hd__nand2_4
X_1197_ _1732_/A _1149_/Y _1196_/X vssd1 vssd1 vccd1 vccd1 _1197_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_46_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_6_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _2208_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_32_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1777__A2 _1135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1718__B _1728_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1934__C1 _1871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1120_ _1344_/A _1335_/B vssd1 vssd1 vccd1 vccd1 _1462_/B sky130_fd_sc_hd__nor2_1
X_1051_ _1377_/A _1106_/A vssd1 vssd1 vccd1 vccd1 _1051_/Y sky130_fd_sc_hd__nor2_1
X_1953_ _1995_/A _2001_/A vssd1 vssd1 vccd1 vccd1 _1954_/B sky130_fd_sc_hd__nor2_1
X_1884_ _1895_/B _1881_/X _1883_/X _2197_/Q vssd1 vssd1 vccd1 vccd1 _1884_/Y sky130_fd_sc_hd__o22ai_2
XFILLER_0_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1217__A1 hold194/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_3_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1909__A _2057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1318_ _1229_/D _1373_/A2 _1285_/B _1317_/Y vssd1 vssd1 vccd1 vccd1 _1418_/A sky130_fd_sc_hd__a22o_1
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1249_ _1728_/B _1249_/B vssd1 vssd1 vccd1 vccd1 _1297_/A sky130_fd_sc_hd__and2_2
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1448__B _1448_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2152_ _2172_/CLK _2152_/D vssd1 vssd1 vccd1 vccd1 _2152_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2221_ _2225_/CLK hold40/X vssd1 vssd1 vccd1 vccd1 hold39/A sky130_fd_sc_hd__dfxtp_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2083_ _2225_/CLK hold66/X vssd1 vssd1 vccd1 vccd1 hold65/A sky130_fd_sc_hd__dfxtp_1
X_1034_ hold93/X vssd1 vssd1 vccd1 vccd1 _1034_/Y sky130_fd_sc_hd__inv_2
X_1103_ _1821_/A _1236_/D _1114_/B _1821_/B vssd1 vssd1 vccd1 vccd1 _1131_/C sky130_fd_sc_hd__and4b_1
X_1867_ _2049_/A _1867_/B vssd1 vssd1 vccd1 vccd1 _2155_/D sky130_fd_sc_hd__and2_1
X_1936_ hold27/X _1920_/Y _1935_/X vssd1 vssd1 vccd1 vccd1 hold28/A sky130_fd_sc_hd__a21o_1
XANTENNA__1610__A1 _2112_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1798_ _1797_/B _1797_/C _1797_/D _1797_/A vssd1 vssd1 vccd1 vccd1 _1804_/A sky130_fd_sc_hd__a31o_1
XFILLER_0_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1284__A _1284_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1721_ _2110_/Q _1765_/B _1776_/B _2143_/Q vssd1 vssd1 vccd1 vccd1 _1726_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_5_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1652_ _1651_/Y _1650_/B _1652_/S vssd1 vssd1 vccd1 vccd1 _1653_/B sky130_fd_sc_hd__mux2_1
X_1583_ _2140_/Q _1776_/A _1808_/A _1469_/X vssd1 vssd1 vccd1 vccd1 _1583_/X sky130_fd_sc_hd__a22o_1
Xhold118 _2133_/Q vssd1 vssd1 vccd1 vccd1 hold118/X sky130_fd_sc_hd__buf_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold107 _1805_/X vssd1 vssd1 vccd1 vccd1 _2131_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold129 _2122_/Q vssd1 vssd1 vccd1 vccd1 _1745_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1922__A _1994_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2204_ _1233_/A _2204_/D vssd1 vssd1 vccd1 vccd1 _2204_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2135_ _2150_/CLK _2135_/D vssd1 vssd1 vccd1 vccd1 _2135_/Q sky130_fd_sc_hd__dfxtp_1
X_2066_ hold45/X _1549_/X _2066_/S vssd1 vssd1 vccd1 vccd1 hold46/A sky130_fd_sc_hd__mux2_1
XFILLER_0_48_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1919_ _1920_/A _1920_/B vssd1 vssd1 vccd1 vccd1 _1933_/B sky130_fd_sc_hd__and2_1
XFILLER_0_44_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1362__A3 _2161_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1510__B1 _1548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1813__A1 _1156_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1704_ hold200/X _1662_/X _1920_/A vssd1 vssd1 vccd1 vccd1 _2112_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_41_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1566_ hold19/X _1542_/X _1567_/S vssd1 vssd1 vccd1 vccd1 hold20/A sky130_fd_sc_hd__mux2_1
X_1497_ _1517_/A _1825_/B _1110_/D _1496_/X _1994_/A vssd1 vssd1 vccd1 vccd1 _1498_/B
+ sky130_fd_sc_hd__o41a_2
X_1635_ _1633_/Y _1634_/X _1635_/S vssd1 vssd1 vccd1 vccd1 _1635_/X sky130_fd_sc_hd__mux2_1
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2118_ _2223_/CLK hold92/X vssd1 vssd1 vccd1 vccd1 hold91/A sky130_fd_sc_hd__dfxtp_1
X_2049_ _2049_/A _2049_/B vssd1 vssd1 vccd1 vccd1 _2205_/D sky130_fd_sc_hd__and2_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout79 input13/X vssd1 vssd1 vccd1 vccd1 _1920_/A sky130_fd_sc_hd__buf_6
Xfanout57 _2054_/A2 vssd1 vssd1 vccd1 vccd1 _1403_/A2 sky130_fd_sc_hd__clkbuf_4
Xfanout68 _2080_/Q vssd1 vssd1 vccd1 vccd1 _1821_/A sky130_fd_sc_hd__buf_4
XFILLER_0_32_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1559__B1 _2003_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_8_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1351_ _1051_/Y _1373_/A2 _1276_/Y _1313_/Y vssd1 vssd1 vccd1 vccd1 _1420_/B sky130_fd_sc_hd__a22o_1
X_1420_ _1420_/A _1420_/B _1420_/C _1420_/D vssd1 vssd1 vccd1 vccd1 _2082_/D sky130_fd_sc_hd__or4_1
X_1282_ _1306_/B _1980_/B _1355_/C _1281_/Y vssd1 vssd1 vccd1 vccd1 _1282_/X sky130_fd_sc_hd__o31a_1
XFILLER_0_73_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1618_ _1611_/Y _1617_/Y _1654_/A vssd1 vssd1 vccd1 vccd1 _1618_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_41_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1549_ _1548_/A _1871_/B _1542_/A _1548_/Y vssd1 vssd1 vccd1 vccd1 _1549_/X sky130_fd_sc_hd__o211a_1
XANTENNA__1722__B1 _1826_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1265_ _1728_/B _1266_/B vssd1 vssd1 vccd1 vccd1 _1995_/A sky130_fd_sc_hd__and2_4
X_1334_ _1391_/A _1417_/A _1405_/A _1334_/D vssd1 vssd1 vccd1 vccd1 _1375_/A sky130_fd_sc_hd__or4_1
X_1403_ _1723_/B _1403_/A2 _1346_/B _1415_/A3 _1333_/C vssd1 vssd1 vccd1 vccd1 _1404_/B
+ sky130_fd_sc_hd__a221o_1
Xinput3 io_in[19] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__1483__A2 _2160_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1196_ hold177/X _1149_/B _1193_/X _1467_/A _1195_/X vssd1 vssd1 vccd1 vccd1 _1196_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__1824__B _1922_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1171__B2 _1868_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1050_ _1377_/A _1338_/A vssd1 vssd1 vccd1 vccd1 _1824_/A sky130_fd_sc_hd__nor2_1
X_1952_ _1980_/A _1285_/B _1984_/C _1306_/A _1995_/A vssd1 vssd1 vccd1 vccd1 _1955_/C
+ sky130_fd_sc_hd__o2111a_1
X_1883_ hold120/X _1882_/Y _1921_/B _1912_/A _2006_/A vssd1 vssd1 vccd1 vccd1 _1883_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1248_ _1796_/A hold1/X _1923_/A vssd1 vssd1 vccd1 vccd1 _1249_/B sky130_fd_sc_hd__mux2_1
X_1317_ _1393_/A _1317_/B vssd1 vssd1 vccd1 vccd1 _1317_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_2_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1208__A2 _1871_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1179_ hold186/X _1149_/C _1827_/B _1796_/A vssd1 vssd1 vccd1 vccd1 _1179_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_2_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1916__A0 _1870_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1835__A _1863_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1931__A3 _1920_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_362 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2220_ _2226_/CLK hold58/X vssd1 vssd1 vccd1 vccd1 hold57/A sky130_fd_sc_hd__dfxtp_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2151_ _2208_/CLK _2151_/D vssd1 vssd1 vccd1 vccd1 _2151_/Q sky130_fd_sc_hd__dfxtp_1
X_1102_ _1377_/A _1102_/B vssd1 vssd1 vccd1 vccd1 _1486_/B sky130_fd_sc_hd__nor2_1
X_2082_ _2210_/CLK _2082_/D vssd1 vssd1 vccd1 vccd1 _2082_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_56_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1033_ _1033_/A vssd1 vssd1 vccd1 vccd1 _1033_/Y sky130_fd_sc_hd__inv_2
X_1935_ _1920_/A _2096_/Q _1920_/B _2003_/A vssd1 vssd1 vccd1 vccd1 _1935_/X sky130_fd_sc_hd__a31o_1
X_1866_ _2049_/A _1866_/B vssd1 vssd1 vccd1 vccd1 _2154_/D sky130_fd_sc_hd__and2_1
X_1797_ _1797_/A _1797_/B _1797_/C _1797_/D vssd1 vssd1 vccd1 vccd1 _1797_/Y sky130_fd_sc_hd__nand4_1
XFILLER_0_12_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold108 _2098_/Q vssd1 vssd1 vccd1 vccd1 hold108/X sky130_fd_sc_hd__dlygate4sd3_1
X_1651_ _1651_/A _1654_/C vssd1 vssd1 vccd1 vccd1 _1651_/Y sky130_fd_sc_hd__nand2_1
X_1720_ _1921_/B _1728_/B vssd1 vssd1 vccd1 vccd1 _1776_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_5_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1582_ _1582_/A _1582_/B _1582_/C vssd1 vssd1 vccd1 vccd1 _1689_/B sky130_fd_sc_hd__and3_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold119 _1816_/X vssd1 vssd1 vccd1 vccd1 _2133_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2065_ hold29/X _1542_/X _2066_/S vssd1 vssd1 vccd1 vccd1 hold30/A sky130_fd_sc_hd__mux2_1
XANTENNA__1922__B _1922_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2203_ _1233_/A _2203_/D vssd1 vssd1 vccd1 vccd1 _2203_/Q sky130_fd_sc_hd__dfxtp_1
X_2134_ _2142_/CLK _2134_/D vssd1 vssd1 vccd1 vccd1 _2134_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1918_ _1918_/A _1918_/B vssd1 vssd1 vccd1 vccd1 _2165_/D sky130_fd_sc_hd__and2_1
XFILLER_0_44_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1849_ _1863_/A _1849_/B vssd1 vssd1 vccd1 vccd1 _2143_/D sky130_fd_sc_hd__and2_1
XFILLER_0_8_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1807__C1 _1717_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1703_ hold177/X _1663_/Y _1920_/A vssd1 vssd1 vccd1 vccd1 _2111_/D sky130_fd_sc_hd__mux2_1
X_1634_ _1669_/A _1474_/B _1638_/S _1632_/X vssd1 vssd1 vccd1 vccd1 _1634_/X sky130_fd_sc_hd__o31a_1
XFILLER_0_26_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1565_ hold31/X _1535_/X _1567_/S vssd1 vssd1 vccd1 vccd1 hold32/A sky130_fd_sc_hd__mux2_1
X_1496_ _2206_/Q _2177_/Q _1922_/B vssd1 vssd1 vccd1 vccd1 _1496_/X sky130_fd_sc_hd__and3b_1
XFILLER_0_39_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2117_ _2223_/CLK _2117_/D vssd1 vssd1 vccd1 vccd1 _2117_/Q sky130_fd_sc_hd__dfxtp_2
X_2048_ _2015_/C _1955_/B _2043_/Y _2043_/B hold196/X vssd1 vssd1 vccd1 vccd1 _2048_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_44_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout58 _2054_/A2 vssd1 vssd1 vccd1 vccd1 _1373_/A2 sky130_fd_sc_hd__buf_4
XFILLER_0_32_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout69 _2079_/Q vssd1 vssd1 vccd1 vccd1 _1236_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_0_32_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1843__A _1863_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1256__A0 _1864_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1281_ _1946_/A _1281_/B vssd1 vssd1 vccd1 vccd1 _1281_/Y sky130_fd_sc_hd__nor2_1
X_1350_ _1392_/A _1375_/A _1419_/A _1350_/D vssd1 vssd1 vccd1 vccd1 _1402_/A sky130_fd_sc_hd__or4_1
XFILLER_0_58_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1247__B1 _1025_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1617_ _1669_/A _1617_/B vssd1 vssd1 vccd1 vccd1 _1617_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_41_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1548_ _1548_/A _1548_/B vssd1 vssd1 vccd1 vccd1 _1548_/Y sky130_fd_sc_hd__nand2_1
X_1479_ _1475_/Y _1476_/X _1477_/Y _1478_/X _1654_/A vssd1 vssd1 vccd1 vccd1 _1479_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_37_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1789__A1 _2112_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1402_ _1402_/A _1402_/B _1402_/C _1402_/D vssd1 vssd1 vccd1 vccd1 _1402_/X sky130_fd_sc_hd__or4_1
XFILLER_0_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput4 io_in[20] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__clkbuf_1
X_1264_ _1808_/A hold27/X _2166_/Q vssd1 vssd1 vccd1 vccd1 _1266_/B sky130_fd_sc_hd__mux2_1
X_1333_ _1389_/A _1333_/B _1333_/C _1390_/A vssd1 vssd1 vccd1 vccd1 _1334_/D sky130_fd_sc_hd__or4_1
X_1195_ _2144_/Q _1149_/C _1827_/B _1784_/A vssd1 vssd1 vccd1 vccd1 _1195_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1815__B1_N _2053_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output27_A _2161_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1882_ _1882_/A _1882_/B vssd1 vssd1 vccd1 vccd1 _1882_/Y sky130_fd_sc_hd__nand2_1
X_1951_ _1955_/B vssd1 vssd1 vccd1 vccd1 _1951_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_3_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1178_ hold228/X _2094_/Q _1994_/A vssd1 vssd1 vccd1 vccd1 _1796_/A sky130_fd_sc_hd__mux2_4
XFILLER_0_47_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1247_ _2163_/Q _1039_/Y _1025_/Y vssd1 vssd1 vccd1 vccd1 _1284_/A sky130_fd_sc_hd__o21a_1
XANTENNA__1941__A _2057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1316_ _1409_/A _1420_/A _1410_/A vssd1 vssd1 vccd1 vccd1 _1392_/A sky130_fd_sc_hd__or3_1
XFILLER_0_2_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1851__A _1863_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1032_ _2185_/Q vssd1 vssd1 vccd1 vccd1 _1032_/Y sky130_fd_sc_hd__inv_2
X_1101_ _1345_/A _1102_/B _1121_/B _1344_/A vssd1 vssd1 vccd1 vccd1 _1441_/B sky130_fd_sc_hd__o22ai_4
X_2081_ _2210_/CLK _2081_/D vssd1 vssd1 vccd1 vccd1 _2081_/Q sky130_fd_sc_hd__dfxtp_2
X_2150_ _2150_/CLK _2150_/D vssd1 vssd1 vccd1 vccd1 _2150_/Q sky130_fd_sc_hd__dfxtp_1
X_1934_ hold96/X _1920_/Y _1933_/X _1871_/A vssd1 vssd1 vccd1 vccd1 hold97/A sky130_fd_sc_hd__o211a_1
XFILLER_0_56_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1700__S _1920_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1865_ _2000_/A _1865_/B vssd1 vssd1 vccd1 vccd1 _2153_/D sky130_fd_sc_hd__and2_1
X_1796_ _1796_/A _1808_/B vssd1 vssd1 vccd1 vccd1 _1797_/D sky130_fd_sc_hd__nand2_1
XFILLER_0_12_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold109 _1568_/X vssd1 vssd1 vccd1 vccd1 _2107_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1650_ _1650_/A _1650_/B vssd1 vssd1 vccd1 vccd1 _1654_/C sky130_fd_sc_hd__nand2_1
X_1581_ _1651_/A _1491_/B _1581_/S vssd1 vssd1 vccd1 vccd1 _1582_/C sky130_fd_sc_hd__mux2_1
X_2202_ _1233_/A _2202_/D vssd1 vssd1 vccd1 vccd1 _2202_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2064_ hold23/X _1535_/X _2066_/S vssd1 vssd1 vccd1 vccd1 hold24/A sky130_fd_sc_hd__mux2_1
XFILLER_0_48_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2133_ _2142_/CLK _2133_/D vssd1 vssd1 vccd1 vccd1 _2133_/Q sky130_fd_sc_hd__dfxtp_1
X_1917_ _1916_/X hold232/X _1917_/S vssd1 vssd1 vccd1 vccd1 _1917_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_29_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1779_ _1780_/B _1780_/C _1780_/D _1780_/A vssd1 vssd1 vccd1 vccd1 _1785_/A sky130_fd_sc_hd__a31o_1
X_1848_ hold176/X _1206_/X _1862_/S vssd1 vssd1 vccd1 vccd1 _1849_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_8_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold160_A _2117_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_300 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1564_ hold15/X _1528_/X _1567_/S vssd1 vssd1 vccd1 vccd1 hold16/A sky130_fd_sc_hd__mux2_1
XFILLER_0_53_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1702_ hold175/X _1701_/Y _1920_/A vssd1 vssd1 vccd1 vccd1 _2110_/D sky130_fd_sc_hd__mux2_1
X_1633_ _1669_/A _1638_/S vssd1 vssd1 vccd1 vccd1 _1633_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_30_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1495_ hold85/X _1494_/Y _1920_/A vssd1 vssd1 vccd1 vccd1 hold86/A sky130_fd_sc_hd__mux2_1
XFILLER_0_39_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2116_ _2223_/CLK _2116_/D vssd1 vssd1 vccd1 vccd1 _2116_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_49_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2047_ _2057_/A _2047_/B vssd1 vssd1 vccd1 vccd1 _2204_/D sky130_fd_sc_hd__and2_1
XFILLER_0_72_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout48 _1923_/B vssd1 vssd1 vccd1 vccd1 _2043_/B sky130_fd_sc_hd__buf_4
Xfanout59 _1243_/Y vssd1 vssd1 vccd1 vccd1 _2054_/A2 sky130_fd_sc_hd__buf_2
XFILLER_0_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout76_A _2057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1280_ _2036_/A _1355_/B _1355_/C _1279_/A _1287_/B vssd1 vssd1 vccd1 vccd1 _1300_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_0_31_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1731__A2 _1717_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1247__A1 _2163_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1547_ _1547_/A _1547_/B vssd1 vssd1 vccd1 vccd1 _1548_/B sky130_fd_sc_hd__xnor2_1
X_1616_ _1632_/A _1614_/X _1615_/Y _1475_/Y vssd1 vssd1 vccd1 vccd1 _1616_/X sky130_fd_sc_hd__a211o_1
X_1478_ _1492_/A _1632_/A _1476_/B vssd1 vssd1 vccd1 vccd1 _1478_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_49_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1789__A2 _1135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_4_12_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1467__C _1920_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1401_ _1401_/A _1401_/B _1408_/C _1401_/D vssd1 vssd1 vccd1 vccd1 _1402_/D sky130_fd_sc_hd__or4_1
XFILLER_0_11_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput5 io_in[21] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__clkbuf_1
X_1194_ hold224/X _2092_/Q _1994_/A vssd1 vssd1 vccd1 vccd1 _1784_/A sky130_fd_sc_hd__mux2_4
X_1263_ _1868_/B hold241/X _1923_/A vssd1 vssd1 vccd1 vccd1 _1980_/B sky130_fd_sc_hd__mux2_2
XANTENNA__1703__S _1920_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1332_ _1776_/A _1365_/A _1331_/X _1340_/B _1135_/A vssd1 vssd1 vccd1 vccd1 _1390_/A
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1631__B2 _1784_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1849__A _1863_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1950_ _2036_/A _1960_/B vssd1 vssd1 vccd1 vccd1 _1955_/B sky130_fd_sc_hd__nor2_2
X_1881_ _1881_/A _1907_/S vssd1 vssd1 vccd1 vccd1 _1881_/X sky130_fd_sc_hd__or2_2
XFILLER_0_22_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1941__B _1941_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1315_ _1116_/C _1296_/B _1241_/A _1373_/A2 _1238_/B vssd1 vssd1 vccd1 vccd1 _1410_/A
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_11_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1177_ _1882_/A _1175_/X _1176_/X vssd1 vssd1 vccd1 vccd1 _1177_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_47_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1246_ _1296_/B _1242_/X _1373_/A2 _1448_/B vssd1 vssd1 vccd1 vccd1 _1312_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_2_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1031_ _1997_/A vssd1 vssd1 vccd1 vccd1 _1031_/Y sky130_fd_sc_hd__inv_2
X_2080_ _2210_/CLK _2080_/D vssd1 vssd1 vccd1 vccd1 _2080_/Q sky130_fd_sc_hd__dfxtp_2
X_1100_ _1345_/A _1102_/B vssd1 vssd1 vccd1 vccd1 _1100_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1933_ _2171_/Q _1933_/B vssd1 vssd1 vccd1 vccd1 _1933_/X sky130_fd_sc_hd__or2_1
X_1864_ _2000_/A _1864_/B vssd1 vssd1 vccd1 vccd1 _2152_/D sky130_fd_sc_hd__and2_1
Xclkbuf_4_5_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _2226_/CLK sky130_fd_sc_hd__clkbuf_8
X_1795_ _2113_/Q _1135_/A _1776_/X _2138_/Q _1717_/B vssd1 vssd1 vccd1 vccd1 _1797_/C
+ sky130_fd_sc_hd__a221oi_2
XFILLER_0_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1163__S _1994_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1229_ _1462_/B _1229_/B _1229_/C _1229_/D vssd1 vssd1 vccd1 vccd1 _1229_/X sky130_fd_sc_hd__or4_2
XFILLER_0_62_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1580_ _1491_/B _1582_/A _1491_/A vssd1 vssd1 vccd1 vccd1 _1582_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_0_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2201_ _2201_/CLK _2201_/D vssd1 vssd1 vccd1 vccd1 _2201_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2132_ _2142_/CLK _2132_/D vssd1 vssd1 vccd1 vccd1 _2132_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2063_ hold63/X _1528_/X _2066_/S vssd1 vssd1 vccd1 vccd1 hold64/A sky130_fd_sc_hd__mux2_1
XANTENNA__1711__S _1920_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1916_ _1870_/B _1914_/X _1922_/B vssd1 vssd1 vccd1 vccd1 _1916_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_44_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1847_ _1863_/A _1847_/B vssd1 vssd1 vccd1 vccd1 _2142_/D sky130_fd_sc_hd__and2_1
X_1778_ _1864_/B _1808_/B vssd1 vssd1 vccd1 vccd1 _1780_/D sky130_fd_sc_hd__nand2_1
XFILLER_0_8_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1752__B1 _1717_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1857__A _1863_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1701_ _1701_/A _1701_/B vssd1 vssd1 vccd1 vccd1 _1701_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_26_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1563_ hold69/X _1525_/X _1567_/S vssd1 vssd1 vccd1 vccd1 hold70/A sky130_fd_sc_hd__mux2_1
X_1494_ _1570_/B vssd1 vssd1 vccd1 vccd1 _1494_/Y sky130_fd_sc_hd__inv_2
X_1632_ _1632_/A _1632_/B _1638_/S vssd1 vssd1 vccd1 vccd1 _1632_/X sky130_fd_sc_hd__or3b_1
XFILLER_0_39_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2115_ _2223_/CLK _2115_/D vssd1 vssd1 vccd1 vccd1 _2115_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout49 _1922_/Y vssd1 vssd1 vccd1 vccd1 _1923_/B sky130_fd_sc_hd__clkbuf_4
X_2046_ _1873_/B _2043_/B _2036_/Y _2043_/Y vssd1 vssd1 vccd1 vccd1 _2047_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1546_ _1913_/A _2117_/Q _1546_/S vssd1 vssd1 vccd1 vccd1 _1547_/B sky130_fd_sc_hd__mux2_1
X_1477_ _1492_/A _1476_/B _1669_/A vssd1 vssd1 vccd1 vccd1 _1477_/Y sky130_fd_sc_hd__a21oi_1
X_1615_ _1611_/A _1611_/B _1617_/B _1632_/B vssd1 vssd1 vccd1 vccd1 _1615_/Y sky130_fd_sc_hd__a211oi_1
X_2029_ _1923_/B _2015_/Y _2028_/X _2000_/A vssd1 vssd1 vccd1 vccd1 _2029_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_37_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1870__A _1871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1331_ _2107_/Q _2108_/Q vssd1 vssd1 vccd1 vccd1 _1331_/X sky130_fd_sc_hd__xor2_2
X_1400_ _1403_/A2 _1724_/A _1413_/C _1417_/D vssd1 vssd1 vccd1 vccd1 _1401_/D sky130_fd_sc_hd__a211o_1
XFILLER_0_11_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput6 io_in[22] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__clkbuf_1
X_1193_ _1191_/X _1192_/X _1499_/A vssd1 vssd1 vccd1 vccd1 _1193_/X sky130_fd_sc_hd__mux2_1
X_1262_ _1946_/A _2015_/B vssd1 vssd1 vccd1 vccd1 _2036_/A sky130_fd_sc_hd__or2_2
XFILLER_0_52_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1529_ hold51/X _1528_/X _1550_/S vssd1 vssd1 vccd1 vccd1 hold52/A sky130_fd_sc_hd__mux2_1
XFILLER_0_45_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1631__A2 _1826_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1147__B2 _1871_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1880_ _2057_/A _1880_/B vssd1 vssd1 vccd1 vccd1 _2160_/D sky130_fd_sc_hd__and2_1
XFILLER_0_28_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1314_ _1824_/A _1373_/A2 _1286_/Y _1313_/Y vssd1 vssd1 vccd1 vccd1 _1420_/A sky130_fd_sc_hd__a22o_1
X_1176_ hold71/A _1499_/B _1174_/X _1499_/A vssd1 vssd1 vccd1 vccd1 _1176_/X sky130_fd_sc_hd__a211o_1
X_1245_ _1245_/A _1245_/B _1245_/C vssd1 vssd1 vccd1 vccd1 _1448_/B sky130_fd_sc_hd__and3_4
XFILLER_0_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2023__C1 _2003_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2014__C1 _2003_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1030_ _2192_/Q vssd1 vssd1 vccd1 vccd1 _1030_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_68_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1932_ hold1/X _1920_/Y _1931_/X vssd1 vssd1 vccd1 vccd1 hold2/A sky130_fd_sc_hd__a21o_1
XFILLER_0_56_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1863_ _1863_/A _1863_/B vssd1 vssd1 vccd1 vccd1 _2150_/D sky130_fd_sc_hd__and2_1
XFILLER_0_58_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1794_ _1794_/A _1806_/B vssd1 vssd1 vccd1 vccd1 _1797_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1531__A1 _2108_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1228_ _1895_/B _1228_/B vssd1 vssd1 vccd1 vccd1 _1228_/Y sky130_fd_sc_hd__nor2_2
X_1159_ _1763_/A _1149_/Y _1158_/X vssd1 vssd1 vccd1 vccd1 _1159_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_15_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2062_ hold71/X _1525_/X _2066_/S vssd1 vssd1 vccd1 vccd1 hold72/A sky130_fd_sc_hd__mux2_1
X_2200_ _2206_/CLK _2200_/D vssd1 vssd1 vccd1 vccd1 _2200_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2131_ _2142_/CLK _2131_/D vssd1 vssd1 vccd1 vccd1 _2131_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_310 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1915_ _1031_/Y _1922_/B _1912_/Y _1893_/Y vssd1 vssd1 vccd1 vccd1 _1917_/S sky130_fd_sc_hd__a31o_1
XFILLER_0_44_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1846_ hold204/X _1209_/X _1862_/S vssd1 vssd1 vccd1 vccd1 _1846_/X sky130_fd_sc_hd__mux2_1
X_1777_ _2110_/Q _1135_/A _1776_/X _2135_/Q _1717_/B vssd1 vssd1 vccd1 vccd1 _1780_/C
+ sky130_fd_sc_hd__a221oi_2
XFILLER_0_4_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1268__A0 _1871_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1807__A2 _1135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1873__A _1912_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1743__A1 _2053_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1259__A0 _1784_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1700_ hold89/X _1707_/B _1920_/A vssd1 vssd1 vccd1 vccd1 hold90/A sky130_fd_sc_hd__mux2_1
X_1631_ _2120_/Q _1826_/D _1460_/Y _1784_/A vssd1 vssd1 vccd1 vccd1 _1638_/S sky130_fd_sc_hd__a22oi_4
XFILLER_0_38_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1562_ hold59/X _1519_/X _1567_/S vssd1 vssd1 vccd1 vccd1 hold60/A sky130_fd_sc_hd__mux2_1
X_1493_ _1650_/B _1492_/A _1490_/X _1492_/Y vssd1 vssd1 vccd1 vccd1 _1570_/B sky130_fd_sc_hd__a211o_1
XTAP_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2114_ _2223_/CLK _2114_/D vssd1 vssd1 vccd1 vccd1 _2114_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_49_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2045_ _2057_/A _2045_/B vssd1 vssd1 vccd1 vccd1 _2203_/D sky130_fd_sc_hd__and2_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1829_ _1829_/A _1829_/B _1829_/C _1829_/D vssd1 vssd1 vccd1 vccd1 _1831_/B sky130_fd_sc_hd__or4_1
XFILLER_0_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1778__A _1864_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1614_ _1611_/A _1611_/B _1617_/B vssd1 vssd1 vccd1 vccd1 _1614_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1545_ _2108_/Q _1545_/B vssd1 vssd1 vccd1 vccd1 _1913_/A sky130_fd_sc_hd__xnor2_1
X_1476_ _1492_/A _1476_/B _1476_/C vssd1 vssd1 vccd1 vccd1 _1476_/X sky130_fd_sc_hd__and3_1
XFILLER_0_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2028_ _2028_/A _2028_/B vssd1 vssd1 vccd1 vccd1 _2028_/X sky130_fd_sc_hd__or2_1
XANTENNA__1891__B1 _1918_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1870__B _1870_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1937__A1 _1920_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1261_ _1281_/B _1306_/B vssd1 vssd1 vccd1 vccd1 _2015_/B sky130_fd_sc_hd__or2_2
X_1330_ _1517_/A _1415_/A3 _1340_/B _1100_/Y vssd1 vssd1 vccd1 vccd1 _1333_/C sky130_fd_sc_hd__a22o_1
Xinput7 io_in[23] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__clkbuf_1
X_1192_ hold9/A hold57/A _1882_/B vssd1 vssd1 vccd1 vccd1 _1192_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_46_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1528_ _2114_/Q _1517_/A _1542_/A _1527_/X vssd1 vssd1 vccd1 vccd1 _1528_/X sky130_fd_sc_hd__o211a_1
X_1459_ _1459_/A _1459_/B _1459_/C _1465_/B vssd1 vssd1 vccd1 vccd1 _1460_/D sky130_fd_sc_hd__or4_1
XANTENNA__1865__B _1865_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1313_ _1393_/A _1313_/B vssd1 vssd1 vccd1 vccd1 _1313_/Y sky130_fd_sc_hd__nor2_1
X_1244_ _1104_/A _1245_/C _1340_/B _1826_/B _1415_/A3 vssd1 vssd1 vccd1 vccd1 _1414_/A
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_2_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1175_ hold33/A hold43/A _1499_/B vssd1 vssd1 vccd1 vccd1 _1175_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_63_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xmax_cap47 _1149_/Y vssd1 vssd1 vccd1 vccd1 _1150_/S sky130_fd_sc_hd__buf_4
XFILLER_0_21_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput10 io_in[26] vssd1 vssd1 vccd1 vccd1 _1558_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1931_ _1920_/A _2094_/Q _1920_/B _2003_/A vssd1 vssd1 vccd1 vccd1 _1931_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_56_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1793_ _2053_/B2 _1797_/A _1792_/Y _1820_/A2 _1788_/A vssd1 vssd1 vccd1 vccd1 _1793_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_3_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1862_ hold195/X _1150_/X _1862_/S vssd1 vssd1 vccd1 vccd1 _1863_/B sky130_fd_sc_hd__mux2_1
XANTENNA__1026__A _1994_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1227_ _1441_/B _1227_/B _1458_/B vssd1 vssd1 vccd1 vccd1 _1228_/B sky130_fd_sc_hd__or3_4
X_1158_ _2116_/Q _1149_/B _1155_/Y _1467_/A _1157_/X vssd1 vssd1 vccd1 vccd1 _1158_/X
+ sky130_fd_sc_hd__a221o_1
X_1089_ hold61/X _1089_/B wire51/X _1089_/D vssd1 vssd1 vccd1 vccd1 _1174_/B sky130_fd_sc_hd__nand4b_4
XFILLER_0_7_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2061_ hold49/X _1519_/X _2066_/S vssd1 vssd1 vccd1 vccd1 hold50/A sky130_fd_sc_hd__mux2_1
X_2130_ _2150_/CLK _2130_/D vssd1 vssd1 vccd1 vccd1 _2130_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1914_ _1911_/Y _1912_/Y _1913_/X hold193/X _1912_/A vssd1 vssd1 vccd1 vccd1 _1914_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_44_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1845_ _1863_/A _1845_/B vssd1 vssd1 vccd1 vccd1 _2141_/D sky130_fd_sc_hd__and2_1
X_1776_ _1776_/A _1776_/B vssd1 vssd1 vccd1 vccd1 _1776_/X sky130_fd_sc_hd__or2_4
XFILLER_0_4_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1630_ _2111_/Q _1460_/A _1468_/A _1193_/X _1629_/X vssd1 vssd1 vccd1 vccd1 _1635_/S
+ sky130_fd_sc_hd__a221o_1
XANTENNA__1431__B2 _2112_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1561_ hold55/X _1511_/X _1567_/S vssd1 vssd1 vccd1 vccd1 hold56/A sky130_fd_sc_hd__mux2_1
X_1492_ _1492_/A _1651_/A vssd1 vssd1 vccd1 vccd1 _1492_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_39_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2113_ _2223_/CLK _2113_/D vssd1 vssd1 vccd1 vccd1 _2113_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_49_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2044_ _1873_/C _2043_/B _2031_/B _2043_/Y vssd1 vssd1 vccd1 vccd1 _2044_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_57_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1828_ _1828_/A _1828_/B _1828_/C _1828_/D vssd1 vssd1 vccd1 vccd1 _1829_/D sky130_fd_sc_hd__or4_1
X_1759_ _2115_/Q _1765_/B vssd1 vssd1 vccd1 vccd1 _1760_/D sky130_fd_sc_hd__nand2_1
XFILLER_0_25_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1868__B _1868_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2045__A _2057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1544_ _1540_/A _1539_/B _1539_/A vssd1 vssd1 vccd1 vccd1 _1547_/A sky130_fd_sc_hd__a21bo_1
X_1613_ _1625_/S vssd1 vssd1 vccd1 vccd1 _1617_/B sky130_fd_sc_hd__inv_2
XFILLER_0_41_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1475_ _1632_/A _1476_/C vssd1 vssd1 vccd1 vccd1 _1475_/Y sky130_fd_sc_hd__nor2_2
X_2027_ _1450_/A _2028_/B _2026_/Y _2000_/A vssd1 vssd1 vccd1 vccd1 _2027_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_60_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold240 _1402_/A vssd1 vssd1 vccd1 vccd1 _2077_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout74_A _1871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput8 io_in[24] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__clkbuf_1
X_1191_ hold13/A hold55/A _1882_/B vssd1 vssd1 vccd1 vccd1 _1191_/X sky130_fd_sc_hd__mux2_1
X_1260_ _1728_/B _1260_/B vssd1 vssd1 vccd1 vccd1 _1306_/B sky130_fd_sc_hd__and2_2
XFILLER_0_52_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1527_ _1548_/A _1868_/B vssd1 vssd1 vccd1 vccd1 _1527_/X sky130_fd_sc_hd__or2_1
X_1458_ _1458_/A _1458_/B _1826_/D _1994_/B vssd1 vssd1 vccd1 vccd1 _1460_/C sky130_fd_sc_hd__or4_1
X_1389_ _1389_/A _1389_/B vssd1 vssd1 vccd1 vccd1 _1404_/A sky130_fd_sc_hd__or2_1
XFILLER_0_60_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1174_ hold69/A _1174_/B _1174_/C vssd1 vssd1 vccd1 vccd1 _1174_/X sky130_fd_sc_hd__and3_1
X_1243_ _1994_/A _1243_/B vssd1 vssd1 vccd1 vccd1 _1243_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_47_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1312_ _1414_/A _1312_/B _1312_/C vssd1 vssd1 vccd1 vccd1 _1409_/A sky130_fd_sc_hd__or3_1
XFILLER_0_63_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1930_ hold102/X _1920_/Y _1929_/X _1871_/A vssd1 vssd1 vccd1 vccd1 _1930_/X sky130_fd_sc_hd__o211a_1
XANTENNA__1132__A _1135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput11 io_in[28] vssd1 vssd1 vccd1 vccd1 _1039_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_71_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1792_ _1792_/A _1792_/B _1792_/C _1792_/D vssd1 vssd1 vccd1 vccd1 _1792_/Y sky130_fd_sc_hd__nand4_1
XFILLER_0_24_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1764__B1 _1717_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1861_ _1863_/A _1861_/B vssd1 vssd1 vccd1 vccd1 _2149_/D sky130_fd_sc_hd__and2_1
X_1226_ _1421_/A _1455_/B vssd1 vssd1 vccd1 vccd1 _1458_/B sky130_fd_sc_hd__or2_1
X_1157_ hold178/X _1149_/C _1827_/B _1156_/X vssd1 vssd1 vccd1 vccd1 _1157_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_62_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1088_ _2179_/Q _1922_/B _1086_/X _1467_/B vssd1 vssd1 vccd1 vccd1 _1499_/A sky130_fd_sc_hd__a211o_4
XANTENNA__1916__S _1922_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1746__B1 _1717_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1210__A2 _1156_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2060_ hold13/X _1511_/X _2066_/S vssd1 vssd1 vccd1 vccd1 hold14/A sky130_fd_sc_hd__mux2_1
XFILLER_0_44_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1913_ _1913_/A _1913_/B vssd1 vssd1 vccd1 vccd1 _1913_/X sky130_fd_sc_hd__or2_1
XFILLER_0_29_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1844_ hold206/X _1211_/X _1862_/S vssd1 vssd1 vccd1 vccd1 _1845_/B sky130_fd_sc_hd__mux2_1
X_1775_ _1775_/A _1806_/B vssd1 vssd1 vccd1 vccd1 _1780_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_4_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2189_ _2201_/CLK _2189_/D vssd1 vssd1 vccd1 vccd1 _2189_/Q sky130_fd_sc_hd__dfxtp_1
X_1209_ _1545_/B _1828_/B _1150_/S hold116/X _1208_/X vssd1 vssd1 vccd1 vccd1 _1209_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__1500__A _2003_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_4_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _2223_/CLK sky130_fd_sc_hd__clkbuf_8
X_1560_ hold77/X _1503_/X _1567_/S vssd1 vssd1 vccd1 vccd1 hold78/A sky130_fd_sc_hd__mux2_1
XANTENNA__1195__B2 _1784_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2112_ _2223_/CLK _2112_/D vssd1 vssd1 vccd1 vccd1 _2112_/Q sky130_fd_sc_hd__dfxtp_4
X_1491_ _1491_/A _1491_/B vssd1 vssd1 vccd1 vccd1 _1651_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_39_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2043_ _2043_/A _2043_/B vssd1 vssd1 vccd1 vccd1 _2043_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_72_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1827_ _1827_/A _1827_/B _1827_/C vssd1 vssd1 vccd1 vccd1 _1828_/D sky130_fd_sc_hd__or3_1
XFILLER_0_29_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1689_ _1689_/A _1689_/B _1694_/A vssd1 vssd1 vccd1 vccd1 _1690_/B sky130_fd_sc_hd__or3_1
X_1758_ _2148_/Q _1776_/B _1717_/B vssd1 vssd1 vccd1 vccd1 _1760_/C sky130_fd_sc_hd__a21oi_1
XFILLER_0_4_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1543_ hold67/X _1501_/Y _1542_/X _1500_/B vssd1 vssd1 vccd1 vccd1 hold68/A sky130_fd_sc_hd__a22o_1
X_1474_ _1462_/Y _1474_/B vssd1 vssd1 vccd1 vccd1 _1632_/B sky130_fd_sc_hd__nand2b_1
X_1612_ _2121_/Q _1826_/D _1460_/Y _1866_/B vssd1 vssd1 vccd1 vccd1 _1625_/S sky130_fd_sc_hd__a22o_1
XFILLER_0_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2026_ _1945_/A _2021_/X _2028_/B vssd1 vssd1 vccd1 vccd1 _2026_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_72_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold241 _2171_/Q vssd1 vssd1 vccd1 vccd1 hold241/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1225__A _1548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold230 _2135_/Q vssd1 vssd1 vccd1 vccd1 hold230/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1937__A3 _1920_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1895__A _1922_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1834__S _1862_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput9 io_in[25] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__1135__A _1135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1190_ hold133/X _1149_/Y _1189_/X vssd1 vssd1 vccd1 vccd1 _1190_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_54_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1526_ hold43/X _1525_/X _1550_/S vssd1 vssd1 vccd1 vccd1 hold44/A sky130_fd_sc_hd__mux2_1
X_1457_ _1486_/A _1486_/D _1462_/B _1776_/A vssd1 vssd1 vccd1 vccd1 _1825_/C sky130_fd_sc_hd__or4_2
XFILLER_0_10_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1388_ _1420_/C _1407_/C _1410_/D _1388_/D vssd1 vssd1 vccd1 vccd1 _1401_/A sky130_fd_sc_hd__or4_1
X_2009_ _2009_/A _2028_/B vssd1 vssd1 vccd1 vccd1 _2009_/X sky130_fd_sc_hd__or2_1
XFILLER_0_18_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1311_ _1311_/A _1393_/B _1311_/C vssd1 vssd1 vccd1 vccd1 _1312_/C sky130_fd_sc_hd__and3_1
X_1242_ _1033_/Y _1229_/X _1238_/X _1241_/Y vssd1 vssd1 vccd1 vccd1 _1242_/X sky130_fd_sc_hd__a211o_1
X_1173_ _1751_/A _1149_/Y _1172_/X vssd1 vssd1 vccd1 vccd1 _1173_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_59_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1231__B1 _2057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1509_ _2111_/Q _1514_/B _1522_/B vssd1 vssd1 vccd1 vccd1 _1509_/Y sky130_fd_sc_hd__nor3_1
XFILLER_0_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1470__B1 _1871_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1525__A1 _1548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1773__A1 _2053_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1860_ hold178/X _1159_/X _1862_/S vssd1 vssd1 vccd1 vccd1 _1860_/X sky130_fd_sc_hd__mux2_1
Xinput12 io_in[29] vssd1 vssd1 vccd1 vccd1 _1941_/B sky130_fd_sc_hd__buf_1
XFILLER_0_71_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1791_ _1792_/B _1792_/C _1792_/D _1792_/A vssd1 vssd1 vccd1 vccd1 _1797_/A sky130_fd_sc_hd__a31o_1
XFILLER_0_24_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1156_ hold216/X _2097_/Q _1994_/A vssd1 vssd1 vccd1 vccd1 _1156_/X sky130_fd_sc_hd__mux2_4
X_1087_ _2179_/Q _1922_/B _1086_/X _1467_/B vssd1 vssd1 vccd1 vccd1 _1882_/A sky130_fd_sc_hd__a211oi_4
X_1225_ _1548_/A _1225_/B vssd1 vssd1 vccd1 vccd1 _1227_/B sky130_fd_sc_hd__nand2_4
XFILLER_0_62_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1989_ hold153/X _2031_/A _1988_/X _2049_/A vssd1 vssd1 vccd1 vccd1 _2185_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_65_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_4_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1842__S _1862_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1912_ _1912_/A _1912_/B vssd1 vssd1 vccd1 vccd1 _1912_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_44_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1843_ _1863_/A _1843_/B vssd1 vssd1 vccd1 vccd1 _2140_/D sky130_fd_sc_hd__and2_1
XFILLER_0_4_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1774_ _1132_/Y _1732_/B _1724_/C vssd1 vssd1 vccd1 vccd1 _1806_/B sky130_fd_sc_hd__a21o_2
XFILLER_0_4_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1208_ _1130_/B _1871_/B _1207_/X hold204/X vssd1 vssd1 vccd1 vccd1 _1208_/X sky130_fd_sc_hd__a22o_1
XANTENNA__1053__A _1548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2188_ _2219_/CLK _2188_/D vssd1 vssd1 vccd1 vccd1 _2188_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1139_ _1469_/A _1378_/C vssd1 vssd1 vccd1 vccd1 _1459_/C sky130_fd_sc_hd__or2_2
XFILLER_0_43_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1898__A _1918_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1490_ _1650_/B _1570_/A _1650_/A vssd1 vssd1 vccd1 vccd1 _1490_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_1_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1 hold1/A vssd1 vssd1 vccd1 vccd1 hold1/X sky130_fd_sc_hd__dlygate4sd3_1
X_2111_ _2208_/CLK _2111_/D vssd1 vssd1 vccd1 vccd1 _2111_/Q sky130_fd_sc_hd__dfxtp_2
X_2042_ _2049_/A _2042_/B vssd1 vssd1 vccd1 vccd1 _2202_/D sky130_fd_sc_hd__and2_1
XFILLER_0_39_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1826_ _1826_/A _1826_/B _1895_/B _1826_/D vssd1 vssd1 vccd1 vccd1 _1827_/C sky130_fd_sc_hd__or4_1
XFILLER_0_25_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1688_ _1689_/B _1694_/A _1689_/A vssd1 vssd1 vccd1 vccd1 _1697_/D sky130_fd_sc_hd__o21ai_1
X_1757_ _1757_/A _1763_/B vssd1 vssd1 vccd1 vccd1 _1760_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_48_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1611_ _1611_/A _1611_/B vssd1 vssd1 vccd1 vccd1 _1611_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_41_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1542_ _1542_/A _1542_/B vssd1 vssd1 vccd1 vccd1 _1542_/X sky130_fd_sc_hd__and2_1
X_1473_ _1462_/Y _1474_/B vssd1 vssd1 vccd1 vccd1 _1476_/C sky130_fd_sc_hd__and2b_2
XFILLER_0_34_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2025_ hold159/X _2028_/B _2024_/Y _2000_/A vssd1 vssd1 vccd1 vccd1 _2195_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_49_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold220 _2152_/Q vssd1 vssd1 vccd1 vccd1 hold220/X sky130_fd_sc_hd__dlygate4sd3_1
X_1809_ _1809_/A _1809_/B _1809_/C _1809_/D vssd1 vssd1 vccd1 vccd1 _1809_/Y sky130_fd_sc_hd__nand4_1
Xhold242 _2176_/Q vssd1 vssd1 vccd1 vccd1 hold93/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold231 _1832_/X vssd1 vssd1 vccd1 vccd1 _1833_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1850__S _1862_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1525_ _1548_/A _1796_/A _1523_/Y _1524_/X _1542_/A vssd1 vssd1 vccd1 vccd1 _1525_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_58_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1456_ _1456_/A _1921_/B vssd1 vssd1 vccd1 vccd1 _1994_/B sky130_fd_sc_hd__nand2_1
X_1387_ _1229_/C _1340_/B _1414_/D _1386_/X vssd1 vssd1 vccd1 vccd1 _1388_/D sky130_fd_sc_hd__a211o_1
XFILLER_0_10_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2008_ _2008_/A _2008_/B vssd1 vssd1 vccd1 vccd1 _2008_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_45_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_9_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1241_ _1241_/A _1241_/B vssd1 vssd1 vccd1 vccd1 _1241_/Y sky130_fd_sc_hd__nor2_1
X_1310_ _1279_/A _1285_/B _2015_/D _1313_/B vssd1 vssd1 vccd1 vccd1 _1311_/C sky130_fd_sc_hd__a31o_1
XFILLER_0_63_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1172_ hold171/X _1149_/B _1169_/X _1467_/A _1171_/X vssd1 vssd1 vccd1 vccd1 _1172_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_59_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1508_ _1514_/B _1522_/B _2111_/Q vssd1 vssd1 vccd1 vccd1 _1515_/A sky130_fd_sc_hd__o21a_1
X_1439_ _2124_/Q _1441_/B _1421_/X _2115_/Q _1423_/X vssd1 vssd1 vccd1 vccd1 _1439_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_69_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1930__C1 _1871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1525__A2 _1796_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput13 io_in[30] vssd1 vssd1 vccd1 vccd1 input13/X sky130_fd_sc_hd__buf_1
XFILLER_0_68_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1461__B2 _1871_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1790_ _1866_/B _1808_/B vssd1 vssd1 vccd1 vccd1 _1792_/D sky130_fd_sc_hd__nand2_1
XFILLER_0_24_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1224_ _1775_/A _1149_/Y _1223_/X vssd1 vssd1 vccd1 vccd1 _1224_/X sky130_fd_sc_hd__a21o_1
X_1155_ _1155_/A vssd1 vssd1 vccd1 vccd1 _1155_/Y sky130_fd_sc_hd__inv_2
X_1086_ hold79/A _1089_/B wire51/X _1089_/D vssd1 vssd1 vccd1 vccd1 _1086_/X sky130_fd_sc_hd__and4_2
XFILLER_0_47_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1988_ _1995_/A _1984_/C _2043_/B vssd1 vssd1 vccd1 vccd1 _1988_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_55_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1204__B2 _1864_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1514__A _2112_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1911_ _1913_/A _1913_/B vssd1 vssd1 vccd1 vccd1 _1911_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__1434__B2 _2164_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1842_ hold211/X _1213_/X _1862_/S vssd1 vssd1 vccd1 vccd1 _1843_/B sky130_fd_sc_hd__mux2_1
X_1773_ _2053_/B2 _1771_/Y _1780_/A _1820_/A2 hold125/X vssd1 vssd1 vccd1 vccd1 _1773_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_69_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2187_ _2219_/CLK _2187_/D vssd1 vssd1 vccd1 vccd1 _2187_/Q sky130_fd_sc_hd__dfxtp_1
X_1207_ _1716_/B _1459_/C _1895_/B vssd1 vssd1 vccd1 vccd1 _1207_/X sky130_fd_sc_hd__or3_4
XFILLER_0_19_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1138_ _1377_/A _1138_/B vssd1 vssd1 vccd1 vccd1 _1901_/S sky130_fd_sc_hd__or2_1
X_1069_ _1377_/B _1126_/A vssd1 vssd1 vccd1 vccd1 _1075_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_70_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1664__B2 _1796_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2 hold2/A vssd1 vssd1 vccd1 vccd1 hold2/X sky130_fd_sc_hd__dlygate4sd3_1
X_2110_ _2208_/CLK _2110_/D vssd1 vssd1 vccd1 vccd1 _2110_/Q sky130_fd_sc_hd__dfxtp_2
X_2041_ _1028_/A _2043_/B _1990_/Y _2036_/Y vssd1 vssd1 vccd1 vccd1 _2042_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_72_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1825_ _1825_/A _1825_/B _1825_/C _1825_/D vssd1 vssd1 vccd1 vccd1 _1828_/C sky130_fd_sc_hd__or4_1
XFILLER_0_32_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1756_ _2053_/B2 _1760_/A _1755_/Y _1820_/A2 _1751_/A vssd1 vssd1 vccd1 vccd1 _1756_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_25_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1687_ _1693_/A _1693_/B _1693_/C vssd1 vssd1 vccd1 vccd1 _1694_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_29_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1848__S _1862_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1610_ _2112_/Q _1460_/A _1609_/X vssd1 vssd1 vccd1 vccd1 _1611_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1541_ _1156_/X _1540_/Y _1548_/A vssd1 vssd1 vccd1 vccd1 _1542_/B sky130_fd_sc_hd__mux2_1
X_1472_ hold83/A _1829_/B vssd1 vssd1 vccd1 vccd1 _1474_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_5_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2024_ _2028_/B _2024_/B vssd1 vssd1 vccd1 vccd1 _2024_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__1331__B _2108_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2053__B2 _2053_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold221 _2154_/Q vssd1 vssd1 vccd1 vccd1 hold221/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold232 _2165_/Q vssd1 vssd1 vccd1 vccd1 hold232/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold243 _2200_/Q vssd1 vssd1 vccd1 vccd1 hold243/X sky130_fd_sc_hd__dlygate4sd3_1
X_1808_ _1808_/A _1808_/B vssd1 vssd1 vccd1 vccd1 _1809_/D sky130_fd_sc_hd__nand2_1
Xhold210 _1838_/X vssd1 vssd1 vccd1 vccd1 _1839_/B sky130_fd_sc_hd__dlygate4sd3_1
X_1739_ _2145_/Q _1776_/B _1738_/X vssd1 vssd1 vccd1 vccd1 _1742_/C sky130_fd_sc_hd__a21oi_1
XFILLER_0_25_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1524_ _1523_/A _1523_/B _1517_/A vssd1 vssd1 vccd1 vccd1 _1524_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_54_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1386_ _1033_/A _1241_/A _1296_/B _1119_/A vssd1 vssd1 vccd1 vccd1 _1386_/X sky130_fd_sc_hd__o211a_1
X_1455_ _1829_/A _1455_/B _1486_/D _1487_/A vssd1 vssd1 vccd1 vccd1 _1460_/A sky130_fd_sc_hd__or4_4
XFILLER_0_10_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2007_ _1923_/B _2019_/A _2006_/X _2000_/A vssd1 vssd1 vccd1 vccd1 _2007_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1234__C1 _1231_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1517__A _1517_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1252__A _1728_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1240_ _1033_/Y _1119_/A _1116_/C vssd1 vssd1 vccd1 vccd1 _1241_/B sky130_fd_sc_hd__a21oi_1
X_1171_ hold182/X _1149_/C _1827_/B _1868_/B vssd1 vssd1 vccd1 vccd1 _1171_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_59_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1507_ hold89/A _1546_/S vssd1 vssd1 vccd1 vccd1 _1522_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_42_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1438_ _2131_/Q _1227_/B _1228_/Y _1169_/X _1437_/X vssd1 vssd1 vccd1 vccd1 _1438_/X
+ sky130_fd_sc_hd__a221o_1
X_1369_ _1408_/A _1390_/C _1391_/B vssd1 vssd1 vccd1 vccd1 _1402_/B sky130_fd_sc_hd__or3_1
XFILLER_0_10_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1470__A2 _1776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold217_A _1156_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1758__B1 _1717_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2055__C_N _1941_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1461__A2 _1826_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput14 rst_n vssd1 vssd1 vccd1 vccd1 _1918_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__1856__S _1862_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1154_ _1499_/A _1151_/X _1152_/Y _1153_/Y vssd1 vssd1 vccd1 vccd1 _1155_/A sky130_fd_sc_hd__a2bb2o_1
X_1223_ _1130_/B _1864_/B _1222_/X _1467_/A vssd1 vssd1 vccd1 vccd1 _1223_/X sky130_fd_sc_hd__a211o_1
XANTENNA__1452__A2 _1776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1085_ _1085_/A _1486_/A _1825_/B _1079_/X vssd1 vssd1 vccd1 vccd1 _1089_/D sky130_fd_sc_hd__nor4b_4
X_1987_ _1033_/A _2031_/A _1986_/X _2057_/A vssd1 vssd1 vccd1 vccd1 _1987_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_15_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold167_A _2163_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1705__A _1921_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1910_ hold85/X hold91/X vssd1 vssd1 vccd1 vccd1 _1913_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_29_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output16_A _2160_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1841_ _1863_/A _1841_/B vssd1 vssd1 vccd1 vccd1 _2139_/D sky130_fd_sc_hd__and2_1
X_1772_ _1772_/A _1772_/B vssd1 vssd1 vccd1 vccd1 _1780_/A sky130_fd_sc_hd__or2_1
X_2186_ _2201_/CLK _2186_/D vssd1 vssd1 vccd1 vccd1 _2186_/Q sky130_fd_sc_hd__dfxtp_1
X_1137_ _1377_/A _1138_/B vssd1 vssd1 vccd1 vccd1 _1378_/C sky130_fd_sc_hd__nor2_2
X_1206_ hold139/X _1149_/Y _1205_/X vssd1 vssd1 vccd1 vccd1 _1206_/X sky130_fd_sc_hd__a21o_2
X_1068_ _2082_/Q _2081_/Q vssd1 vssd1 vccd1 vccd1 _1126_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_70_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1189__A1 _2112_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1260__A _1728_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1664__A2 _1826_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1352__A1 _1517_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3 hold3/A vssd1 vssd1 vccd1 vccd1 hold3/X sky130_fd_sc_hd__dlygate4sd3_1
X_2040_ _2049_/A _2040_/B vssd1 vssd1 vccd1 vccd1 _2201_/D sky130_fd_sc_hd__and2_1
XFILLER_0_72_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1812__C1 _1717_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1686_ _1689_/B _1686_/B vssd1 vssd1 vccd1 vccd1 _1693_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_40_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1824_ _1824_/A _1922_/B _1823_/X vssd1 vssd1 vccd1 vccd1 _1825_/D sky130_fd_sc_hd__or3b_1
X_1755_ _1755_/A _1755_/B _1755_/C _1755_/D vssd1 vssd1 vccd1 vccd1 _1755_/Y sky130_fd_sc_hd__nand4_1
XFILLER_0_25_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2169_ _2182_/CLK _2169_/D vssd1 vssd1 vccd1 vccd1 _2169_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1239__B _1239_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1540_ _1540_/A _1540_/B vssd1 vssd1 vccd1 vccd1 _1540_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_54_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1471_ _2117_/Q _1460_/A _1468_/A _1096_/X _1470_/X vssd1 vssd1 vccd1 vccd1 _1476_/B
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_5_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2023_ hold83/X _1923_/B _2022_/X _2003_/A vssd1 vssd1 vccd1 vccd1 hold84/A sky130_fd_sc_hd__a211o_1
XANTENNA__2038__C1 _2057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1807_ _2115_/Q _1135_/A _1776_/X _2140_/Q _1717_/B vssd1 vssd1 vccd1 vccd1 _1809_/C
+ sky130_fd_sc_hd__a221oi_2
XFILLER_0_9_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold222 _2157_/Q vssd1 vssd1 vccd1 vccd1 hold222/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold233 _1917_/X vssd1 vssd1 vccd1 vccd1 _1918_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold244 _2189_/Q vssd1 vssd1 vccd1 vccd1 hold244/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold200 _2112_/Q vssd1 vssd1 vccd1 vccd1 hold200/X sky130_fd_sc_hd__dlygate4sd3_1
X_1669_ _1669_/A _1669_/B vssd1 vssd1 vccd1 vccd1 _1669_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_40_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold211 _2140_/Q vssd1 vssd1 vccd1 vccd1 hold211/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_4_3_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _2209_/CLK sky130_fd_sc_hd__clkbuf_8
X_1738_ _1025_/Y hold93/X _1455_/B vssd1 vssd1 vccd1 vccd1 _1738_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_25_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1523_ _1523_/A _1523_/B vssd1 vssd1 vccd1 vccd1 _1523_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__1546__A1 _2117_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1454_ _2009_/A _1829_/B vssd1 vssd1 vccd1 vccd1 _1654_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_10_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1385_ _1486_/B _1365_/A _1403_/A2 _1826_/B vssd1 vssd1 vccd1 vccd1 _1414_/D sky130_fd_sc_hd__a22o_1
X_2006_ _2006_/A _2028_/B vssd1 vssd1 vccd1 vccd1 _2006_/X sky130_fd_sc_hd__or2_1
XFILLER_0_45_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1517__B _1866_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1708__A _1921_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1170_ hold212/X hold96/X _1994_/A vssd1 vssd1 vccd1 vccd1 _1868_/B sky130_fd_sc_hd__mux2_4
XFILLER_0_47_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1506_ _2188_/Q _2151_/Q vssd1 vssd1 vccd1 vccd1 _1546_/S sky130_fd_sc_hd__nand2b_1
X_1437_ _2123_/Q _1441_/B _1421_/X _2114_/Q _1436_/X vssd1 vssd1 vccd1 vccd1 _1437_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_2_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1299_ _1299_/A _1336_/B _1299_/C vssd1 vssd1 vccd1 vccd1 _1300_/C sky130_fd_sc_hd__and3_1
X_1368_ _1408_/B _1413_/A _1407_/B vssd1 vssd1 vccd1 vccd1 _1391_/B sky130_fd_sc_hd__or3_1
XANTENNA_clkbuf_4_13_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1153_ hold67/A _1499_/B _1882_/A vssd1 vssd1 vccd1 vccd1 _1153_/Y sky130_fd_sc_hd__a21oi_1
X_1084_ _1084_/A _1141_/B vssd1 vssd1 vccd1 vccd1 _1486_/A sky130_fd_sc_hd__nor2_2
X_1222_ _2110_/Q _1828_/B _1207_/X _2135_/Q _1130_/A vssd1 vssd1 vccd1 vccd1 _1222_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_59_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1986_ _1980_/A _2001_/C _1973_/A _2043_/B vssd1 vssd1 vccd1 vccd1 _1986_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_70_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1530__B _2108_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1258__A _1728_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1840_ hold207/X _1215_/X _1862_/S vssd1 vssd1 vccd1 vccd1 _1840_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_29_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1771_ _1772_/A _1772_/B vssd1 vssd1 vccd1 vccd1 _1771_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2185_ _2201_/CLK _2185_/D vssd1 vssd1 vccd1 vccd1 _2185_/Q sky130_fd_sc_hd__dfxtp_1
X_1136_ _1377_/A _1136_/B vssd1 vssd1 vccd1 vccd1 _1469_/A sky130_fd_sc_hd__nor2_1
X_1205_ hold175/X _1149_/B _1202_/Y _1467_/A _1204_/X vssd1 vssd1 vccd1 vccd1 _1205_/X
+ sky130_fd_sc_hd__a221o_1
X_1067_ _1821_/A _2079_/Q _2078_/Q _2077_/Q vssd1 vssd1 vccd1 vccd1 _1377_/B sky130_fd_sc_hd__or4_2
XFILLER_0_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1969_ hold202/X _1923_/B _2003_/A vssd1 vssd1 vccd1 vccd1 _1969_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_50_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4 hold4/A vssd1 vssd1 vccd1 vccd1 hold4/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1823_ _2082_/Q _2081_/Q _1822_/X vssd1 vssd1 vccd1 vccd1 _1823_/X sky130_fd_sc_hd__a21o_1
X_1685_ _1582_/B _1582_/C _1582_/A vssd1 vssd1 vccd1 vccd1 _1686_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_40_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1754_ _1755_/B _1755_/C _1755_/D _1755_/A vssd1 vssd1 vccd1 vccd1 _1760_/A sky130_fd_sc_hd__a31o_1
XFILLER_0_25_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2168_ _2214_/CLK hold4/X vssd1 vssd1 vccd1 vccd1 hold3/A sky130_fd_sc_hd__dfxtp_1
X_2099_ _2214_/CLK hold78/X vssd1 vssd1 vccd1 vccd1 hold77/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1119_ _1119_/A _1716_/A vssd1 vssd1 vccd1 vccd1 _1828_/A sky130_fd_sc_hd__or2_1
XFILLER_0_63_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_300 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1470_ _2142_/Q _1776_/A _1871_/B _1469_/X vssd1 vssd1 vccd1 vccd1 _1470_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_1_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2022_ _2043_/A _2001_/C _2024_/B _2031_/A vssd1 vssd1 vccd1 vccd1 _2022_/X sky130_fd_sc_hd__o31a_1
XFILLER_0_9_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1806_ _1806_/A _1806_/B vssd1 vssd1 vccd1 vccd1 _1809_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_31_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold201 _2144_/Q vssd1 vssd1 vccd1 vccd1 hold201/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_17_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold223 _1808_/A vssd1 vssd1 vccd1 vccd1 _1869_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold212 _2156_/Q vssd1 vssd1 vccd1 vccd1 hold212/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold245 _2166_/Q vssd1 vssd1 vccd1 vccd1 hold245/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold234 _2162_/Q vssd1 vssd1 vccd1 vccd1 hold234/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1668_ _1632_/A _1666_/X _1667_/Y _1475_/Y vssd1 vssd1 vccd1 vccd1 _1668_/X sky130_fd_sc_hd__a211o_1
X_1599_ _1632_/A _1603_/B _1595_/X vssd1 vssd1 vccd1 vccd1 _1599_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1737_ _1732_/B _1724_/C hold133/X vssd1 vssd1 vccd1 vccd1 _1742_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_0_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1266__A _1728_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1522_ _2113_/Q _1522_/B vssd1 vssd1 vccd1 vccd1 _1523_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_50_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1453_ _2009_/A _1829_/B vssd1 vssd1 vccd1 vccd1 _1697_/A sky130_fd_sc_hd__and2_2
XFILLER_0_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2005_ _2005_/A _2005_/B vssd1 vssd1 vccd1 vccd1 _2019_/A sky130_fd_sc_hd__nor2_1
X_1384_ _1128_/A _1365_/A _1403_/A2 _1116_/C _1405_/C vssd1 vssd1 vccd1 vccd1 _1410_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_26_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1528__A2 _1517_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output39_A _2162_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1505_ _2188_/Q _2151_/Q hold89/A vssd1 vssd1 vccd1 vccd1 _1514_/B sky130_fd_sc_hd__and3_1
XFILLER_0_56_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1436_ _1025_/Y _1039_/Y _1455_/B _1421_/A _2205_/Q vssd1 vssd1 vccd1 vccd1 _1436_/X
+ sky130_fd_sc_hd__a32o_1
X_1367_ _1776_/A _1403_/A2 _1365_/X _1414_/C vssd1 vssd1 vccd1 vccd1 _1390_/C sky130_fd_sc_hd__a211o_1
XFILLER_0_2_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1298_ _1996_/A _2001_/B _1360_/C _1317_/B vssd1 vssd1 vccd1 vccd1 _1299_/C sky130_fd_sc_hd__o211a_1
XFILLER_0_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_328 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1221_ hold177/X _1828_/B _1150_/S hold98/X _1220_/X vssd1 vssd1 vccd1 vccd1 _1221_/X
+ sky130_fd_sc_hd__a221o_2
X_1152_ hold47/A _1882_/B vssd1 vssd1 vccd1 vccd1 _1152_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_59_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1083_ _1345_/A _1080_/B _1102_/B _1344_/A vssd1 vssd1 vccd1 vccd1 _1825_/B sky130_fd_sc_hd__o22ai_4
X_1985_ _1239_/A _2028_/B _1978_/B _1984_/X _2000_/A vssd1 vssd1 vccd1 vccd1 _1985_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_7_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1419_ _1419_/A _1419_/B vssd1 vssd1 vccd1 vccd1 _1420_/D sky130_fd_sc_hd__or2_1
Xwire51 wire51/A vssd1 vssd1 vccd1 vccd1 wire51/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_21_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1770_ hold125/X _1763_/B _1769_/X vssd1 vssd1 vccd1 vccd1 _1772_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__1912__A _1912_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2184_ _2210_/CLK _2184_/D vssd1 vssd1 vccd1 vccd1 _2184_/Q sky130_fd_sc_hd__dfxtp_1
X_1204_ hold176/X _1149_/C _1827_/B _1864_/B vssd1 vssd1 vccd1 vccd1 _1204_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
X_1135_ _1135_/A _1238_/B _1229_/C vssd1 vssd1 vccd1 vccd1 _1828_/B sky130_fd_sc_hd__or3_4
X_1066_ _1821_/A _1236_/D _1114_/B vssd1 vssd1 vccd1 vccd1 _1826_/A sky130_fd_sc_hd__nor3_1
XFILLER_0_62_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1968_ _1995_/A _2001_/C _1984_/C _1964_/Y _1967_/Y vssd1 vssd1 vccd1 vccd1 _1968_/X
+ sky130_fd_sc_hd__a311o_1
X_1899_ _1903_/B _1378_/C _1881_/X _1071_/Y _1912_/A vssd1 vssd1 vccd1 vccd1 _1899_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_0_43_353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1594__B1 _1868_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1269__A _1728_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5 hold5/A vssd1 vssd1 vccd1 vccd1 hold5/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1753_ _2114_/Q _1765_/B vssd1 vssd1 vccd1 vccd1 _1755_/D sky130_fd_sc_hd__nand2_1
X_1822_ _1245_/B _1821_/X _1345_/B _1106_/A vssd1 vssd1 vccd1 vccd1 _1822_/X sky130_fd_sc_hd__o211a_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1684_ _1691_/A _1708_/B _1691_/C vssd1 vssd1 vccd1 vccd1 _1693_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_40_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2167_ _2182_/CLK hold95/X vssd1 vssd1 vccd1 vccd1 _2167_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2098_ _2182_/CLK _2098_/D vssd1 vssd1 vccd1 vccd1 _2098_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2056__A1 _1025_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1049_ _1821_/A _1114_/B _1821_/B _1236_/D vssd1 vssd1 vccd1 vccd1 _1338_/A sky130_fd_sc_hd__or4bb_4
XFILLER_0_35_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1118_ _1245_/A _2081_/Q _1131_/C vssd1 vssd1 vccd1 vccd1 _1716_/A sky130_fd_sc_hd__and3_1
XFILLER_0_43_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2021_ _2043_/A _2008_/B _2024_/B vssd1 vssd1 vccd1 vccd1 _2021_/X sky130_fd_sc_hd__o21a_1
XANTENNA__1462__A _1922_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold224 _2153_/Q vssd1 vssd1 vccd1 vccd1 hold224/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold202 _2179_/Q vssd1 vssd1 vccd1 vccd1 hold202/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold235 _1897_/X vssd1 vssd1 vccd1 vccd1 _1898_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold213 _2202_/Q vssd1 vssd1 vccd1 vccd1 _1028_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_1805_ _2053_/B2 _1809_/A _1804_/Y _1820_/A2 _1800_/A vssd1 vssd1 vccd1 vccd1 _1805_/X
+ sky130_fd_sc_hd__a32o_1
X_1736_ _1734_/X _1735_/Y _1732_/A _1820_/A2 vssd1 vssd1 vccd1 vccd1 _1736_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_25_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1667_ _1622_/A _1622_/B _1669_/B _1632_/B vssd1 vssd1 vccd1 vccd1 _1667_/Y sky130_fd_sc_hd__a211oi_1
X_1598_ _1476_/C _1595_/X _1603_/B _1475_/Y vssd1 vssd1 vccd1 vccd1 _1598_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2219_ _2219_/CLK hold38/X vssd1 vssd1 vccd1 vccd1 hold37/A sky130_fd_sc_hd__dfxtp_1
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1712__A0 _1545_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1521_ _2112_/Q _1514_/B _1515_/X vssd1 vssd1 vccd1 vccd1 _1523_/A sky130_fd_sc_hd__a21o_1
X_1452_ _2107_/Q _1776_/A _1829_/B _2195_/Q _1228_/B vssd1 vssd1 vccd1 vccd1 _1650_/B
+ sky130_fd_sc_hd__a221o_2
X_1383_ _1100_/Y _1415_/A3 _1340_/B _1458_/A vssd1 vssd1 vccd1 vccd1 _1405_/C sky130_fd_sc_hd__a22o_1
XFILLER_0_22_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1920__A _1920_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2004_ _1255_/Y _2015_/B _1960_/B _1996_/A _1995_/A vssd1 vssd1 vccd1 vccd1 _2005_/B
+ sky130_fd_sc_hd__o32a_1
XFILLER_0_42_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1942__B1 _2003_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1719_ _1732_/B _1724_/C hold139/X vssd1 vssd1 vccd1 vccd1 _1726_/A sky130_fd_sc_hd__o21a_1
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1830__A _1921_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1740__A _2112_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1216__A2 _1796_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1504_ hold65/X _1503_/X _1550_/S vssd1 vssd1 vccd1 vccd1 hold66/A sky130_fd_sc_hd__mux2_1
XANTENNA__1924__B1 _2003_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1435_ _1177_/X _1228_/Y _1422_/Y _2113_/Q _1434_/X vssd1 vssd1 vccd1 vccd1 _1435_/X
+ sky130_fd_sc_hd__a221o_1
X_1366_ _1824_/A _1365_/A _1403_/A2 _1486_/D vssd1 vssd1 vccd1 vccd1 _1414_/C sky130_fd_sc_hd__a22o_1
XFILLER_0_10_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1297_ _1297_/A _2015_/A vssd1 vssd1 vccd1 vccd1 _1317_/B sky130_fd_sc_hd__or2_1
XFILLER_0_73_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1151_ hold19/A hold29/A _1499_/B vssd1 vssd1 vccd1 vccd1 _1151_/X sky130_fd_sc_hd__mux2_1
X_1220_ _1130_/B _1865_/B _1207_/X hold227/X vssd1 vssd1 vccd1 vccd1 _1220_/X sky130_fd_sc_hd__a22o_1
XANTENNA__1382__A1 _1922_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1082_ _1344_/A _1102_/B vssd1 vssd1 vccd1 vccd1 _1903_/B sky130_fd_sc_hd__nor2_2
X_1984_ _2015_/C _1984_/B _1984_/C vssd1 vssd1 vccd1 vccd1 _1984_/X sky130_fd_sc_hd__and3_1
XFILLER_0_55_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1418_ _1418_/A _1418_/B _1418_/C _1418_/D vssd1 vssd1 vccd1 vccd1 _1419_/B sky130_fd_sc_hd__or4_1
X_1349_ _1390_/B _1406_/A _1411_/A _1349_/D vssd1 vssd1 vccd1 vccd1 _1350_/D sky130_fd_sc_hd__or4_1
XFILLER_0_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1203_ hold220/X hold94/X _1994_/A vssd1 vssd1 vccd1 vccd1 _1864_/B sky130_fd_sc_hd__mux2_4
X_2183_ _2219_/CLK _2183_/D vssd1 vssd1 vccd1 vccd1 _2183_/Q sky130_fd_sc_hd__dfxtp_1
X_1134_ _1344_/A _1138_/B vssd1 vssd1 vccd1 vccd1 _1229_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_18_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1065_ _1345_/A _1136_/B vssd1 vssd1 vccd1 vccd1 _1128_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1967_ _1948_/B _1951_/Y _2005_/A vssd1 vssd1 vccd1 vccd1 _1967_/Y sky130_fd_sc_hd__a21oi_1
X_1898_ _1918_/A _1898_/B vssd1 vssd1 vccd1 vccd1 _2162_/D sky130_fd_sc_hd__and2_1
XFILLER_0_50_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1585__B2 _1808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6 hold6/A vssd1 vssd1 vccd1 vccd1 hold6/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_71_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1812__A2 _1135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1683_ _1693_/A _1683_/B vssd1 vssd1 vccd1 vccd1 _1691_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_40_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1752_ _2147_/Q _1776_/B _1717_/B vssd1 vssd1 vccd1 vccd1 _1755_/C sky130_fd_sc_hd__a21oi_1
X_1821_ _1821_/A _1821_/B _1236_/D vssd1 vssd1 vccd1 vccd1 _1821_/X sky130_fd_sc_hd__or3b_1
XFILLER_0_20_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2097_ _2172_/CLK _2097_/D vssd1 vssd1 vccd1 vccd1 _2097_/Q sky130_fd_sc_hd__dfxtp_1
X_2166_ _2214_/CLK _2166_/D vssd1 vssd1 vccd1 vccd1 _2166_/Q sky130_fd_sc_hd__dfxtp_2
X_1117_ _1344_/A _1136_/B vssd1 vssd1 vccd1 vccd1 _1119_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_63_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1264__A0 _1808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1048_ _1084_/A _1106_/A vssd1 vssd1 vccd1 vccd1 _1548_/A sky130_fd_sc_hd__or2_4
XFILLER_0_0_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1833__A _1863_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2020_ _2005_/A _2016_/X _2019_/Y vssd1 vssd1 vccd1 vccd1 _2024_/B sky130_fd_sc_hd__o21a_1
XANTENNA__1918__A _1918_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold225 _1784_/A vssd1 vssd1 vccd1 vccd1 _1865_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__1549__A1 _1548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold203 _2192_/Q vssd1 vssd1 vccd1 vccd1 hold203/X sky130_fd_sc_hd__dlygate4sd3_1
X_1666_ _1622_/A _1622_/B _1669_/B vssd1 vssd1 vccd1 vccd1 _1666_/X sky130_fd_sc_hd__a21o_1
Xhold236 _2160_/Q vssd1 vssd1 vccd1 vccd1 hold236/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold214 _2164_/Q vssd1 vssd1 vccd1 vccd1 hold214/X sky130_fd_sc_hd__dlygate4sd3_1
X_1804_ _1804_/A _1804_/B _1804_/C _1804_/D vssd1 vssd1 vccd1 vccd1 _1804_/Y sky130_fd_sc_hd__nand4_1
X_1735_ _1735_/A _1742_/A vssd1 vssd1 vccd1 vccd1 _1735_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_25_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1597_ _1595_/X _1603_/B _1669_/A vssd1 vssd1 vccd1 vccd1 _1597_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__1075__D _1922_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2218_ _2226_/CLK hold46/X vssd1 vssd1 vccd1 vccd1 hold45/A sky130_fd_sc_hd__dfxtp_1
X_2149_ _2150_/CLK _2149_/D vssd1 vssd1 vccd1 vccd1 _2149_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1520_ hold75/X _1501_/Y _1519_/X _1500_/B vssd1 vssd1 vccd1 vccd1 hold76/A sky130_fd_sc_hd__a22o_1
XFILLER_0_42_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1451_ _2107_/Q _1776_/A _1829_/B _2195_/Q _1228_/B vssd1 vssd1 vccd1 vccd1 _1491_/B
+ sky130_fd_sc_hd__a221oi_4
X_1382_ _1922_/B _1340_/B _1381_/X _1415_/A3 vssd1 vssd1 vccd1 vccd1 _1407_/C sky130_fd_sc_hd__a22o_1
XANTENNA__1920__B _1920_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2003_ _2003_/A _2003_/B vssd1 vssd1 vccd1 vccd1 _2189_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_9_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1649_ _1697_/A _1635_/S _1647_/X _1648_/Y vssd1 vssd1 vccd1 vccd1 _1653_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_41_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1718_ _1922_/B _1728_/B vssd1 vssd1 vccd1 vccd1 _1724_/C sky130_fd_sc_hd__and2_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_2_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _2164_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_67_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1503_ _2110_/Q _1517_/A _1542_/A _1502_/X vssd1 vssd1 vccd1 vccd1 _1503_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_50_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1296_ _1922_/B _1296_/B vssd1 vssd1 vccd1 vccd1 _1393_/A sky130_fd_sc_hd__nand2_2
X_1434_ _2130_/Q _1227_/B _1423_/X _2164_/Q _1433_/X vssd1 vssd1 vccd1 vccd1 _1434_/X
+ sky130_fd_sc_hd__a221o_1
X_1365_ _1365_/A _1826_/D _1365_/C vssd1 vssd1 vccd1 vccd1 _1365_/X sky130_fd_sc_hd__and3_1
XFILLER_0_53_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout63_A _2053_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1841__A _1863_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1906__A1 hold194/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1150_ _1148_/X hold125/X _1150_/S vssd1 vssd1 vccd1 vccd1 _1150_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1081_ _1236_/D _1114_/B _1821_/B _1821_/A vssd1 vssd1 vccd1 vccd1 _1102_/B sky130_fd_sc_hd__nand4b_4
XFILLER_0_7_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1983_ _1923_/B _1980_/X _1981_/X _1982_/X _1871_/A vssd1 vssd1 vccd1 vccd1 _1983_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_2_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1417_ _1417_/A _1417_/B _1417_/C _1417_/D vssd1 vssd1 vccd1 vccd1 _1418_/D sky130_fd_sc_hd__or4_1
XFILLER_0_2_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1279_ _1279_/A _1287_/B vssd1 vssd1 vccd1 vccd1 _1279_/Y sky130_fd_sc_hd__nor2_1
X_1348_ _1123_/C _1403_/A2 _1346_/X _1415_/A3 _1389_/B vssd1 vssd1 vccd1 vccd1 _1349_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_73_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2182_ _2182_/CLK _2182_/D vssd1 vssd1 vccd1 vccd1 _2182_/Q sky130_fd_sc_hd__dfxtp_1
X_1202_ _1202_/A _1202_/B vssd1 vssd1 vccd1 vccd1 _1202_/Y sky130_fd_sc_hd__nand2_1
X_1064_ _2080_/Q _1236_/D _1114_/B _1821_/B vssd1 vssd1 vccd1 vccd1 _1136_/B sky130_fd_sc_hd__or4bb_2
X_1133_ _1345_/A _1338_/A vssd1 vssd1 vccd1 vccd1 _1238_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_18_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1966_ _1923_/B _1964_/Y _1965_/X _2000_/A vssd1 vssd1 vccd1 vccd1 _2178_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_47_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1897_ _1896_/X hold234/X _1897_/S vssd1 vssd1 vccd1 vccd1 _1897_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_50_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1594__A2 _1776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1585__A2 _1826_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold7 hold7/A vssd1 vssd1 vccd1 vccd1 hold7/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_71_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1820_ hold116/X _1820_/A2 _1819_/Y _2053_/B2 vssd1 vssd1 vccd1 vccd1 _1820_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_29_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1682_ _1593_/B _1593_/C _1593_/A vssd1 vssd1 vccd1 vccd1 _1683_/B sky130_fd_sc_hd__a21oi_1
X_1751_ _1751_/A _1763_/B vssd1 vssd1 vccd1 vccd1 _1755_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_20_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2096_ _2172_/CLK _2096_/D vssd1 vssd1 vccd1 vccd1 _2096_/Q sky130_fd_sc_hd__dfxtp_1
X_2165_ _2208_/CLK _2165_/D vssd1 vssd1 vccd1 vccd1 _2165_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_45_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1116_ _1238_/A _1723_/A _1116_/C vssd1 vssd1 vccd1 vccd1 _1123_/A sky130_fd_sc_hd__or3_1
X_1047_ _1345_/A _1106_/A vssd1 vssd1 vccd1 vccd1 _1517_/A sky130_fd_sc_hd__nor2_4
XFILLER_0_71_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_15_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _2172_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_63_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1949_ _2015_/C _1281_/Y _1984_/C _1948_/Y vssd1 vssd1 vccd1 vccd1 _1978_/A sky130_fd_sc_hd__a31o_1
XFILLER_0_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1296__A _1922_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1246__B2 _1448_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1803_ _1804_/B _1804_/C _1804_/D _1804_/A vssd1 vssd1 vccd1 vccd1 _1809_/A sky130_fd_sc_hd__a31o_1
XANTENNA__1549__A2 _1871_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold226 _2159_/Q vssd1 vssd1 vccd1 vccd1 hold226/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold215 _1999_/X vssd1 vssd1 vccd1 vccd1 _2000_/B sky130_fd_sc_hd__dlygate4sd3_1
X_1665_ _1673_/S vssd1 vssd1 vccd1 vccd1 _1669_/B sky130_fd_sc_hd__inv_2
Xhold237 _1879_/X vssd1 vssd1 vccd1 vccd1 _1880_/B sky130_fd_sc_hd__dlygate4sd3_1
X_1596_ _2123_/Q _1826_/D _1460_/Y _1868_/B vssd1 vssd1 vccd1 vccd1 _1603_/B sky130_fd_sc_hd__a22o_1
Xhold204 _2142_/Q vssd1 vssd1 vccd1 vccd1 hold204/X sky130_fd_sc_hd__dlygate4sd3_1
X_1734_ _1734_/A _1734_/B _1734_/C _1734_/D vssd1 vssd1 vccd1 vccd1 _1734_/X sky130_fd_sc_hd__and4_1
XFILLER_0_21_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2217_ _2225_/CLK hold30/X vssd1 vssd1 vccd1 vccd1 hold29/A sky130_fd_sc_hd__dfxtp_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1485__A1 _1448_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2079_ _2164_/CLK _2079_/D vssd1 vssd1 vccd1 vccd1 _2079_/Q sky130_fd_sc_hd__dfxtp_1
X_2148_ _2150_/CLK _2148_/D vssd1 vssd1 vccd1 vccd1 _2148_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1450_ _1450_/A _1829_/B vssd1 vssd1 vccd1 vccd1 _1491_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_35_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1381_ _1826_/D _1364_/Y _1378_/X _1724_/B vssd1 vssd1 vccd1 vccd1 _1381_/X sky130_fd_sc_hd__a211o_1
X_2002_ _1874_/B _2043_/B _2001_/X vssd1 vssd1 vccd1 vccd1 _2003_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1648_ _1697_/C _1652_/S _1654_/A vssd1 vssd1 vccd1 vccd1 _1648_/Y sky130_fd_sc_hd__o21ai_1
X_1579_ _1697_/A _1476_/B _1576_/X _1578_/Y vssd1 vssd1 vccd1 vccd1 _1582_/A sky130_fd_sc_hd__a22o_1
X_1717_ _1922_/B _1717_/B _1765_/B vssd1 vssd1 vccd1 vccd1 _1732_/B sky130_fd_sc_hd__nor3_2
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1839__A _1863_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_0_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1502_ _1548_/A _1864_/B vssd1 vssd1 vccd1 vccd1 _1502_/X sky130_fd_sc_hd__or2_1
X_1433_ _2122_/Q _1441_/B vssd1 vssd1 vccd1 vccd1 _1433_/X sky130_fd_sc_hd__and2_1
X_1295_ _1881_/A _1296_/B vssd1 vssd1 vccd1 vccd1 _1360_/C sky130_fd_sc_hd__and2_1
X_1364_ _1365_/C vssd1 vssd1 vccd1 vccd1 _1364_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_73_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1915__A2 _1922_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1612__B2 _1866_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output37_A _2163_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1080_ _1345_/A _1080_/B vssd1 vssd1 vccd1 vccd1 _1458_/A sky130_fd_sc_hd__nor2_2
X_1982_ _1982_/A _2028_/B vssd1 vssd1 vccd1 vccd1 _1982_/X sky130_fd_sc_hd__or2_1
XFILLER_0_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1416_ _1416_/A _1416_/B _1416_/C _1416_/D vssd1 vssd1 vccd1 vccd1 _1418_/C sky130_fd_sc_hd__or4_1
X_1347_ _1044_/X _1245_/C _1340_/B _1458_/A _1415_/A3 vssd1 vssd1 vccd1 vccd1 _1389_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_2_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1278_ _2015_/B _1278_/B vssd1 vssd1 vccd1 vccd1 _1287_/B sky130_fd_sc_hd__or2_1
XFILLER_0_38_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1201_ hold37/A _1499_/B _1199_/X _1499_/A vssd1 vssd1 vccd1 vccd1 _1202_/B sky130_fd_sc_hd__o211ai_2
XFILLER_0_20_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2181_ _2219_/CLK hold80/X vssd1 vssd1 vccd1 vccd1 hold79/A sky130_fd_sc_hd__dfxtp_1
X_1063_ _1143_/A _1141_/B _1344_/A vssd1 vssd1 vccd1 vccd1 _1825_/A sky130_fd_sc_hd__a21oi_1
X_1132_ _1135_/A vssd1 vssd1 vccd1 vccd1 _1132_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_18_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1965_ _1965_/A _2028_/B vssd1 vssd1 vccd1 vccd1 _1965_/X sky130_fd_sc_hd__or2_1
XFILLER_0_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1896_ _1545_/B _1871_/B _1896_/S vssd1 vssd1 vccd1 vccd1 _1896_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_43_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1847__A _1863_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold8 hold8/A vssd1 vssd1 vccd1 vccd1 hold8/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1750_ _2053_/B2 _1755_/A _1749_/Y _1820_/A2 _1745_/A vssd1 vssd1 vccd1 vccd1 _1750_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_52_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1681_ _1680_/A _1680_/B _1705_/B _1707_/A vssd1 vssd1 vccd1 vccd1 _1708_/B sky130_fd_sc_hd__o31a_1
XFILLER_0_40_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2164_ _2164_/CLK _2164_/D vssd1 vssd1 vccd1 vccd1 _2164_/Q sky130_fd_sc_hd__dfxtp_2
X_2095_ _2172_/CLK _2095_/D vssd1 vssd1 vccd1 vccd1 hold96/A sky130_fd_sc_hd__dfxtp_1
X_1115_ _1345_/A _1138_/B vssd1 vssd1 vccd1 vccd1 _1116_/C sky130_fd_sc_hd__nor2_2
X_1046_ _1236_/D _1821_/B _1114_/B _1821_/A vssd1 vssd1 vccd1 vccd1 _1106_/A sky130_fd_sc_hd__or4bb_4
XFILLER_0_63_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1948_ _2005_/A _1948_/B vssd1 vssd1 vccd1 vccd1 _1948_/Y sky130_fd_sc_hd__nor2_1
X_1879_ hold236/X _1878_/X _1879_/S vssd1 vssd1 vccd1 vccd1 _1879_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_16_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_5_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1802_ _1868_/B _1808_/B vssd1 vssd1 vccd1 vccd1 _1804_/D sky130_fd_sc_hd__nand2_1
X_1733_ _1734_/B _1734_/C _1734_/D _1734_/A vssd1 vssd1 vccd1 vccd1 _1742_/A sky130_fd_sc_hd__a31o_1
Xhold216 _2158_/Q vssd1 vssd1 vccd1 vccd1 hold216/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1595_ _2114_/Q _1460_/A _1468_/A _1169_/X _1594_/X vssd1 vssd1 vccd1 vccd1 _1595_/X
+ sky130_fd_sc_hd__a221o_1
X_1664_ _2122_/Q _1826_/D _1460_/Y _1796_/A vssd1 vssd1 vccd1 vccd1 _1673_/S sky130_fd_sc_hd__a22o_1
Xhold205 _1846_/X vssd1 vssd1 vccd1 vccd1 _1847_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold238 _2082_/Q vssd1 vssd1 vccd1 vccd1 _1040_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold227 _2136_/Q vssd1 vssd1 vccd1 vccd1 hold227/X sky130_fd_sc_hd__dlygate4sd3_1
X_2216_ _2226_/CLK hold24/X vssd1 vssd1 vccd1 vccd1 hold23/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2147_ _2150_/CLK _2147_/D vssd1 vssd1 vccd1 vccd1 _2147_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1029_ _1029_/A vssd1 vssd1 vccd1 vccd1 _1029_/Y sky130_fd_sc_hd__inv_2
X_2078_ _2210_/CLK _2078_/D vssd1 vssd1 vccd1 vccd1 _2078_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1457__D _1776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1380_ _1245_/A _1131_/C _1448_/B _1379_/X vssd1 vssd1 vccd1 vccd1 _1724_/B sky130_fd_sc_hd__a211o_1
XFILLER_0_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2001_ _2001_/A _2001_/B _2001_/C _2028_/B vssd1 vssd1 vccd1 vccd1 _2001_/X sky130_fd_sc_hd__and4_1
XANTENNA__1164__B2 _1808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1927__B1 _2003_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1716_ _1716_/A _1716_/B _1829_/C vssd1 vssd1 vccd1 vccd1 _1765_/B sky130_fd_sc_hd__or3_4
XFILLER_0_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1156__S _1994_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1647_ _1697_/C _1646_/X _1645_/X _1669_/A vssd1 vssd1 vccd1 vccd1 _1647_/X sky130_fd_sc_hd__o2bb2a_1
X_1578_ _1697_/A _1578_/B vssd1 vssd1 vccd1 vccd1 _1578_/Y sky130_fd_sc_hd__nor2_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1830__D _1920_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1855__A _1863_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1501_ _1550_/S vssd1 vssd1 vccd1 vccd1 _1501_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1704__S _1920_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1363_ hold87/X _1363_/B vssd1 vssd1 vccd1 vccd1 _1365_/C sky130_fd_sc_hd__xnor2_1
X_1432_ _1186_/Y _1228_/Y _1430_/X _1431_/X vssd1 vssd1 vccd1 vccd1 _1432_/X sky130_fd_sc_hd__a211o_1
X_1294_ _1297_/A _1980_/A vssd1 vssd1 vccd1 vccd1 _2001_/B sky130_fd_sc_hd__or2_1
XFILLER_0_73_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1612__A2 _1826_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1367__A1 _1776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1981_ _1297_/A _1960_/B _1984_/B _2015_/A vssd1 vssd1 vccd1 vccd1 _1981_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_7_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1415_ _1057_/A _1085_/A _1415_/A3 _1340_/X _1396_/B vssd1 vssd1 vccd1 vccd1 _1416_/D
+ sky130_fd_sc_hd__a311o_1
X_1346_ _1724_/A _1346_/B vssd1 vssd1 vccd1 vccd1 _1346_/X sky130_fd_sc_hd__or2_1
X_1277_ _1297_/A _1980_/A vssd1 vssd1 vccd1 vccd1 _1278_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_61_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1521__A1 _2112_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1200_ hold77/A _1499_/B _1198_/X _1882_/A vssd1 vssd1 vccd1 vccd1 _1202_/A sky130_fd_sc_hd__o211ai_2
X_2180_ _2219_/CLK hold62/X vssd1 vssd1 vccd1 vccd1 hold61/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1062_ _1143_/A _1344_/A vssd1 vssd1 vccd1 vccd1 _1062_/Y sky130_fd_sc_hd__nor2_1
X_1131_ _1245_/A _1245_/B _1131_/C vssd1 vssd1 vccd1 vccd1 _1135_/A sky130_fd_sc_hd__and3_4
X_1964_ _1964_/A _1964_/B vssd1 vssd1 vccd1 vccd1 _1964_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_55_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1895_ _1922_/B _1895_/B vssd1 vssd1 vccd1 vccd1 _1896_/S sky130_fd_sc_hd__nor2_1
XFILLER_0_28_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1329_ _1062_/Y _1415_/A3 _1340_/B _1119_/A _1410_/C vssd1 vssd1 vccd1 vccd1 _1333_/B
+ sky130_fd_sc_hd__a221o_1
XANTENNA__1863__A _1863_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold9 hold9/A vssd1 vssd1 vccd1 vccd1 hold9/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_57_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1680_ _1680_/A _1680_/B _1705_/B vssd1 vssd1 vccd1 vccd1 _1707_/B sky130_fd_sc_hd__or3_1
XFILLER_0_20_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1497__B1 _1994_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1712__S _1920_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2163_ _2209_/CLK _2163_/D vssd1 vssd1 vccd1 vccd1 _2163_/Q sky130_fd_sc_hd__dfxtp_2
X_1114_ _2080_/Q _1114_/B _1821_/B _2079_/Q vssd1 vssd1 vccd1 vccd1 _1138_/B sky130_fd_sc_hd__or4b_2
X_2094_ _2172_/CLK _2094_/D vssd1 vssd1 vccd1 vccd1 _2094_/Q sky130_fd_sc_hd__dfxtp_1
X_1045_ _2082_/Q _2081_/Q vssd1 vssd1 vccd1 vccd1 _1084_/A sky130_fd_sc_hd__nand2b_2
XFILLER_0_71_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1947_ _1947_/A _1973_/B vssd1 vssd1 vccd1 vccd1 _1948_/B sky130_fd_sc_hd__or2_1
X_1878_ _1877_/X _1864_/B _1907_/S vssd1 vssd1 vccd1 vccd1 _1878_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_43_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold217 _1156_/X vssd1 vssd1 vccd1 vccd1 _1870_/B sky130_fd_sc_hd__buf_1
XFILLER_0_53_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1663_ _1663_/A _1663_/B vssd1 vssd1 vccd1 vccd1 _1663_/Y sky130_fd_sc_hd__xnor2_1
Xhold206 _2141_/Q vssd1 vssd1 vccd1 vccd1 hold206/X sky130_fd_sc_hd__dlygate4sd3_1
X_1801_ _2114_/Q _1135_/A _1776_/X _2139_/Q _1717_/B vssd1 vssd1 vccd1 vccd1 _1804_/C
+ sky130_fd_sc_hd__a221oi_2
X_1732_ _1732_/A _1732_/B vssd1 vssd1 vccd1 vccd1 _1734_/D sky130_fd_sc_hd__nand2_1
XFILLER_0_25_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold228 _2155_/Q vssd1 vssd1 vccd1 vccd1 hold228/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1706__A1 _1921_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1594_ _2139_/Q _1776_/A _1868_/B _1469_/X vssd1 vssd1 vccd1 vccd1 _1594_/X sky130_fd_sc_hd__a22o_1
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold239 _2077_/Q vssd1 vssd1 vccd1 vccd1 _1111_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2215_ _2223_/CLK hold64/X vssd1 vssd1 vccd1 vccd1 hold63/A sky130_fd_sc_hd__dfxtp_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2077_ _2210_/CLK _2077_/D vssd1 vssd1 vccd1 vccd1 _2077_/Q sky130_fd_sc_hd__dfxtp_1
X_2146_ _2150_/CLK _2146_/D vssd1 vssd1 vccd1 vccd1 _2146_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1028_ _1028_/A vssd1 vssd1 vccd1 vccd1 _1028_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_36_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2000_ _2000_/A _2000_/B vssd1 vssd1 vccd1 vccd1 _2188_/D sky130_fd_sc_hd__and2_1
XFILLER_0_26_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1498__A _1918_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1927__A1 _1994_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1646_ _1476_/C _1652_/S _1475_/Y vssd1 vssd1 vccd1 vccd1 _1646_/X sky130_fd_sc_hd__a21o_1
X_1715_ _1716_/A _1829_/C vssd1 vssd1 vccd1 vccd1 _1808_/B sky130_fd_sc_hd__or2_4
XFILLER_0_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1577_ _1632_/A _1581_/S _1573_/X vssd1 vssd1 vccd1 vccd1 _1578_/B sky130_fd_sc_hd__a21oi_1
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2129_ _2209_/CLK _2129_/D vssd1 vssd1 vccd1 vccd1 _2129_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1871__A _1871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1500_ _2003_/A _1500_/B vssd1 vssd1 vccd1 vccd1 _1550_/S sky130_fd_sc_hd__or2_4
XFILLER_0_50_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1293_ _1297_/A _1980_/A vssd1 vssd1 vccd1 vccd1 _1360_/B sky130_fd_sc_hd__nor2_1
X_1362_ _2162_/Q _2160_/Q _2165_/Q _2161_/Q hold81/A hold73/A vssd1 vssd1 vccd1 vccd1
+ _1363_/B sky130_fd_sc_hd__mux4_1
X_1431_ _2129_/Q _1227_/B _1422_/Y _2112_/Q vssd1 vssd1 vccd1 vccd1 _1431_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_58_330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1629_ _2136_/Q _1776_/A _1784_/A _1469_/X vssd1 vssd1 vccd1 vccd1 _1629_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_41_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1980_ _1980_/A _1980_/B _2001_/C _1984_/C vssd1 vssd1 vccd1 vccd1 _1980_/X sky130_fd_sc_hd__and4_1
XFILLER_0_55_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1776__A _1776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1276_ _1279_/A vssd1 vssd1 vccd1 vccd1 _1276_/Y sky130_fd_sc_hd__inv_2
X_1414_ _1414_/A _1414_/B _1414_/C _1414_/D vssd1 vssd1 vccd1 vccd1 _1416_/C sky130_fd_sc_hd__or4_1
X_1345_ _1345_/A _1345_/B vssd1 vssd1 vccd1 vccd1 _1346_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_1_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _2142_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_69_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1130_ _1130_/A _1130_/B _1130_/C vssd1 vssd1 vccd1 vccd1 _1149_/B sky130_fd_sc_hd__or3_4
XFILLER_0_20_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1061_ _1344_/A _1141_/B vssd1 vssd1 vccd1 vccd1 _1061_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_28_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1963_ _1955_/B _1954_/B _1962_/X _1973_/A vssd1 vssd1 vccd1 vccd1 _1964_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_55_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1894_ _1141_/X _1893_/Y _1883_/X vssd1 vssd1 vccd1 vccd1 _1897_/S sky130_fd_sc_hd__a21bo_1
XFILLER_0_43_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1259_ _1784_/A hold3/X _2166_/Q vssd1 vssd1 vccd1 vccd1 _1260_/B sky130_fd_sc_hd__mux2_1
XANTENNA__1503__A2 _1517_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1328_ _1487_/B _1415_/A3 _1340_/B _1128_/A vssd1 vssd1 vccd1 vccd1 _1410_/C sky130_fd_sc_hd__a22o_1
XFILLER_0_34_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1975__C1 _2003_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1430__B2 _2163_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2093_ _2172_/CLK _2093_/D vssd1 vssd1 vccd1 vccd1 _2093_/Q sky130_fd_sc_hd__dfxtp_1
X_2162_ _2208_/CLK _2162_/D vssd1 vssd1 vccd1 vccd1 _2162_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__1497__A1 _1517_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1113_ _1377_/A _1121_/B vssd1 vssd1 vccd1 vccd1 _1723_/A sky130_fd_sc_hd__nor2_1
X_1044_ _2082_/Q _2081_/Q vssd1 vssd1 vccd1 vccd1 _1044_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_61_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1946_ _1946_/A _2008_/B vssd1 vssd1 vccd1 vccd1 _1973_/B sky130_fd_sc_hd__or2_1
X_1877_ _1876_/X _1239_/B _1877_/S vssd1 vssd1 vccd1 vccd1 _1877_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_43_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwrapped_6502_80 vssd1 vssd1 vccd1 vccd1 wrapped_6502_80/HI io_out[28] sky130_fd_sc_hd__conb_1
XFILLER_0_39_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2035__A _2057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1800_ _1800_/A _1806_/B vssd1 vssd1 vccd1 vccd1 _1804_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_25_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold229 _1796_/A vssd1 vssd1 vccd1 vccd1 _1867_/B sky130_fd_sc_hd__buf_1
X_1662_ _1662_/A _1662_/B vssd1 vssd1 vccd1 vccd1 _1662_/X sky130_fd_sc_hd__xor2_1
XANTENNA__1784__A _1784_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold207 _2139_/Q vssd1 vssd1 vccd1 vccd1 hold207/X sky130_fd_sc_hd__dlygate4sd3_1
X_1731_ _1034_/Y _1717_/B _1765_/B _2111_/Q vssd1 vssd1 vccd1 vccd1 _1734_/C sky130_fd_sc_hd__a22oi_2
Xhold218 _2137_/Q vssd1 vssd1 vccd1 vccd1 hold218/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2214_ _2214_/CLK hold72/X vssd1 vssd1 vccd1 vccd1 hold71/A sky130_fd_sc_hd__dfxtp_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1706__A2 hold194/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1593_ _1593_/A _1593_/B _1593_/C vssd1 vssd1 vccd1 vccd1 _1693_/A sky130_fd_sc_hd__and3_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2076_ _2223_/CLK hold86/X vssd1 vssd1 vccd1 vccd1 hold85/A sky130_fd_sc_hd__dfxtp_1
X_1027_ _1873_/B vssd1 vssd1 vccd1 vccd1 _1027_/Y sky130_fd_sc_hd__inv_2
X_2145_ _2164_/CLK _2145_/D vssd1 vssd1 vccd1 vccd1 _2145_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1929_ _2169_/Q _1933_/B vssd1 vssd1 vccd1 vccd1 _1929_/X sky130_fd_sc_hd__or2_1
XFILLER_0_48_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1869__A _1871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_14_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _2182_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold90 hold90/A vssd1 vssd1 vccd1 vccd1 hold90/X sky130_fd_sc_hd__dlygate4sd3_1
X_1645_ _1643_/A _1643_/B _1652_/S vssd1 vssd1 vccd1 vccd1 _1645_/X sky130_fd_sc_hd__o21a_1
X_1576_ _1476_/C _1573_/X _1581_/S _1575_/Y _1475_/Y vssd1 vssd1 vccd1 vccd1 _1576_/X
+ sky130_fd_sc_hd__a311o_1
X_1714_ _1104_/A _1044_/X _1097_/X _1245_/C vssd1 vssd1 vccd1 vccd1 _1829_/C sky130_fd_sc_hd__o22a_1
XFILLER_0_13_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2059_ hold35/X _1503_/X _2066_/S vssd1 vssd1 vccd1 vccd1 hold36/A sky130_fd_sc_hd__mux2_1
X_2128_ _2209_/CLK hold99/X vssd1 vssd1 vccd1 vccd1 hold98/A sky130_fd_sc_hd__dfxtp_1
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1871__B _1871_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1430_ _2121_/Q _1441_/B _1423_/X _2163_/Q vssd1 vssd1 vccd1 vccd1 _1430_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1292_ _1980_/A _2015_/B _1355_/C _1947_/A vssd1 vssd1 vccd1 vccd1 _1336_/B sky130_fd_sc_hd__or4_1
X_1361_ _1061_/Y _1373_/A2 _1285_/B _1360_/X vssd1 vssd1 vccd1 vccd1 _1407_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_58_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1559_ _1882_/A _1882_/B _1498_/B _2003_/A vssd1 vssd1 vccd1 vccd1 _1567_/S sky130_fd_sc_hd__a31o_4
X_1628_ _1628_/A _1628_/B vssd1 vssd1 vccd1 vccd1 _1662_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_1_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1866__B _1866_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold236_A _2160_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1524__B1 _1517_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_356 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1413_ _1413_/A _1413_/B _1413_/C _1413_/D vssd1 vssd1 vccd1 vccd1 _2081_/D sky130_fd_sc_hd__or4_1
XFILLER_0_64_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1275_ _1355_/B _2008_/A vssd1 vssd1 vccd1 vccd1 _1279_/A sky130_fd_sc_hd__or2_1
XANTENNA__1818__A1 _1871_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1344_ _1344_/A _1377_/B vssd1 vssd1 vccd1 vccd1 _1724_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_73_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1178__S _1994_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1906__S _1912_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1060_ _1821_/B _1114_/B _2079_/Q _2080_/Q vssd1 vssd1 vccd1 vccd1 _1141_/B sky130_fd_sc_hd__nand4b_4
XANTENNA_output35_A _1234_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1962_ _2015_/A _1980_/B _2015_/C _2015_/B vssd1 vssd1 vccd1 vccd1 _1962_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_28_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1893_ _2028_/A _1448_/B _1881_/X vssd1 vssd1 vccd1 vccd1 _1893_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_28_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_14_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1258_ _1728_/B _1258_/B vssd1 vssd1 vccd1 vccd1 _1306_/A sky130_fd_sc_hd__nand2_2
X_1189_ _2112_/Q _1149_/B _1186_/Y _1467_/A _1188_/X vssd1 vssd1 vccd1 vccd1 _1189_/X
+ sky130_fd_sc_hd__a221o_1
X_1327_ _1486_/A _1415_/A3 _1340_/B _1830_/B vssd1 vssd1 vccd1 vccd1 _1389_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_61_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2092_ _2172_/CLK _2092_/D vssd1 vssd1 vccd1 vccd1 _2092_/Q sky130_fd_sc_hd__dfxtp_1
X_2161_ _2209_/CLK _2161_/D vssd1 vssd1 vccd1 vccd1 _2161_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_45_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1043_ _1377_/A _1143_/A vssd1 vssd1 vccd1 vccd1 _1421_/A sky130_fd_sc_hd__nor2_2
X_1112_ _1345_/A _1335_/B vssd1 vssd1 vccd1 vccd1 _1238_/A sky130_fd_sc_hd__nor2_1
X_1945_ _1945_/A _1995_/B vssd1 vssd1 vccd1 vccd1 _2005_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_43_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1876_ _1027_/Y hold175/X _1912_/A vssd1 vssd1 vccd1 vccd1 _1876_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_43_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwrapped_6502_81 vssd1 vssd1 vccd1 vccd1 wrapped_6502_81/HI io_out[29] sky130_fd_sc_hd__conb_1
XFILLER_0_39_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1939__B1 _2003_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1661_ _1662_/A _1662_/B vssd1 vssd1 vccd1 vccd1 _1661_/X sky130_fd_sc_hd__and2_1
X_1592_ _1651_/A _1491_/B _1592_/S vssd1 vssd1 vccd1 vccd1 _1593_/C sky130_fd_sc_hd__mux2_1
Xhold208 _1840_/X vssd1 vssd1 vccd1 vccd1 _1841_/B sky130_fd_sc_hd__dlygate4sd3_1
X_1730_ _1728_/Y _1729_/X _1921_/B vssd1 vssd1 vccd1 vccd1 _1734_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_13_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold219 _1836_/X vssd1 vssd1 vccd1 vccd1 _1837_/B sky130_fd_sc_hd__dlygate4sd3_1
X_2213_ _2225_/CLK hold50/X vssd1 vssd1 vccd1 vccd1 hold49/A sky130_fd_sc_hd__dfxtp_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2144_ _2164_/CLK _2144_/D vssd1 vssd1 vccd1 vccd1 _2144_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2075_ hold17/X _1549_/X _2075_/S vssd1 vssd1 vccd1 vccd1 hold18/A sky130_fd_sc_hd__mux2_1
X_1026_ _1994_/A vssd1 vssd1 vccd1 vccd1 _1921_/A sky130_fd_sc_hd__inv_2
XFILLER_0_8_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1928_ hold3/X _1920_/Y _1927_/X vssd1 vssd1 vccd1 vccd1 hold4/A sky130_fd_sc_hd__a21o_1
XFILLER_0_44_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1859_ _1863_/A _1859_/B vssd1 vssd1 vccd1 vccd1 _2148_/D sky130_fd_sc_hd__and2_1
XANTENNA__1330__A1 _1517_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold91 hold91/A vssd1 vssd1 vccd1 vccd1 hold91/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold80 hold80/A vssd1 vssd1 vccd1 vccd1 hold80/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1927__A3 _1920_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1713_ hold91/X _1476_/B _1920_/A vssd1 vssd1 vccd1 vccd1 hold92/A sky130_fd_sc_hd__mux2_1
XFILLER_0_26_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1575_ _1573_/X _1581_/S _1669_/A vssd1 vssd1 vccd1 vccd1 _1575_/Y sky130_fd_sc_hd__a21oi_1
X_1644_ _2119_/Q _1826_/D _1460_/Y _1864_/B vssd1 vssd1 vccd1 vccd1 _1652_/S sky130_fd_sc_hd__a22o_1
XFILLER_0_6_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2127_ _2209_/CLK _2127_/D vssd1 vssd1 vccd1 vccd1 _2127_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2058_ _1882_/A _1499_/B _1542_/A _2003_/A vssd1 vssd1 vccd1 vccd1 _2066_/S sky130_fd_sc_hd__a31o_4
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1360_ _1984_/B _1360_/B _1360_/C vssd1 vssd1 vccd1 vccd1 _1360_/X sky130_fd_sc_hd__and3_1
XFILLER_0_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1291_ _2015_/A _1996_/A _1285_/B _1336_/A vssd1 vssd1 vccd1 vccd1 _1299_/A sky130_fd_sc_hd__a211o_1
XFILLER_0_37_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1558_ _2049_/A _1558_/B vssd1 vssd1 vccd1 vccd1 _2098_/D sky130_fd_sc_hd__and2_1
X_1627_ _1626_/B _1626_/C _1626_/A vssd1 vssd1 vccd1 vccd1 _1628_/B sky130_fd_sc_hd__a21oi_1
X_1489_ _1697_/A _1654_/B _1479_/X vssd1 vssd1 vccd1 vccd1 _1570_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__1781__A1 _2053_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold229_A _1796_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1412_ _1412_/A _1412_/B _1412_/C vssd1 vssd1 vccd1 vccd1 _1413_/D sky130_fd_sc_hd__or3_1
X_1343_ _1129_/B _1365_/A _1403_/A2 _1238_/A _1416_/B vssd1 vssd1 vccd1 vccd1 _1411_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_11_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1274_ _1945_/A _1995_/B vssd1 vssd1 vccd1 vccd1 _2008_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_3_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1194__S _1994_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1832__S _1862_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1961_ _1973_/A _1973_/B _2036_/B _1336_/B _1336_/A vssd1 vssd1 vccd1 vccd1 _1964_/A
+ sky130_fd_sc_hd__o32a_1
X_1892_ hold147/X _1884_/Y _1891_/Y vssd1 vssd1 vccd1 vccd1 _1892_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_28_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_168 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1326_ _1717_/B _1365_/A _1403_/A2 _1903_/B _1416_/A vssd1 vssd1 vccd1 vccd1 _1405_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_11_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1257_ _1728_/B _1258_/B vssd1 vssd1 vccd1 vccd1 _1281_/B sky130_fd_sc_hd__and2_1
X_1188_ hold190/X _1149_/C _1827_/B _1866_/B vssd1 vssd1 vccd1 vccd1 _1188_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_338 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1888__A _2112_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2160_ _2210_/CLK _2160_/D vssd1 vssd1 vccd1 vccd1 _2160_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_0_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2091_ _2172_/CLK _2091_/D vssd1 vssd1 vccd1 vccd1 hold94/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1042_ _1821_/A _1236_/D _1821_/B _1114_/B vssd1 vssd1 vccd1 vccd1 _1143_/A sky130_fd_sc_hd__or4b_2
X_1111_ _1111_/A _1826_/A vssd1 vssd1 vccd1 vccd1 _1335_/B sky130_fd_sc_hd__nand2_1
X_1944_ _2001_/A _1995_/B vssd1 vssd1 vccd1 vccd1 _1973_/A sky130_fd_sc_hd__or2_1
X_1875_ _1873_/X _1877_/S _1872_/X vssd1 vssd1 vccd1 vccd1 _1879_/S sky130_fd_sc_hd__o21a_1
XFILLER_0_0_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1709__B2 _1921_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwrapped_6502_82 vssd1 vssd1 vccd1 vccd1 wrapped_6502_82/HI io_out[30] sky130_fd_sc_hd__conb_1
X_1309_ _2015_/B _2001_/B vssd1 vssd1 vccd1 vccd1 _1313_/B sky130_fd_sc_hd__or2_1
XFILLER_0_47_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1939__A1 _1994_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1660_ _1663_/A _1659_/B _1639_/X vssd1 vssd1 vccd1 vccd1 _1662_/B sky130_fd_sc_hd__a21o_1
X_1591_ _1491_/B _1593_/A _1491_/A vssd1 vssd1 vccd1 vccd1 _1593_/B sky130_fd_sc_hd__a21o_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold209 _2138_/Q vssd1 vssd1 vccd1 vccd1 hold209/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2212_ _2226_/CLK hold14/X vssd1 vssd1 vccd1 vccd1 hold13/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2143_ _2164_/CLK _2143_/D vssd1 vssd1 vccd1 vccd1 _2143_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2074_ hold47/X _1542_/X _2075_/S vssd1 vssd1 vccd1 vccd1 hold48/A sky130_fd_sc_hd__mux2_1
XFILLER_0_48_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1025_ _2210_/Q vssd1 vssd1 vccd1 vccd1 _1025_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_29_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1927_ _1994_/A _2092_/Q _1920_/B _2003_/A vssd1 vssd1 vccd1 vccd1 _1927_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_44_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1858_ hold183/X _1166_/X _1862_/S vssd1 vssd1 vccd1 vccd1 _1859_/B sky130_fd_sc_hd__mux2_1
X_1789_ _2112_/Q _1135_/A _1776_/X _2137_/Q _1717_/B vssd1 vssd1 vccd1 vccd1 _1792_/C
+ sky130_fd_sc_hd__a221oi_2
XFILLER_0_12_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold70 hold70/A vssd1 vssd1 vccd1 vccd1 hold70/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold92 hold92/A vssd1 vssd1 vccd1 vccd1 hold92/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold81 hold81/A vssd1 vssd1 vccd1 vccd1 hold81/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1840__S _1862_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1609__B1 _1866_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1712_ _1545_/B _1690_/X _1920_/A vssd1 vssd1 vccd1 vccd1 _2117_/D sky130_fd_sc_hd__mux2_1
X_1643_ _1643_/A _1643_/B vssd1 vssd1 vccd1 vccd1 _1697_/C sky130_fd_sc_hd__or2_1
XANTENNA_1 hold175/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1574_ _2125_/Q _1826_/D _1460_/Y _1156_/X vssd1 vssd1 vccd1 vccd1 _1581_/S sky130_fd_sc_hd__a22o_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2057_ _2057_/A _2057_/B vssd1 vssd1 vccd1 vccd1 _2210_/D sky130_fd_sc_hd__and2_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2126_ _2142_/CLK _2126_/D vssd1 vssd1 vccd1 vccd1 _2126_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout77_A _1918_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2057__A _2057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1290_ _1306_/A _1306_/B vssd1 vssd1 vccd1 vccd1 _1996_/A sky130_fd_sc_hd__or2_2
XFILLER_0_37_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1626_ _1626_/A _1626_/B _1626_/C vssd1 vssd1 vccd1 vccd1 _1628_/A sky130_fd_sc_hd__and3_1
XFILLER_0_5_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1557_ _2049_/A input9/X vssd1 vssd1 vccd1 vccd1 _2097_/D sky130_fd_sc_hd__and2_1
X_1488_ _1488_/A _1488_/B _1488_/C vssd1 vssd1 vccd1 vccd1 _1654_/B sky130_fd_sc_hd__or3_1
XTAP_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2109_ _2223_/CLK hold90/X vssd1 vssd1 vccd1 vccd1 hold89/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1273_ _1945_/A _1995_/B vssd1 vssd1 vccd1 vccd1 _1273_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_48_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1342_ _1075_/C _1365_/A _1340_/B _1229_/B vssd1 vssd1 vccd1 vccd1 _1416_/B sky130_fd_sc_hd__a22o_1
X_1411_ _1411_/A _1411_/B _1411_/C _1411_/D vssd1 vssd1 vccd1 vccd1 _1412_/C sky130_fd_sc_hd__or4_1
XFILLER_0_3_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1987__C1 _2057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1609_ _2137_/Q _1776_/A _1866_/B _1469_/X vssd1 vssd1 vccd1 vccd1 _1609_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_1_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1442__B2 _2165_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1960_ _2015_/C _1960_/B vssd1 vssd1 vccd1 vccd1 _2036_/B sky130_fd_sc_hd__nand2_1
X_1891_ _1884_/Y _1890_/X _1918_/A vssd1 vssd1 vccd1 vccd1 _1891_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1256_ _1864_/B _2167_/Q _2166_/Q vssd1 vssd1 vccd1 vccd1 _1258_/B sky130_fd_sc_hd__mux2_1
X_1325_ _1051_/Y _1365_/A _1403_/A2 _1486_/B vssd1 vssd1 vccd1 vccd1 _1416_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_59_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1187_ hold221/X hold102/X _1994_/A vssd1 vssd1 vccd1 vccd1 _1866_/B sky130_fd_sc_hd__mux2_4
XFILLER_0_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1994__A _1994_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1424__B2 _2160_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold191_A _2108_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2090_ _2226_/CLK hold22/X vssd1 vssd1 vccd1 vccd1 hold21/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1110_ _1829_/A _1455_/B _1486_/D _1110_/D vssd1 vssd1 vccd1 vccd1 _1130_/A sky130_fd_sc_hd__or4_1
Xclkbuf_4_0_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _2150_/CLK sky130_fd_sc_hd__clkbuf_8
X_1041_ _2081_/Q _2082_/Q vssd1 vssd1 vccd1 vccd1 _1041_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_0_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1943_ _2001_/A _1995_/B vssd1 vssd1 vccd1 vccd1 _1984_/C sky130_fd_sc_hd__nor2_2
X_1874_ _2006_/A _1874_/B _1997_/A vssd1 vssd1 vccd1 vccd1 _1877_/S sky130_fd_sc_hd__or3_1
XFILLER_0_43_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapped_6502_83 vssd1 vssd1 vccd1 vccd1 wrapped_6502_83/HI io_out[34] sky130_fd_sc_hd__conb_1
X_1308_ _1278_/B _1960_/B _1307_/Y _1304_/X _1287_/B vssd1 vssd1 vccd1 vccd1 _1393_/B
+ sky130_fd_sc_hd__o32a_1
X_1239_ _1239_/A _1239_/B vssd1 vssd1 vccd1 vccd1 _1241_/A sky130_fd_sc_hd__or2_1
XFILLER_0_62_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1838__S _1862_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1590_ _1697_/A _1573_/X _1589_/X vssd1 vssd1 vccd1 vccd1 _1593_/A sky130_fd_sc_hd__a21o_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1572__B1 _1156_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2073_ hold25/X _1535_/X _2075_/S vssd1 vssd1 vccd1 vccd1 hold26/A sky130_fd_sc_hd__mux2_1
X_2211_ _2214_/CLK hold36/X vssd1 vssd1 vccd1 vccd1 hold35/A sky130_fd_sc_hd__dfxtp_1
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2142_ _2142_/CLK _2142_/D vssd1 vssd1 vccd1 vccd1 _2142_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1926_ hold94/X _1920_/Y _1925_/X _1871_/A vssd1 vssd1 vccd1 vccd1 hold95/A sky130_fd_sc_hd__o211a_1
XFILLER_0_44_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1788_ _1788_/A _1806_/B vssd1 vssd1 vccd1 vccd1 _1792_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_24_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1857_ _1863_/A _1857_/B vssd1 vssd1 vccd1 vccd1 _2147_/D sky130_fd_sc_hd__and2_1
XFILLER_0_47_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold71 hold71/A vssd1 vssd1 vccd1 vccd1 hold71/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold60 hold60/A vssd1 vssd1 vccd1 vccd1 hold60/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 hold82/A vssd1 vssd1 vccd1 vccd1 hold82/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold93 hold93/A vssd1 vssd1 vccd1 vccd1 hold93/X sky130_fd_sc_hd__buf_1
XANTENNA__1568__S _1994_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1711_ hold193/X _1694_/Y _1920_/A vssd1 vssd1 vccd1 vccd1 _2116_/D sky130_fd_sc_hd__mux2_1
X_1642_ _2110_/Q _1460_/A _1641_/X vssd1 vssd1 vccd1 vccd1 _1643_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_26_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1573_ _2116_/Q _1460_/A _1468_/A _1155_/Y _1572_/X vssd1 vssd1 vccd1 vccd1 _1573_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2056_ _1025_/Y _1903_/B hold164/X vssd1 vssd1 vccd1 vccd1 _2056_/Y sky130_fd_sc_hd__o21ai_1
X_2125_ _2150_/CLK _2125_/D vssd1 vssd1 vccd1 vccd1 _2125_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1909_ _2057_/A _1909_/B vssd1 vssd1 vccd1 vccd1 _2164_/D sky130_fd_sc_hd__and2_1
XFILLER_0_8_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1556_ _2049_/A input8/X vssd1 vssd1 vccd1 vccd1 _2096_/D sky130_fd_sc_hd__and2_1
X_1625_ _1651_/A _1491_/B _1625_/S vssd1 vssd1 vccd1 vccd1 _1626_/C sky130_fd_sc_hd__mux2_1
XFILLER_0_5_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1487_ _1487_/A _1487_/B _1487_/C _1054_/C vssd1 vssd1 vccd1 vccd1 _1488_/C sky130_fd_sc_hd__or4b_1
XTAP_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2108_ _2223_/CLK _2108_/D vssd1 vssd1 vccd1 vccd1 _2108_/Q sky130_fd_sc_hd__dfxtp_2
X_2039_ hold188/X _2043_/B _1990_/Y _2031_/B vssd1 vssd1 vccd1 vccd1 _2039_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_49_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_4_13_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _2214_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_32_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1846__S _1862_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1410_ _1410_/A _1410_/B _1410_/C _1410_/D vssd1 vssd1 vccd1 vccd1 _1411_/D sky130_fd_sc_hd__or4_1
XFILLER_0_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1212__A2 _1808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1272_ _1728_/B _1272_/B vssd1 vssd1 vccd1 vccd1 _1995_/B sky130_fd_sc_hd__and2_4
XFILLER_0_48_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1341_ _1085_/A _1415_/A3 _1340_/B _1459_/B _1340_/X vssd1 vssd1 vccd1 vccd1 _1406_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_3_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1451__A2 _1776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1608_ _1186_/A _1186_/B _1468_/Y vssd1 vssd1 vccd1 vccd1 _1611_/A sky130_fd_sc_hd__a21o_1
X_1539_ _1539_/A _1539_/B vssd1 vssd1 vccd1 vccd1 _1540_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold234_A _2162_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold190 _2145_/Q vssd1 vssd1 vccd1 vccd1 hold190/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1969__B1 _2003_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1890_ _1887_/X _1888_/X _1889_/X _1886_/Y _1895_/B vssd1 vssd1 vccd1 vccd1 _1890_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_0_11_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1186_ _1186_/A _1186_/B vssd1 vssd1 vccd1 vccd1 _1186_/Y sky130_fd_sc_hd__nand2_1
X_1255_ _1946_/A vssd1 vssd1 vccd1 vccd1 _1255_/Y sky130_fd_sc_hd__inv_2
X_1324_ _1033_/A _1229_/X _1296_/B _1373_/A2 _1469_/A vssd1 vssd1 vccd1 vccd1 _1417_/A
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_34_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1188__B2 _1866_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout52_A _1284_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1179__B2 _1796_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1040_ _2081_/Q _1040_/B vssd1 vssd1 vccd1 vccd1 _1104_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_68_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1942_ hold93/X _1921_/B _2003_/A vssd1 vssd1 vccd1 vccd1 _2176_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_28_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1873_ _1912_/A _1873_/B _1873_/C _2080_/Q vssd1 vssd1 vccd1 vccd1 _1873_/X sky130_fd_sc_hd__or4b_1
XFILLER_0_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapped_6502_84 vssd1 vssd1 vccd1 vccd1 wrapped_6502_84/HI io_out[35] sky130_fd_sc_hd__conb_1
XANTENNA__1054__B _1548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1169_ _1167_/X _1168_/X _1499_/A vssd1 vssd1 vccd1 vccd1 _1169_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1893__A2 _1448_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1307_ _1984_/B _2001_/C vssd1 vssd1 vccd1 vccd1 _1307_/Y sky130_fd_sc_hd__nor2_1
X_1238_ _1238_/A _1238_/B _1895_/B _1238_/D vssd1 vssd1 vccd1 vccd1 _1238_/X sky130_fd_sc_hd__or4_1
XFILLER_0_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1939__A3 _1920_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1854__S _1862_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2210_ _2210_/CLK _2210_/D vssd1 vssd1 vccd1 vccd1 _2210_/Q sky130_fd_sc_hd__dfxtp_1
X_2072_ hold11/X _1528_/X _2075_/S vssd1 vssd1 vccd1 vccd1 hold12/A sky130_fd_sc_hd__mux2_1
X_2141_ _2142_/CLK _2141_/D vssd1 vssd1 vccd1 vccd1 _2141_/Q sky130_fd_sc_hd__dfxtp_1
X_1925_ _2167_/Q _1933_/B vssd1 vssd1 vccd1 vccd1 _1925_/X sky130_fd_sc_hd__or2_1
XFILLER_0_56_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1787_ _2053_/B2 _1785_/Y _1792_/A _1820_/A2 hold98/X vssd1 vssd1 vccd1 vccd1 hold99/A
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_12_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1856_ hold182/X _1173_/X _1862_/S vssd1 vssd1 vccd1 vccd1 _1857_/B sky130_fd_sc_hd__mux2_1
XANTENNA_hold147_A _2161_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1251__A0 _1866_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold94 hold94/A vssd1 vssd1 vccd1 vccd1 hold94/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 hold72/A vssd1 vssd1 vccd1 vccd1 hold72/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold50 hold50/A vssd1 vssd1 vccd1 vccd1 hold50/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold61 hold61/A vssd1 vssd1 vccd1 vccd1 hold61/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 hold83/A vssd1 vssd1 vccd1 vccd1 hold83/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1609__A2 _1776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1710_ hold180/X _1692_/Y _1920_/A vssd1 vssd1 vccd1 vccd1 _1710_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_53_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1572_ _2141_/Q _1776_/A _1156_/X _1469_/X vssd1 vssd1 vccd1 vccd1 _1572_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_41_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1641_ _2135_/Q _1776_/A _1864_/B _1469_/X vssd1 vssd1 vccd1 vccd1 _1641_/X sky130_fd_sc_hd__a22o_1
XANTENNA__1793__A1 _2053_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2124_ _2150_/CLK _2124_/D vssd1 vssd1 vccd1 vccd1 _2124_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1481__B1 _2160_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2055_ _2210_/Q _2055_/B _1941_/B vssd1 vssd1 vccd1 vccd1 _2055_/X sky130_fd_sc_hd__or3b_1
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1908_ hold214/X _1907_/X _1908_/S vssd1 vssd1 vccd1 vccd1 _1909_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_44_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1839_ _1863_/A _1839_/B vssd1 vssd1 vccd1 vccd1 _2138_/D sky130_fd_sc_hd__and2_1
XFILLER_0_8_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput40 _1206_/X vssd1 vssd1 vccd1 vccd1 io_out[3] sky130_fd_sc_hd__buf_12
XFILLER_0_41_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1555_ _2049_/A input7/X vssd1 vssd1 vccd1 vccd1 _2095_/D sky130_fd_sc_hd__and2_1
XANTENNA__1518__A1 _1517_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1624_ _1491_/B _1626_/A _1491_/A vssd1 vssd1 vccd1 vccd1 _1626_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_41_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2107_ _2214_/CLK _2107_/D vssd1 vssd1 vccd1 vccd1 _2107_/Q sky130_fd_sc_hd__dfxtp_2
X_1486_ _1486_/A _1486_/B _1907_/S _1486_/D vssd1 vssd1 vccd1 vccd1 _1487_/C sky130_fd_sc_hd__or4_1
XTAP_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2038_ _1029_/A _2028_/B _2037_/X _2057_/A vssd1 vssd1 vccd1 vccd1 _2200_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_43_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1253__A _1728_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1340_ _1723_/A _1340_/B vssd1 vssd1 vccd1 vccd1 _1340_/X sky130_fd_sc_hd__and2_1
XANTENNA__1862__S _1862_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1271_ _1156_/X hold53/X _2166_/Q vssd1 vssd1 vccd1 vccd1 _1272_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_3_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1538_ _2116_/Q _1538_/B vssd1 vssd1 vccd1 vccd1 _1539_/B sky130_fd_sc_hd__or2_1
X_1607_ _1691_/A _1607_/B vssd1 vssd1 vccd1 vccd1 _1707_/A sky130_fd_sc_hd__nor2_1
X_1469_ _1469_/A _1826_/D vssd1 vssd1 vccd1 vccd1 _1469_/X sky130_fd_sc_hd__or2_4
XFILLER_0_38_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold180 _2115_/Q vssd1 vssd1 vccd1 vccd1 hold180/X sky130_fd_sc_hd__buf_1
XFILLER_0_45_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_1_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold191 _2108_/Q vssd1 vssd1 vccd1 vccd1 _1239_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__1902__A1 _1866_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1323_ _1407_/A _1410_/B _1414_/B vssd1 vssd1 vccd1 vccd1 _1391_/A sky130_fd_sc_hd__or3_1
XFILLER_0_11_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1185_ hold39/A _1499_/B _1183_/X _1499_/A vssd1 vssd1 vccd1 vccd1 _1186_/B sky130_fd_sc_hd__o211ai_1
X_1254_ _1297_/A _2015_/A vssd1 vssd1 vccd1 vccd1 _1946_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_46_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1896__A0 _1545_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1888__D _2117_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1872_ _1033_/Y _1881_/A _1895_/B _1874_/B _1907_/S vssd1 vssd1 vccd1 vccd1 _1872_/X
+ sky130_fd_sc_hd__a221o_1
X_1941_ _2057_/A _1941_/B vssd1 vssd1 vccd1 vccd1 _2175_/D sky130_fd_sc_hd__and2_1
XFILLER_0_9_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1306_ _1306_/A _1306_/B vssd1 vssd1 vccd1 vccd1 _2008_/B sky130_fd_sc_hd__nand2_1
X_1168_ hold11/A hold51/A _1499_/B vssd1 vssd1 vccd1 vccd1 _1168_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_59_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1099_ _1344_/A _1121_/B vssd1 vssd1 vccd1 vccd1 _1459_/B sky130_fd_sc_hd__nor2_1
X_1237_ _1104_/A _1044_/X _1245_/C vssd1 vssd1 vccd1 vccd1 _1238_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_19_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1572__A2 _1776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2140_ _2142_/CLK _2140_/D vssd1 vssd1 vccd1 vccd1 _2140_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2071_ hold33/X _1525_/X _2075_/S vssd1 vssd1 vccd1 vccd1 hold34/A sky130_fd_sc_hd__mux2_1
X_1924_ _1920_/Y _1923_/Y _2003_/A vssd1 vssd1 vccd1 vccd1 _2166_/D sky130_fd_sc_hd__a21oi_1
X_1855_ _1863_/A _1855_/B vssd1 vssd1 vccd1 vccd1 _2146_/D sky130_fd_sc_hd__and2_1
X_1786_ _1785_/B _1785_/C _1785_/D _1785_/A vssd1 vssd1 vccd1 vccd1 _1792_/A sky130_fd_sc_hd__a31o_1
XFILLER_0_12_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold40 hold40/A vssd1 vssd1 vccd1 vccd1 hold40/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold95 hold95/A vssd1 vssd1 vccd1 vccd1 hold95/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 hold51/A vssd1 vssd1 vccd1 vccd1 hold51/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 hold62/A vssd1 vssd1 vccd1 vccd1 hold62/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 hold73/A vssd1 vssd1 vccd1 vccd1 hold73/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 hold84/A vssd1 vssd1 vccd1 vccd1 hold84/X sky130_fd_sc_hd__dlygate4sd3_1
X_1640_ _1202_/A _1202_/B _1468_/Y vssd1 vssd1 vccd1 vccd1 _1643_/A sky130_fd_sc_hd__a21oi_1
X_1571_ _1697_/B _1571_/B vssd1 vssd1 vccd1 vccd1 _1689_/A sky130_fd_sc_hd__and2_1
XFILLER_0_41_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2123_ _2150_/CLK _2123_/D vssd1 vssd1 vccd1 vccd1 _2123_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2054_ hold81/X _2054_/A2 _1355_/C _1735_/A vssd1 vssd1 vccd1 vccd1 hold82/A sky130_fd_sc_hd__a22o_1
XFILLER_0_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1907_ _1906_/X _1867_/B _1907_/S vssd1 vssd1 vccd1 vccd1 _1907_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_32_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1838_ hold209/X _1217_/X _1862_/S vssd1 vssd1 vccd1 vccd1 _1838_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1769__C1 _1717_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_6_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1769_ _2117_/Q _1765_/B _1776_/B _2150_/Q _1717_/B vssd1 vssd1 vccd1 vccd1 _1769_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_12_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput30 _1435_/X vssd1 vssd1 vccd1 vccd1 io_out[22] sky130_fd_sc_hd__buf_12
XFILLER_0_31_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput41 _1197_/X vssd1 vssd1 vccd1 vccd1 io_out[4] sky130_fd_sc_hd__buf_12
XFILLER_0_23_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1554_ _2049_/A input6/X vssd1 vssd1 vccd1 vccd1 _2094_/D sky130_fd_sc_hd__and2_1
X_1485_ _1448_/B _1481_/X _1483_/X _1459_/C vssd1 vssd1 vccd1 vccd1 _1488_/B sky130_fd_sc_hd__a22o_1
X_1623_ _1616_/X _1618_/X _1622_/Y _1697_/A vssd1 vssd1 vccd1 vccd1 _1626_/A sky130_fd_sc_hd__a22o_1
XTAP_166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
.ends

