VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO vliw
  CLASS BLOCK ;
  FOREIGN vliw ;
  ORIGIN 0.000 0.000 ;
  SIZE 2200.000 BY 800.000 ;
  PIN cache_PC[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.721000 ;
    PORT
      LAYER met2 ;
        RECT 41.950 796.000 42.230 800.000 ;
    END
  END cache_PC[0]
  PIN cache_PC[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 92.550 796.000 92.830 800.000 ;
    END
  END cache_PC[10]
  PIN cache_PC[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 97.610 796.000 97.890 800.000 ;
    END
  END cache_PC[11]
  PIN cache_PC[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 102.670 796.000 102.950 800.000 ;
    END
  END cache_PC[12]
  PIN cache_PC[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 107.730 796.000 108.010 800.000 ;
    END
  END cache_PC[13]
  PIN cache_PC[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 112.790 796.000 113.070 800.000 ;
    END
  END cache_PC[14]
  PIN cache_PC[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 117.850 796.000 118.130 800.000 ;
    END
  END cache_PC[15]
  PIN cache_PC[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 122.910 796.000 123.190 800.000 ;
    END
  END cache_PC[16]
  PIN cache_PC[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 127.970 796.000 128.250 800.000 ;
    END
  END cache_PC[17]
  PIN cache_PC[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 133.030 796.000 133.310 800.000 ;
    END
  END cache_PC[18]
  PIN cache_PC[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 138.090 796.000 138.370 800.000 ;
    END
  END cache_PC[19]
  PIN cache_PC[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 47.010 796.000 47.290 800.000 ;
    END
  END cache_PC[1]
  PIN cache_PC[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 143.150 796.000 143.430 800.000 ;
    END
  END cache_PC[20]
  PIN cache_PC[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 148.210 796.000 148.490 800.000 ;
    END
  END cache_PC[21]
  PIN cache_PC[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 153.270 796.000 153.550 800.000 ;
    END
  END cache_PC[22]
  PIN cache_PC[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 158.330 796.000 158.610 800.000 ;
    END
  END cache_PC[23]
  PIN cache_PC[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 163.390 796.000 163.670 800.000 ;
    END
  END cache_PC[24]
  PIN cache_PC[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 168.450 796.000 168.730 800.000 ;
    END
  END cache_PC[25]
  PIN cache_PC[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 173.510 796.000 173.790 800.000 ;
    END
  END cache_PC[26]
  PIN cache_PC[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 178.570 796.000 178.850 800.000 ;
    END
  END cache_PC[27]
  PIN cache_PC[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 52.070 796.000 52.350 800.000 ;
    END
  END cache_PC[2]
  PIN cache_PC[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 57.130 796.000 57.410 800.000 ;
    END
  END cache_PC[3]
  PIN cache_PC[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 62.190 796.000 62.470 800.000 ;
    END
  END cache_PC[4]
  PIN cache_PC[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 67.250 796.000 67.530 800.000 ;
    END
  END cache_PC[5]
  PIN cache_PC[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 72.310 796.000 72.590 800.000 ;
    END
  END cache_PC[6]
  PIN cache_PC[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 77.370 796.000 77.650 800.000 ;
    END
  END cache_PC[7]
  PIN cache_PC[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 82.430 796.000 82.710 800.000 ;
    END
  END cache_PC[8]
  PIN cache_PC[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 87.490 796.000 87.770 800.000 ;
    END
  END cache_PC[9]
  PIN cache_entry[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 183.630 796.000 183.910 800.000 ;
    END
  END cache_entry[0]
  PIN cache_entry[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 689.630 796.000 689.910 800.000 ;
    END
  END cache_entry[100]
  PIN cache_entry[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 694.690 796.000 694.970 800.000 ;
    END
  END cache_entry[101]
  PIN cache_entry[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 699.750 796.000 700.030 800.000 ;
    END
  END cache_entry[102]
  PIN cache_entry[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 704.810 796.000 705.090 800.000 ;
    END
  END cache_entry[103]
  PIN cache_entry[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met2 ;
        RECT 709.870 796.000 710.150 800.000 ;
    END
  END cache_entry[104]
  PIN cache_entry[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 714.930 796.000 715.210 800.000 ;
    END
  END cache_entry[105]
  PIN cache_entry[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 719.990 796.000 720.270 800.000 ;
    END
  END cache_entry[106]
  PIN cache_entry[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 725.050 796.000 725.330 800.000 ;
    END
  END cache_entry[107]
  PIN cache_entry[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 730.110 796.000 730.390 800.000 ;
    END
  END cache_entry[108]
  PIN cache_entry[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 735.170 796.000 735.450 800.000 ;
    END
  END cache_entry[109]
  PIN cache_entry[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 234.230 796.000 234.510 800.000 ;
    END
  END cache_entry[10]
  PIN cache_entry[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 740.230 796.000 740.510 800.000 ;
    END
  END cache_entry[110]
  PIN cache_entry[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 745.290 796.000 745.570 800.000 ;
    END
  END cache_entry[111]
  PIN cache_entry[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 750.350 796.000 750.630 800.000 ;
    END
  END cache_entry[112]
  PIN cache_entry[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 755.410 796.000 755.690 800.000 ;
    END
  END cache_entry[113]
  PIN cache_entry[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 760.470 796.000 760.750 800.000 ;
    END
  END cache_entry[114]
  PIN cache_entry[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met2 ;
        RECT 765.530 796.000 765.810 800.000 ;
    END
  END cache_entry[115]
  PIN cache_entry[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met2 ;
        RECT 770.590 796.000 770.870 800.000 ;
    END
  END cache_entry[116]
  PIN cache_entry[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 775.650 796.000 775.930 800.000 ;
    END
  END cache_entry[117]
  PIN cache_entry[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 780.710 796.000 780.990 800.000 ;
    END
  END cache_entry[118]
  PIN cache_entry[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 785.770 796.000 786.050 800.000 ;
    END
  END cache_entry[119]
  PIN cache_entry[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 239.290 796.000 239.570 800.000 ;
    END
  END cache_entry[11]
  PIN cache_entry[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 790.830 796.000 791.110 800.000 ;
    END
  END cache_entry[120]
  PIN cache_entry[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 795.890 796.000 796.170 800.000 ;
    END
  END cache_entry[121]
  PIN cache_entry[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met2 ;
        RECT 800.950 796.000 801.230 800.000 ;
    END
  END cache_entry[122]
  PIN cache_entry[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met2 ;
        RECT 806.010 796.000 806.290 800.000 ;
    END
  END cache_entry[123]
  PIN cache_entry[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 811.070 796.000 811.350 800.000 ;
    END
  END cache_entry[124]
  PIN cache_entry[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 816.130 796.000 816.410 800.000 ;
    END
  END cache_entry[125]
  PIN cache_entry[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.120500 ;
    ANTENNADIFFAREA 2.173500 ;
    PORT
      LAYER met2 ;
        RECT 821.190 796.000 821.470 800.000 ;
    END
  END cache_entry[126]
  PIN cache_entry[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.747000 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met2 ;
        RECT 826.250 796.000 826.530 800.000 ;
    END
  END cache_entry[127]
  PIN cache_entry[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 244.350 796.000 244.630 800.000 ;
    END
  END cache_entry[12]
  PIN cache_entry[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 249.410 796.000 249.690 800.000 ;
    END
  END cache_entry[13]
  PIN cache_entry[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 254.470 796.000 254.750 800.000 ;
    END
  END cache_entry[14]
  PIN cache_entry[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 259.530 796.000 259.810 800.000 ;
    END
  END cache_entry[15]
  PIN cache_entry[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 264.590 796.000 264.870 800.000 ;
    END
  END cache_entry[16]
  PIN cache_entry[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 269.650 796.000 269.930 800.000 ;
    END
  END cache_entry[17]
  PIN cache_entry[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 274.710 796.000 274.990 800.000 ;
    END
  END cache_entry[18]
  PIN cache_entry[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 279.770 796.000 280.050 800.000 ;
    END
  END cache_entry[19]
  PIN cache_entry[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 188.690 796.000 188.970 800.000 ;
    END
  END cache_entry[1]
  PIN cache_entry[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 284.830 796.000 285.110 800.000 ;
    END
  END cache_entry[20]
  PIN cache_entry[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 289.890 796.000 290.170 800.000 ;
    END
  END cache_entry[21]
  PIN cache_entry[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 294.950 796.000 295.230 800.000 ;
    END
  END cache_entry[22]
  PIN cache_entry[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 300.010 796.000 300.290 800.000 ;
    END
  END cache_entry[23]
  PIN cache_entry[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 305.070 796.000 305.350 800.000 ;
    END
  END cache_entry[24]
  PIN cache_entry[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 310.130 796.000 310.410 800.000 ;
    END
  END cache_entry[25]
  PIN cache_entry[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 315.190 796.000 315.470 800.000 ;
    END
  END cache_entry[26]
  PIN cache_entry[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 320.250 796.000 320.530 800.000 ;
    END
  END cache_entry[27]
  PIN cache_entry[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 325.310 796.000 325.590 800.000 ;
    END
  END cache_entry[28]
  PIN cache_entry[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 330.370 796.000 330.650 800.000 ;
    END
  END cache_entry[29]
  PIN cache_entry[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 193.750 796.000 194.030 800.000 ;
    END
  END cache_entry[2]
  PIN cache_entry[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 335.430 796.000 335.710 800.000 ;
    END
  END cache_entry[30]
  PIN cache_entry[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 340.490 796.000 340.770 800.000 ;
    END
  END cache_entry[31]
  PIN cache_entry[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 345.550 796.000 345.830 800.000 ;
    END
  END cache_entry[32]
  PIN cache_entry[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 350.610 796.000 350.890 800.000 ;
    END
  END cache_entry[33]
  PIN cache_entry[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 355.670 796.000 355.950 800.000 ;
    END
  END cache_entry[34]
  PIN cache_entry[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 360.730 796.000 361.010 800.000 ;
    END
  END cache_entry[35]
  PIN cache_entry[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 365.790 796.000 366.070 800.000 ;
    END
  END cache_entry[36]
  PIN cache_entry[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 370.850 796.000 371.130 800.000 ;
    END
  END cache_entry[37]
  PIN cache_entry[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 375.910 796.000 376.190 800.000 ;
    END
  END cache_entry[38]
  PIN cache_entry[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 380.970 796.000 381.250 800.000 ;
    END
  END cache_entry[39]
  PIN cache_entry[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 198.810 796.000 199.090 800.000 ;
    END
  END cache_entry[3]
  PIN cache_entry[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 386.030 796.000 386.310 800.000 ;
    END
  END cache_entry[40]
  PIN cache_entry[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 391.090 796.000 391.370 800.000 ;
    END
  END cache_entry[41]
  PIN cache_entry[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 396.150 796.000 396.430 800.000 ;
    END
  END cache_entry[42]
  PIN cache_entry[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 401.210 796.000 401.490 800.000 ;
    END
  END cache_entry[43]
  PIN cache_entry[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 406.270 796.000 406.550 800.000 ;
    END
  END cache_entry[44]
  PIN cache_entry[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 411.330 796.000 411.610 800.000 ;
    END
  END cache_entry[45]
  PIN cache_entry[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 416.390 796.000 416.670 800.000 ;
    END
  END cache_entry[46]
  PIN cache_entry[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 421.450 796.000 421.730 800.000 ;
    END
  END cache_entry[47]
  PIN cache_entry[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 426.510 796.000 426.790 800.000 ;
    END
  END cache_entry[48]
  PIN cache_entry[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 431.570 796.000 431.850 800.000 ;
    END
  END cache_entry[49]
  PIN cache_entry[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 203.870 796.000 204.150 800.000 ;
    END
  END cache_entry[4]
  PIN cache_entry[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 436.630 796.000 436.910 800.000 ;
    END
  END cache_entry[50]
  PIN cache_entry[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 441.690 796.000 441.970 800.000 ;
    END
  END cache_entry[51]
  PIN cache_entry[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 446.750 796.000 447.030 800.000 ;
    END
  END cache_entry[52]
  PIN cache_entry[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 451.810 796.000 452.090 800.000 ;
    END
  END cache_entry[53]
  PIN cache_entry[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 456.870 796.000 457.150 800.000 ;
    END
  END cache_entry[54]
  PIN cache_entry[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 461.930 796.000 462.210 800.000 ;
    END
  END cache_entry[55]
  PIN cache_entry[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 466.990 796.000 467.270 800.000 ;
    END
  END cache_entry[56]
  PIN cache_entry[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 472.050 796.000 472.330 800.000 ;
    END
  END cache_entry[57]
  PIN cache_entry[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 477.110 796.000 477.390 800.000 ;
    END
  END cache_entry[58]
  PIN cache_entry[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 482.170 796.000 482.450 800.000 ;
    END
  END cache_entry[59]
  PIN cache_entry[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 208.930 796.000 209.210 800.000 ;
    END
  END cache_entry[5]
  PIN cache_entry[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 487.230 796.000 487.510 800.000 ;
    END
  END cache_entry[60]
  PIN cache_entry[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 492.290 796.000 492.570 800.000 ;
    END
  END cache_entry[61]
  PIN cache_entry[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 497.350 796.000 497.630 800.000 ;
    END
  END cache_entry[62]
  PIN cache_entry[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 502.410 796.000 502.690 800.000 ;
    END
  END cache_entry[63]
  PIN cache_entry[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 507.470 796.000 507.750 800.000 ;
    END
  END cache_entry[64]
  PIN cache_entry[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 512.530 796.000 512.810 800.000 ;
    END
  END cache_entry[65]
  PIN cache_entry[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 517.590 796.000 517.870 800.000 ;
    END
  END cache_entry[66]
  PIN cache_entry[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 522.650 796.000 522.930 800.000 ;
    END
  END cache_entry[67]
  PIN cache_entry[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 527.710 796.000 527.990 800.000 ;
    END
  END cache_entry[68]
  PIN cache_entry[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 532.770 796.000 533.050 800.000 ;
    END
  END cache_entry[69]
  PIN cache_entry[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 213.990 796.000 214.270 800.000 ;
    END
  END cache_entry[6]
  PIN cache_entry[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 537.830 796.000 538.110 800.000 ;
    END
  END cache_entry[70]
  PIN cache_entry[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 542.890 796.000 543.170 800.000 ;
    END
  END cache_entry[71]
  PIN cache_entry[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 547.950 796.000 548.230 800.000 ;
    END
  END cache_entry[72]
  PIN cache_entry[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 553.010 796.000 553.290 800.000 ;
    END
  END cache_entry[73]
  PIN cache_entry[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 558.070 796.000 558.350 800.000 ;
    END
  END cache_entry[74]
  PIN cache_entry[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 563.130 796.000 563.410 800.000 ;
    END
  END cache_entry[75]
  PIN cache_entry[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 568.190 796.000 568.470 800.000 ;
    END
  END cache_entry[76]
  PIN cache_entry[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 573.250 796.000 573.530 800.000 ;
    END
  END cache_entry[77]
  PIN cache_entry[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 578.310 796.000 578.590 800.000 ;
    END
  END cache_entry[78]
  PIN cache_entry[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 583.370 796.000 583.650 800.000 ;
    END
  END cache_entry[79]
  PIN cache_entry[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 219.050 796.000 219.330 800.000 ;
    END
  END cache_entry[7]
  PIN cache_entry[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 588.430 796.000 588.710 800.000 ;
    END
  END cache_entry[80]
  PIN cache_entry[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 593.490 796.000 593.770 800.000 ;
    END
  END cache_entry[81]
  PIN cache_entry[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 598.550 796.000 598.830 800.000 ;
    END
  END cache_entry[82]
  PIN cache_entry[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 603.610 796.000 603.890 800.000 ;
    END
  END cache_entry[83]
  PIN cache_entry[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 608.670 796.000 608.950 800.000 ;
    END
  END cache_entry[84]
  PIN cache_entry[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 613.730 796.000 614.010 800.000 ;
    END
  END cache_entry[85]
  PIN cache_entry[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 618.790 796.000 619.070 800.000 ;
    END
  END cache_entry[86]
  PIN cache_entry[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 623.850 796.000 624.130 800.000 ;
    END
  END cache_entry[87]
  PIN cache_entry[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 628.910 796.000 629.190 800.000 ;
    END
  END cache_entry[88]
  PIN cache_entry[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 633.970 796.000 634.250 800.000 ;
    END
  END cache_entry[89]
  PIN cache_entry[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 224.110 796.000 224.390 800.000 ;
    END
  END cache_entry[8]
  PIN cache_entry[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 639.030 796.000 639.310 800.000 ;
    END
  END cache_entry[90]
  PIN cache_entry[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 644.090 796.000 644.370 800.000 ;
    END
  END cache_entry[91]
  PIN cache_entry[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 649.150 796.000 649.430 800.000 ;
    END
  END cache_entry[92]
  PIN cache_entry[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 654.210 796.000 654.490 800.000 ;
    END
  END cache_entry[93]
  PIN cache_entry[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 659.270 796.000 659.550 800.000 ;
    END
  END cache_entry[94]
  PIN cache_entry[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 664.330 796.000 664.610 800.000 ;
    END
  END cache_entry[95]
  PIN cache_entry[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 669.390 796.000 669.670 800.000 ;
    END
  END cache_entry[96]
  PIN cache_entry[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 674.450 796.000 674.730 800.000 ;
    END
  END cache_entry[97]
  PIN cache_entry[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 679.510 796.000 679.790 800.000 ;
    END
  END cache_entry[98]
  PIN cache_entry[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 684.570 796.000 684.850 800.000 ;
    END
  END cache_entry[99]
  PIN cache_entry[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 229.170 796.000 229.450 800.000 ;
    END
  END cache_entry[9]
  PIN cache_entry_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.934000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 84.360 2200.000 84.960 ;
    END
  END cache_entry_valid
  PIN cache_hit
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 76.200 2200.000 76.800 ;
    END
  END cache_hit
  PIN cache_invalidate
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 78.920 2200.000 79.520 ;
    END
  END cache_invalidate
  PIN cache_new_entry[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 9.628200 ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END cache_new_entry[0]
  PIN cache_new_entry[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.489500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 915.950 0.000 916.230 4.000 ;
    END
  END cache_new_entry[100]
  PIN cache_new_entry[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.489500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 924.690 0.000 924.970 4.000 ;
    END
  END cache_new_entry[101]
  PIN cache_new_entry[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.489500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 933.430 0.000 933.710 4.000 ;
    END
  END cache_new_entry[102]
  PIN cache_new_entry[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.489500 ;
    ANTENNADIFFAREA 1.325700 ;
    PORT
      LAYER met2 ;
        RECT 942.170 0.000 942.450 4.000 ;
    END
  END cache_new_entry[103]
  PIN cache_new_entry[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.489500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 950.910 0.000 951.190 4.000 ;
    END
  END cache_new_entry[104]
  PIN cache_new_entry[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.489500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 959.650 0.000 959.930 4.000 ;
    END
  END cache_new_entry[105]
  PIN cache_new_entry[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.489500 ;
    ANTENNADIFFAREA 1.325700 ;
    PORT
      LAYER met2 ;
        RECT 968.390 0.000 968.670 4.000 ;
    END
  END cache_new_entry[106]
  PIN cache_new_entry[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.489500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 977.130 0.000 977.410 4.000 ;
    END
  END cache_new_entry[107]
  PIN cache_new_entry[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.489500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 985.870 0.000 986.150 4.000 ;
    END
  END cache_new_entry[108]
  PIN cache_new_entry[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.489500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 994.610 0.000 994.890 4.000 ;
    END
  END cache_new_entry[109]
  PIN cache_new_entry[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.363500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 129.350 0.000 129.630 4.000 ;
    END
  END cache_new_entry[10]
  PIN cache_new_entry[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.621000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1003.350 0.000 1003.630 4.000 ;
    END
  END cache_new_entry[110]
  PIN cache_new_entry[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.747000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1012.090 0.000 1012.370 4.000 ;
    END
  END cache_new_entry[111]
  PIN cache_new_entry[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1020.830 0.000 1021.110 4.000 ;
    END
  END cache_new_entry[112]
  PIN cache_new_entry[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1029.570 0.000 1029.850 4.000 ;
    END
  END cache_new_entry[113]
  PIN cache_new_entry[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1038.310 0.000 1038.590 4.000 ;
    END
  END cache_new_entry[114]
  PIN cache_new_entry[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1047.050 0.000 1047.330 4.000 ;
    END
  END cache_new_entry[115]
  PIN cache_new_entry[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1055.790 0.000 1056.070 4.000 ;
    END
  END cache_new_entry[116]
  PIN cache_new_entry[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1064.530 0.000 1064.810 4.000 ;
    END
  END cache_new_entry[117]
  PIN cache_new_entry[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1073.270 0.000 1073.550 4.000 ;
    END
  END cache_new_entry[118]
  PIN cache_new_entry[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1082.010 0.000 1082.290 4.000 ;
    END
  END cache_new_entry[119]
  PIN cache_new_entry[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.186500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 138.090 0.000 138.370 4.000 ;
    END
  END cache_new_entry[11]
  PIN cache_new_entry[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1090.750 0.000 1091.030 4.000 ;
    END
  END cache_new_entry[120]
  PIN cache_new_entry[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1099.490 0.000 1099.770 4.000 ;
    END
  END cache_new_entry[121]
  PIN cache_new_entry[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1108.230 0.000 1108.510 4.000 ;
    END
  END cache_new_entry[122]
  PIN cache_new_entry[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1116.970 0.000 1117.250 4.000 ;
    END
  END cache_new_entry[123]
  PIN cache_new_entry[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1125.710 0.000 1125.990 4.000 ;
    END
  END cache_new_entry[124]
  PIN cache_new_entry[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1134.450 0.000 1134.730 4.000 ;
    END
  END cache_new_entry[125]
  PIN cache_new_entry[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1143.190 0.000 1143.470 4.000 ;
    END
  END cache_new_entry[126]
  PIN cache_new_entry[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1151.930 0.000 1152.210 4.000 ;
    END
  END cache_new_entry[127]
  PIN cache_new_entry[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.186500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 146.830 0.000 147.110 4.000 ;
    END
  END cache_new_entry[12]
  PIN cache_new_entry[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.363500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 155.570 0.000 155.850 4.000 ;
    END
  END cache_new_entry[13]
  PIN cache_new_entry[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.186500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 4.000 ;
    END
  END cache_new_entry[14]
  PIN cache_new_entry[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 173.050 0.000 173.330 4.000 ;
    END
  END cache_new_entry[15]
  PIN cache_new_entry[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.186500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 181.790 0.000 182.070 4.000 ;
    END
  END cache_new_entry[16]
  PIN cache_new_entry[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.186500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 190.530 0.000 190.810 4.000 ;
    END
  END cache_new_entry[17]
  PIN cache_new_entry[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 199.270 0.000 199.550 4.000 ;
    END
  END cache_new_entry[18]
  PIN cache_new_entry[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 208.010 0.000 208.290 4.000 ;
    END
  END cache_new_entry[19]
  PIN cache_new_entry[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.186500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 50.690 0.000 50.970 4.000 ;
    END
  END cache_new_entry[1]
  PIN cache_new_entry[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.186500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 216.750 0.000 217.030 4.000 ;
    END
  END cache_new_entry[20]
  PIN cache_new_entry[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 4.000 ;
    END
  END cache_new_entry[21]
  PIN cache_new_entry[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.186500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 234.230 0.000 234.510 4.000 ;
    END
  END cache_new_entry[22]
  PIN cache_new_entry[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.186500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 242.970 0.000 243.250 4.000 ;
    END
  END cache_new_entry[23]
  PIN cache_new_entry[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.186500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 251.710 0.000 251.990 4.000 ;
    END
  END cache_new_entry[24]
  PIN cache_new_entry[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.186500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 260.450 0.000 260.730 4.000 ;
    END
  END cache_new_entry[25]
  PIN cache_new_entry[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.048500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 269.190 0.000 269.470 4.000 ;
    END
  END cache_new_entry[26]
  PIN cache_new_entry[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.186500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 277.930 0.000 278.210 4.000 ;
    END
  END cache_new_entry[27]
  PIN cache_new_entry[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.186500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 286.670 0.000 286.950 4.000 ;
    END
  END cache_new_entry[28]
  PIN cache_new_entry[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.363500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 295.410 0.000 295.690 4.000 ;
    END
  END cache_new_entry[29]
  PIN cache_new_entry[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.363500 ;
    ANTENNADIFFAREA 2.629800 ;
    PORT
      LAYER met2 ;
        RECT 59.430 0.000 59.710 4.000 ;
    END
  END cache_new_entry[2]
  PIN cache_new_entry[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.186500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 304.150 0.000 304.430 4.000 ;
    END
  END cache_new_entry[30]
  PIN cache_new_entry[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.363500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 312.890 0.000 313.170 4.000 ;
    END
  END cache_new_entry[31]
  PIN cache_new_entry[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.363500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 321.630 0.000 321.910 4.000 ;
    END
  END cache_new_entry[32]
  PIN cache_new_entry[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.363500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 330.370 0.000 330.650 4.000 ;
    END
  END cache_new_entry[33]
  PIN cache_new_entry[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.363500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 339.110 0.000 339.390 4.000 ;
    END
  END cache_new_entry[34]
  PIN cache_new_entry[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.363500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 347.850 0.000 348.130 4.000 ;
    END
  END cache_new_entry[35]
  PIN cache_new_entry[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.363500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 356.590 0.000 356.870 4.000 ;
    END
  END cache_new_entry[36]
  PIN cache_new_entry[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.363500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 365.330 0.000 365.610 4.000 ;
    END
  END cache_new_entry[37]
  PIN cache_new_entry[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.363500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 374.070 0.000 374.350 4.000 ;
    END
  END cache_new_entry[38]
  PIN cache_new_entry[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.363500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 382.810 0.000 383.090 4.000 ;
    END
  END cache_new_entry[39]
  PIN cache_new_entry[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.186500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 68.170 0.000 68.450 4.000 ;
    END
  END cache_new_entry[3]
  PIN cache_new_entry[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 391.550 0.000 391.830 4.000 ;
    END
  END cache_new_entry[40]
  PIN cache_new_entry[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.363500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 400.290 0.000 400.570 4.000 ;
    END
  END cache_new_entry[41]
  PIN cache_new_entry[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.186500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 409.030 0.000 409.310 4.000 ;
    END
  END cache_new_entry[42]
  PIN cache_new_entry[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.186500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 417.770 0.000 418.050 4.000 ;
    END
  END cache_new_entry[43]
  PIN cache_new_entry[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.363500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 426.510 0.000 426.790 4.000 ;
    END
  END cache_new_entry[44]
  PIN cache_new_entry[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.203000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 435.250 0.000 435.530 4.000 ;
    END
  END cache_new_entry[45]
  PIN cache_new_entry[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.363500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 443.990 0.000 444.270 4.000 ;
    END
  END cache_new_entry[46]
  PIN cache_new_entry[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.203000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 452.730 0.000 453.010 4.000 ;
    END
  END cache_new_entry[47]
  PIN cache_new_entry[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.203000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 461.470 0.000 461.750 4.000 ;
    END
  END cache_new_entry[48]
  PIN cache_new_entry[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.186500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 470.210 0.000 470.490 4.000 ;
    END
  END cache_new_entry[49]
  PIN cache_new_entry[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.363500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 76.910 0.000 77.190 4.000 ;
    END
  END cache_new_entry[4]
  PIN cache_new_entry[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.186500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 478.950 0.000 479.230 4.000 ;
    END
  END cache_new_entry[50]
  PIN cache_new_entry[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.149000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 487.690 0.000 487.970 4.000 ;
    END
  END cache_new_entry[51]
  PIN cache_new_entry[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 496.430 0.000 496.710 4.000 ;
    END
  END cache_new_entry[52]
  PIN cache_new_entry[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.186500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 505.170 0.000 505.450 4.000 ;
    END
  END cache_new_entry[53]
  PIN cache_new_entry[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.186500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 513.910 0.000 514.190 4.000 ;
    END
  END cache_new_entry[54]
  PIN cache_new_entry[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.186500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 522.650 0.000 522.930 4.000 ;
    END
  END cache_new_entry[55]
  PIN cache_new_entry[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 531.390 0.000 531.670 4.000 ;
    END
  END cache_new_entry[56]
  PIN cache_new_entry[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.186500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 540.130 0.000 540.410 4.000 ;
    END
  END cache_new_entry[57]
  PIN cache_new_entry[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.363500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 548.870 0.000 549.150 4.000 ;
    END
  END cache_new_entry[58]
  PIN cache_new_entry[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.363500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 557.610 0.000 557.890 4.000 ;
    END
  END cache_new_entry[59]
  PIN cache_new_entry[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.186500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 85.650 0.000 85.930 4.000 ;
    END
  END cache_new_entry[5]
  PIN cache_new_entry[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.363500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 566.350 0.000 566.630 4.000 ;
    END
  END cache_new_entry[60]
  PIN cache_new_entry[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.363500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 575.090 0.000 575.370 4.000 ;
    END
  END cache_new_entry[61]
  PIN cache_new_entry[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.363500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 583.830 0.000 584.110 4.000 ;
    END
  END cache_new_entry[62]
  PIN cache_new_entry[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.186500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 592.570 0.000 592.850 4.000 ;
    END
  END cache_new_entry[63]
  PIN cache_new_entry[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.363500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 601.310 0.000 601.590 4.000 ;
    END
  END cache_new_entry[64]
  PIN cache_new_entry[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.149000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 610.050 0.000 610.330 4.000 ;
    END
  END cache_new_entry[65]
  PIN cache_new_entry[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.149000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 618.790 0.000 619.070 4.000 ;
    END
  END cache_new_entry[66]
  PIN cache_new_entry[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 627.530 0.000 627.810 4.000 ;
    END
  END cache_new_entry[67]
  PIN cache_new_entry[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.203000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 636.270 0.000 636.550 4.000 ;
    END
  END cache_new_entry[68]
  PIN cache_new_entry[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.149000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 645.010 0.000 645.290 4.000 ;
    END
  END cache_new_entry[69]
  PIN cache_new_entry[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.186500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 94.390 0.000 94.670 4.000 ;
    END
  END cache_new_entry[6]
  PIN cache_new_entry[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 1.760400 ;
    PORT
      LAYER met2 ;
        RECT 653.750 0.000 654.030 4.000 ;
    END
  END cache_new_entry[70]
  PIN cache_new_entry[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.149000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 662.490 0.000 662.770 4.000 ;
    END
  END cache_new_entry[71]
  PIN cache_new_entry[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.485000 ;
    ANTENNADIFFAREA 1.325700 ;
    PORT
      LAYER met2 ;
        RECT 671.230 0.000 671.510 4.000 ;
    END
  END cache_new_entry[72]
  PIN cache_new_entry[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.203000 ;
    ANTENNADIFFAREA 1.325700 ;
    PORT
      LAYER met2 ;
        RECT 679.970 0.000 680.250 4.000 ;
    END
  END cache_new_entry[73]
  PIN cache_new_entry[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.149000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 688.710 0.000 688.990 4.000 ;
    END
  END cache_new_entry[74]
  PIN cache_new_entry[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.149000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 697.450 0.000 697.730 4.000 ;
    END
  END cache_new_entry[75]
  PIN cache_new_entry[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.485000 ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 706.190 0.000 706.470 4.000 ;
    END
  END cache_new_entry[76]
  PIN cache_new_entry[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.203000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 714.930 0.000 715.210 4.000 ;
    END
  END cache_new_entry[77]
  PIN cache_new_entry[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 723.670 0.000 723.950 4.000 ;
    END
  END cache_new_entry[78]
  PIN cache_new_entry[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 1.760400 ;
    PORT
      LAYER met2 ;
        RECT 732.410 0.000 732.690 4.000 ;
    END
  END cache_new_entry[79]
  PIN cache_new_entry[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.186500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END cache_new_entry[7]
  PIN cache_new_entry[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 741.150 0.000 741.430 4.000 ;
    END
  END cache_new_entry[80]
  PIN cache_new_entry[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.737000 ;
    ANTENNADIFFAREA 2.629800 ;
    PORT
      LAYER met2 ;
        RECT 749.890 0.000 750.170 4.000 ;
    END
  END cache_new_entry[81]
  PIN cache_new_entry[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.737000 ;
    ANTENNADIFFAREA 2.629800 ;
    PORT
      LAYER met2 ;
        RECT 758.630 0.000 758.910 4.000 ;
    END
  END cache_new_entry[82]
  PIN cache_new_entry[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.737000 ;
    ANTENNADIFFAREA 1.325700 ;
    PORT
      LAYER met2 ;
        RECT 767.370 0.000 767.650 4.000 ;
    END
  END cache_new_entry[83]
  PIN cache_new_entry[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.737000 ;
    ANTENNADIFFAREA 1.760400 ;
    PORT
      LAYER met2 ;
        RECT 776.110 0.000 776.390 4.000 ;
    END
  END cache_new_entry[84]
  PIN cache_new_entry[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.737000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 784.850 0.000 785.130 4.000 ;
    END
  END cache_new_entry[85]
  PIN cache_new_entry[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.737000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 793.590 0.000 793.870 4.000 ;
    END
  END cache_new_entry[86]
  PIN cache_new_entry[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 802.330 0.000 802.610 4.000 ;
    END
  END cache_new_entry[87]
  PIN cache_new_entry[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.737000 ;
    ANTENNADIFFAREA 2.195100 ;
    PORT
      LAYER met2 ;
        RECT 811.070 0.000 811.350 4.000 ;
    END
  END cache_new_entry[88]
  PIN cache_new_entry[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.737000 ;
    ANTENNADIFFAREA 1.325700 ;
    PORT
      LAYER met2 ;
        RECT 819.810 0.000 820.090 4.000 ;
    END
  END cache_new_entry[89]
  PIN cache_new_entry[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.186500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 111.870 0.000 112.150 4.000 ;
    END
  END cache_new_entry[8]
  PIN cache_new_entry[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.737000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 828.550 0.000 828.830 4.000 ;
    END
  END cache_new_entry[90]
  PIN cache_new_entry[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.737000 ;
    ANTENNADIFFAREA 1.760400 ;
    PORT
      LAYER met2 ;
        RECT 837.290 0.000 837.570 4.000 ;
    END
  END cache_new_entry[91]
  PIN cache_new_entry[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 846.030 0.000 846.310 4.000 ;
    END
  END cache_new_entry[92]
  PIN cache_new_entry[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.737000 ;
    ANTENNADIFFAREA 2.629800 ;
    PORT
      LAYER met2 ;
        RECT 854.770 0.000 855.050 4.000 ;
    END
  END cache_new_entry[93]
  PIN cache_new_entry[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.737000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 863.510 0.000 863.790 4.000 ;
    END
  END cache_new_entry[94]
  PIN cache_new_entry[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.351500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 872.250 0.000 872.530 4.000 ;
    END
  END cache_new_entry[95]
  PIN cache_new_entry[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.368000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 880.990 0.000 881.270 4.000 ;
    END
  END cache_new_entry[96]
  PIN cache_new_entry[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.489500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 889.730 0.000 890.010 4.000 ;
    END
  END cache_new_entry[97]
  PIN cache_new_entry[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.489500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 898.470 0.000 898.750 4.000 ;
    END
  END cache_new_entry[98]
  PIN cache_new_entry[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.489500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 907.210 0.000 907.490 4.000 ;
    END
  END cache_new_entry[99]
  PIN cache_new_entry[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.186500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 120.610 0.000 120.890 4.000 ;
    END
  END cache_new_entry[9]
  PIN cache_rst
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 81.640 2200.000 82.240 ;
    END
  END cache_rst
  PIN curr_PC[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.343500 ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 836.370 796.000 836.650 800.000 ;
    END
  END curr_PC[0]
  PIN curr_PC[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.223500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 886.970 796.000 887.250 800.000 ;
    END
  END curr_PC[10]
  PIN curr_PC[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.486500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 892.030 796.000 892.310 800.000 ;
    END
  END curr_PC[11]
  PIN curr_PC[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.365000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 897.090 796.000 897.370 800.000 ;
    END
  END curr_PC[12]
  PIN curr_PC[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.608000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 902.150 796.000 902.430 800.000 ;
    END
  END curr_PC[13]
  PIN curr_PC[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.971500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 907.210 796.000 907.490 800.000 ;
    END
  END curr_PC[14]
  PIN curr_PC[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.368000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 912.270 796.000 912.550 800.000 ;
    END
  END curr_PC[15]
  PIN curr_PC[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.084500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 917.330 796.000 917.610 800.000 ;
    END
  END curr_PC[16]
  PIN curr_PC[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.104500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 922.390 796.000 922.670 800.000 ;
    END
  END curr_PC[17]
  PIN curr_PC[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.837000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 927.450 796.000 927.730 800.000 ;
    END
  END curr_PC[18]
  PIN curr_PC[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.857000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 932.510 796.000 932.790 800.000 ;
    END
  END curr_PC[19]
  PIN curr_PC[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.608000 ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 841.430 796.000 841.710 800.000 ;
    END
  END curr_PC[1]
  PIN curr_PC[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.103000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 937.570 796.000 937.850 800.000 ;
    END
  END curr_PC[20]
  PIN curr_PC[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 942.630 796.000 942.910 800.000 ;
    END
  END curr_PC[21]
  PIN curr_PC[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.983000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 947.690 796.000 947.970 800.000 ;
    END
  END curr_PC[22]
  PIN curr_PC[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.081500 ;
    ANTENNADIFFAREA 1.760400 ;
    PORT
      LAYER met2 ;
        RECT 952.750 796.000 953.030 800.000 ;
    END
  END curr_PC[23]
  PIN curr_PC[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.204500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 957.810 796.000 958.090 800.000 ;
    END
  END curr_PC[24]
  PIN curr_PC[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.242000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 962.870 796.000 963.150 800.000 ;
    END
  END curr_PC[25]
  PIN curr_PC[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.727000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 967.930 796.000 968.210 800.000 ;
    END
  END curr_PC[26]
  PIN curr_PC[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.612500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 972.990 796.000 973.270 800.000 ;
    END
  END curr_PC[27]
  PIN curr_PC[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.967000 ;
    ANTENNADIFFAREA 3.542400 ;
    PORT
      LAYER met2 ;
        RECT 846.490 796.000 846.770 800.000 ;
    END
  END curr_PC[2]
  PIN curr_PC[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    ANTENNADIFFAREA 3.977100 ;
    PORT
      LAYER met2 ;
        RECT 851.550 796.000 851.830 800.000 ;
    END
  END curr_PC[3]
  PIN curr_PC[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.845500 ;
    ANTENNADIFFAREA 3.542400 ;
    PORT
      LAYER met2 ;
        RECT 856.610 796.000 856.890 800.000 ;
    END
  END curr_PC[4]
  PIN curr_PC[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.751500 ;
    ANTENNADIFFAREA 2.195100 ;
    PORT
      LAYER met2 ;
        RECT 861.670 796.000 861.950 800.000 ;
    END
  END curr_PC[5]
  PIN curr_PC[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.353500 ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 866.730 796.000 867.010 800.000 ;
    END
  END curr_PC[6]
  PIN curr_PC[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.789000 ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 871.790 796.000 872.070 800.000 ;
    END
  END curr_PC[7]
  PIN curr_PC[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.961500 ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 876.850 796.000 877.130 800.000 ;
    END
  END curr_PC[8]
  PIN curr_PC[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.984500 ;
    ANTENNADIFFAREA 4.846500 ;
    PORT
      LAYER met2 ;
        RECT 881.910 796.000 882.190 800.000 ;
    END
  END curr_PC[9]
  PIN custom_settings[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 2122.070 0.000 2122.350 4.000 ;
    END
  END custom_settings[0]
  PIN custom_settings[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met2 ;
        RECT 2130.810 0.000 2131.090 4.000 ;
    END
  END custom_settings[1]
  PIN custom_settings[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.719500 ;
    PORT
      LAYER met2 ;
        RECT 2139.550 0.000 2139.830 4.000 ;
    END
  END custom_settings[2]
  PIN custom_settings[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.719500 ;
    PORT
      LAYER met2 ;
        RECT 2148.290 0.000 2148.570 4.000 ;
    END
  END custom_settings[3]
  PIN custom_settings[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 2157.030 0.000 2157.310 4.000 ;
    END
  END custom_settings[4]
  PIN dest_idx0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1210.810 796.000 1211.090 800.000 ;
    END
  END dest_idx0[0]
  PIN dest_idx0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met2 ;
        RECT 1215.870 796.000 1216.150 800.000 ;
    END
  END dest_idx0[1]
  PIN dest_idx0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 1220.930 796.000 1221.210 800.000 ;
    END
  END dest_idx0[2]
  PIN dest_idx0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.237500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1225.990 796.000 1226.270 800.000 ;
    END
  END dest_idx0[3]
  PIN dest_idx0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 6.070500 ;
    PORT
      LAYER met2 ;
        RECT 1231.050 796.000 1231.330 800.000 ;
    END
  END dest_idx0[4]
  PIN dest_idx0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 6.691500 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met2 ;
        RECT 1236.110 796.000 1236.390 800.000 ;
    END
  END dest_idx0[5]
  PIN dest_idx1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 212.200 2200.000 212.800 ;
    END
  END dest_idx1[0]
  PIN dest_idx1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 7.308000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 214.920 2200.000 215.520 ;
    END
  END dest_idx1[1]
  PIN dest_idx1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 7.308000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 217.640 2200.000 218.240 ;
    END
  END dest_idx1[2]
  PIN dest_idx1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.242000 ;
    ANTENNADIFFAREA 7.824600 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 220.360 2200.000 220.960 ;
    END
  END dest_idx1[3]
  PIN dest_idx1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 223.080 2200.000 223.680 ;
    END
  END dest_idx1[4]
  PIN dest_idx1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 225.800 2200.000 226.400 ;
    END
  END dest_idx1[5]
  PIN dest_idx2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.901500 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.760 4.000 207.360 ;
    END
  END dest_idx2[0]
  PIN dest_idx2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.139000 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 209.480 4.000 210.080 ;
    END
  END dest_idx2[1]
  PIN dest_idx2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.017500 ;
    ANTENNADIFFAREA 2.173500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.200 4.000 212.800 ;
    END
  END dest_idx2[2]
  PIN dest_idx2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.353500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.920 4.000 215.520 ;
    END
  END dest_idx2[3]
  PIN dest_idx2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.611000 ;
    ANTENNADIFFAREA 2.173500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END dest_idx2[4]
  PIN dest_idx2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.858500 ;
    ANTENNADIFFAREA 4.347000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 220.360 4.000 220.960 ;
    END
  END dest_idx2[5]
  PIN dest_mask0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.485000 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met2 ;
        RECT 1200.690 796.000 1200.970 800.000 ;
    END
  END dest_mask0[0]
  PIN dest_mask0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.732500 ;
    PORT
      LAYER met2 ;
        RECT 1205.750 796.000 1206.030 800.000 ;
    END
  END dest_mask0[1]
  PIN dest_mask1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.485000 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 206.760 2200.000 207.360 ;
    END
  END dest_mask1[0]
  PIN dest_mask1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.732500 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 209.480 2200.000 210.080 ;
    END
  END dest_mask1[1]
  PIN dest_mask2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.207500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 201.320 4.000 201.920 ;
    END
  END dest_mask2[0]
  PIN dest_mask2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.838500 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
    END
  END dest_mask2[1]
  PIN dest_pred0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.882000 ;
    ANTENNADIFFAREA 3.042900 ;
    PORT
      LAYER met2 ;
        RECT 1256.350 796.000 1256.630 800.000 ;
    END
  END dest_pred0[0]
  PIN dest_pred0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.882000 ;
    ANTENNADIFFAREA 3.042900 ;
    PORT
      LAYER met2 ;
        RECT 1261.410 796.000 1261.690 800.000 ;
    END
  END dest_pred0[1]
  PIN dest_pred0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.882000 ;
    ANTENNADIFFAREA 3.042900 ;
    PORT
      LAYER met2 ;
        RECT 1266.470 796.000 1266.750 800.000 ;
    END
  END dest_pred0[2]
  PIN dest_pred1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.756000 ;
    ANTENNADIFFAREA 2.608200 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 236.680 2200.000 237.280 ;
    END
  END dest_pred1[0]
  PIN dest_pred1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.368000 ;
    ANTENNADIFFAREA 2.608200 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 239.400 2200.000 240.000 ;
    END
  END dest_pred1[1]
  PIN dest_pred1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.756000 ;
    ANTENNADIFFAREA 2.608200 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 242.120 2200.000 242.720 ;
    END
  END dest_pred1[2]
  PIN dest_pred2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.882000 ;
    ANTENNADIFFAREA 3.042900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.240 4.000 231.840 ;
    END
  END dest_pred2[0]
  PIN dest_pred2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.999000 ;
    ANTENNADIFFAREA 2.173500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 233.960 4.000 234.560 ;
    END
  END dest_pred2[1]
  PIN dest_pred2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.882000 ;
    ANTENNADIFFAREA 3.042900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.680 4.000 237.280 ;
    END
  END dest_pred2[2]
  PIN dest_pred_val0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.882000 ;
    ANTENNADIFFAREA 3.042900 ;
    PORT
      LAYER met2 ;
        RECT 1271.530 796.000 1271.810 800.000 ;
    END
  END dest_pred_val0
  PIN dest_pred_val1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.611000 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 244.840 2200.000 245.440 ;
    END
  END dest_pred_val1
  PIN dest_pred_val2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 3.042900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 239.400 4.000 240.000 ;
    END
  END dest_pred_val2
  PIN dest_val0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.485000 ;
    ANTENNADIFFAREA 3.477600 ;
    PORT
      LAYER met2 ;
        RECT 1038.770 796.000 1039.050 800.000 ;
    END
  END dest_val0[0]
  PIN dest_val0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.485000 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met2 ;
        RECT 1089.370 796.000 1089.650 800.000 ;
    END
  END dest_val0[10]
  PIN dest_val0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 1094.430 796.000 1094.710 800.000 ;
    END
  END dest_val0[11]
  PIN dest_val0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1099.490 796.000 1099.770 800.000 ;
    END
  END dest_val0[12]
  PIN dest_val0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.237500 ;
    PORT
      LAYER met2 ;
        RECT 1104.550 796.000 1104.830 800.000 ;
    END
  END dest_val0[13]
  PIN dest_val0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.327500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1109.610 796.000 1109.890 800.000 ;
    END
  END dest_val0[14]
  PIN dest_val0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.698000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1114.670 796.000 1114.950 800.000 ;
    END
  END dest_val0[15]
  PIN dest_val0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1119.730 796.000 1120.010 800.000 ;
    END
  END dest_val0[16]
  PIN dest_val0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.079500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1124.790 796.000 1125.070 800.000 ;
    END
  END dest_val0[17]
  PIN dest_val0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.594500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1129.850 796.000 1130.130 800.000 ;
    END
  END dest_val0[18]
  PIN dest_val0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1134.910 796.000 1135.190 800.000 ;
    END
  END dest_val0[19]
  PIN dest_val0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.594500 ;
    ANTENNADIFFAREA 4.347000 ;
    PORT
      LAYER met2 ;
        RECT 1043.830 796.000 1044.110 800.000 ;
    END
  END dest_val0[1]
  PIN dest_val0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.077500 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met2 ;
        RECT 1139.970 796.000 1140.250 800.000 ;
    END
  END dest_val0[20]
  PIN dest_val0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.945500 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met2 ;
        RECT 1145.030 796.000 1145.310 800.000 ;
    END
  END dest_val0[21]
  PIN dest_val0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.079500 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met2 ;
        RECT 1150.090 796.000 1150.370 800.000 ;
    END
  END dest_val0[22]
  PIN dest_val0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1155.150 796.000 1155.430 800.000 ;
    END
  END dest_val0[23]
  PIN dest_val0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.842000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1160.210 796.000 1160.490 800.000 ;
    END
  END dest_val0[24]
  PIN dest_val0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.079500 ;
    PORT
      LAYER met2 ;
        RECT 1165.270 796.000 1165.550 800.000 ;
    END
  END dest_val0[25]
  PIN dest_val0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.227500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1170.330 796.000 1170.610 800.000 ;
    END
  END dest_val0[26]
  PIN dest_val0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.694000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1175.390 796.000 1175.670 800.000 ;
    END
  END dest_val0[27]
  PIN dest_val0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.694000 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met2 ;
        RECT 1180.450 796.000 1180.730 800.000 ;
    END
  END dest_val0[28]
  PIN dest_val0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.832000 ;
    PORT
      LAYER met2 ;
        RECT 1185.510 796.000 1185.790 800.000 ;
    END
  END dest_val0[29]
  PIN dest_val0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.128500 ;
    ANTENNADIFFAREA 5.651100 ;
    PORT
      LAYER met2 ;
        RECT 1048.890 796.000 1049.170 800.000 ;
    END
  END dest_val0[2]
  PIN dest_val0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.217500 ;
    PORT
      LAYER met2 ;
        RECT 1190.570 796.000 1190.850 800.000 ;
    END
  END dest_val0[30]
  PIN dest_val0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.258000 ;
    PORT
      LAYER met2 ;
        RECT 1195.630 796.000 1195.910 800.000 ;
    END
  END dest_val0[31]
  PIN dest_val0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.242000 ;
    ANTENNADIFFAREA 2.608200 ;
    PORT
      LAYER met2 ;
        RECT 1053.950 796.000 1054.230 800.000 ;
    END
  END dest_val0[3]
  PIN dest_val0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1059.010 796.000 1059.290 800.000 ;
    END
  END dest_val0[4]
  PIN dest_val0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1064.070 796.000 1064.350 800.000 ;
    END
  END dest_val0[5]
  PIN dest_val0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.732500 ;
    ANTENNADIFFAREA 2.173500 ;
    PORT
      LAYER met2 ;
        RECT 1069.130 796.000 1069.410 800.000 ;
    END
  END dest_val0[6]
  PIN dest_val0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.485000 ;
    PORT
      LAYER met2 ;
        RECT 1074.190 796.000 1074.470 800.000 ;
    END
  END dest_val0[7]
  PIN dest_val0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.737000 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met2 ;
        RECT 1079.250 796.000 1079.530 800.000 ;
    END
  END dest_val0[8]
  PIN dest_val0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.789500 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met2 ;
        RECT 1084.310 796.000 1084.590 800.000 ;
    END
  END dest_val0[9]
  PIN dest_val1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.980000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 119.720 2200.000 120.320 ;
    END
  END dest_val1[0]
  PIN dest_val1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.732500 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 146.920 2200.000 147.520 ;
    END
  END dest_val1[10]
  PIN dest_val1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 149.640 2200.000 150.240 ;
    END
  END dest_val1[11]
  PIN dest_val1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.237500 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 152.360 2200.000 152.960 ;
    END
  END dest_val1[12]
  PIN dest_val1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.921000 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 155.080 2200.000 155.680 ;
    END
  END dest_val1[13]
  PIN dest_val1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.901500 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 157.800 2200.000 158.400 ;
    END
  END dest_val1[14]
  PIN dest_val1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.149000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 160.520 2200.000 161.120 ;
    END
  END dest_val1[15]
  PIN dest_val1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.958000 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 163.240 2200.000 163.840 ;
    END
  END dest_val1[16]
  PIN dest_val1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 165.960 2200.000 166.560 ;
    END
  END dest_val1[17]
  PIN dest_val1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.347000 ;
    ANTENNADIFFAREA 4.347000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 168.680 2200.000 169.280 ;
    END
  END dest_val1[18]
  PIN dest_val1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.465000 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 171.400 2200.000 172.000 ;
    END
  END dest_val1[19]
  PIN dest_val1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.089500 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 122.440 2200.000 123.040 ;
    END
  END dest_val1[1]
  PIN dest_val1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.164500 ;
    ANTENNADIFFAREA 5.216400 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 174.120 2200.000 174.720 ;
    END
  END dest_val1[20]
  PIN dest_val1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.945500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 176.840 2200.000 177.440 ;
    END
  END dest_val1[21]
  PIN dest_val1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.079500 ;
    ANTENNADIFFAREA 2.608200 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 179.560 2200.000 180.160 ;
    END
  END dest_val1[22]
  PIN dest_val1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807500 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 182.280 2200.000 182.880 ;
    END
  END dest_val1[23]
  PIN dest_val1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.732500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 185.000 2200.000 185.600 ;
    END
  END dest_val1[24]
  PIN dest_val1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.079500 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 187.720 2200.000 188.320 ;
    END
  END dest_val1[25]
  PIN dest_val1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.475000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 190.440 2200.000 191.040 ;
    END
  END dest_val1[26]
  PIN dest_val1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.584500 ;
    ANTENNADIFFAREA 3.912300 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 193.160 2200.000 193.760 ;
    END
  END dest_val1[27]
  PIN dest_val1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.694000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 195.880 2200.000 196.480 ;
    END
  END dest_val1[28]
  PIN dest_val1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.832000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 198.600 2200.000 199.200 ;
    END
  END dest_val1[29]
  PIN dest_val1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.950000 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 125.160 2200.000 125.760 ;
    END
  END dest_val1[2]
  PIN dest_val1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.327000 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 201.320 2200.000 201.920 ;
    END
  END dest_val1[30]
  PIN dest_val1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.258000 ;
    ANTENNADIFFAREA 2.608200 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 204.040 2200.000 204.640 ;
    END
  END dest_val1[31]
  PIN dest_val1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.420500 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 127.880 2200.000 128.480 ;
    END
  END dest_val1[3]
  PIN dest_val1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 130.600 2200.000 131.200 ;
    END
  END dest_val1[4]
  PIN dest_val1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.416000 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 133.320 2200.000 133.920 ;
    END
  END dest_val1[5]
  PIN dest_val1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 136.040 2200.000 136.640 ;
    END
  END dest_val1[6]
  PIN dest_val1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.485000 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 138.760 2200.000 139.360 ;
    END
  END dest_val1[7]
  PIN dest_val1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.737000 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 141.480 2200.000 142.080 ;
    END
  END dest_val1[8]
  PIN dest_val1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.037000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 144.200 2200.000 144.800 ;
    END
  END dest_val1[9]
  PIN dest_val2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 10.867499 ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.280 4.000 114.880 ;
    END
  END dest_val2[0]
  PIN dest_val2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 141.480 4.000 142.080 ;
    END
  END dest_val2[10]
  PIN dest_val2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 144.200 4.000 144.800 ;
    END
  END dest_val2[11]
  PIN dest_val2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 3.477600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.920 4.000 147.520 ;
    END
  END dest_val2[12]
  PIN dest_val2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END dest_val2[13]
  PIN dest_val2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 3.042900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 152.360 4.000 152.960 ;
    END
  END dest_val2[14]
  PIN dest_val2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 3.477600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.080 4.000 155.680 ;
    END
  END dest_val2[15]
  PIN dest_val2[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.800 4.000 158.400 ;
    END
  END dest_val2[16]
  PIN dest_val2[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 160.520 4.000 161.120 ;
    END
  END dest_val2[17]
  PIN dest_val2[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END dest_val2[18]
  PIN dest_val2[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.960 4.000 166.560 ;
    END
  END dest_val2[19]
  PIN dest_val2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    ANTENNADIFFAREA 3.912300 ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.000 4.000 117.600 ;
    END
  END dest_val2[1]
  PIN dest_val2[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.680 4.000 169.280 ;
    END
  END dest_val2[20]
  PIN dest_val2[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 2.608200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 171.400 4.000 172.000 ;
    END
  END dest_val2[21]
  PIN dest_val2[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 2.608200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.120 4.000 174.720 ;
    END
  END dest_val2[22]
  PIN dest_val2[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END dest_val2[23]
  PIN dest_val2[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 0.000 179.560 4.000 180.160 ;
    END
  END dest_val2[24]
  PIN dest_val2[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 182.280 4.000 182.880 ;
    END
  END dest_val2[25]
  PIN dest_val2[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.000 4.000 185.600 ;
    END
  END dest_val2[26]
  PIN dest_val2[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 2.173500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.720 4.000 188.320 ;
    END
  END dest_val2[27]
  PIN dest_val2[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 4.000 191.040 ;
    END
  END dest_val2[28]
  PIN dest_val2[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    ANTENNADIFFAREA 2.608200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.160 4.000 193.760 ;
    END
  END dest_val2[29]
  PIN dest_val2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.720 4.000 120.320 ;
    END
  END dest_val2[2]
  PIN dest_val2[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 2.608200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.880 4.000 196.480 ;
    END
  END dest_val2[30]
  PIN dest_val2[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 198.600 4.000 199.200 ;
    END
  END dest_val2[31]
  PIN dest_val2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    ANTENNADIFFAREA 3.912300 ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END dest_val2[3]
  PIN dest_val2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.160 4.000 125.760 ;
    END
  END dest_val2[4]
  PIN dest_val2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    ANTENNADIFFAREA 3.912300 ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.880 4.000 128.480 ;
    END
  END dest_val2[5]
  PIN dest_val2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    ANTENNADIFFAREA 3.042900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.600 4.000 131.200 ;
    END
  END dest_val2[6]
  PIN dest_val2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 0.000 133.320 4.000 133.920 ;
    END
  END dest_val2[7]
  PIN dest_val2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END dest_val2[8]
  PIN dest_val2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.760 4.000 139.360 ;
    END
  END dest_val2[9]
  PIN eu0_busy
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.621000 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met2 ;
        RECT 1610.550 796.000 1610.830 800.000 ;
    END
  END eu0_busy
  PIN eu0_instruction[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 15.670799 ;
    PORT
      LAYER met2 ;
        RECT 1615.610 796.000 1615.890 800.000 ;
    END
  END eu0_instruction[0]
  PIN eu0_instruction[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 10.454400 ;
    PORT
      LAYER met2 ;
        RECT 1666.210 796.000 1666.490 800.000 ;
    END
  END eu0_instruction[10]
  PIN eu0_instruction[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 10.454400 ;
    PORT
      LAYER met2 ;
        RECT 1671.270 796.000 1671.550 800.000 ;
    END
  END eu0_instruction[11]
  PIN eu0_instruction[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1676.330 796.000 1676.610 800.000 ;
    END
  END eu0_instruction[12]
  PIN eu0_instruction[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 10.454400 ;
    PORT
      LAYER met2 ;
        RECT 1681.390 796.000 1681.670 800.000 ;
    END
  END eu0_instruction[13]
  PIN eu0_instruction[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 10.454400 ;
    PORT
      LAYER met2 ;
        RECT 1686.450 796.000 1686.730 800.000 ;
    END
  END eu0_instruction[14]
  PIN eu0_instruction[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1691.510 796.000 1691.790 800.000 ;
    END
  END eu0_instruction[15]
  PIN eu0_instruction[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1696.570 796.000 1696.850 800.000 ;
    END
  END eu0_instruction[16]
  PIN eu0_instruction[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1701.630 796.000 1701.910 800.000 ;
    END
  END eu0_instruction[17]
  PIN eu0_instruction[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1706.690 796.000 1706.970 800.000 ;
    END
  END eu0_instruction[18]
  PIN eu0_instruction[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1711.750 796.000 1712.030 800.000 ;
    END
  END eu0_instruction[19]
  PIN eu0_instruction[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 41.752800 ;
    PORT
      LAYER met2 ;
        RECT 1620.670 796.000 1620.950 800.000 ;
    END
  END eu0_instruction[1]
  PIN eu0_instruction[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1716.810 796.000 1717.090 800.000 ;
    END
  END eu0_instruction[20]
  PIN eu0_instruction[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1721.870 796.000 1722.150 800.000 ;
    END
  END eu0_instruction[21]
  PIN eu0_instruction[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1726.930 796.000 1727.210 800.000 ;
    END
  END eu0_instruction[22]
  PIN eu0_instruction[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1731.990 796.000 1732.270 800.000 ;
    END
  END eu0_instruction[23]
  PIN eu0_instruction[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1737.050 796.000 1737.330 800.000 ;
    END
  END eu0_instruction[24]
  PIN eu0_instruction[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1742.110 796.000 1742.390 800.000 ;
    END
  END eu0_instruction[25]
  PIN eu0_instruction[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1747.170 796.000 1747.450 800.000 ;
    END
  END eu0_instruction[26]
  PIN eu0_instruction[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1752.230 796.000 1752.510 800.000 ;
    END
  END eu0_instruction[27]
  PIN eu0_instruction[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1757.290 796.000 1757.570 800.000 ;
    END
  END eu0_instruction[28]
  PIN eu0_instruction[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1762.350 796.000 1762.630 800.000 ;
    END
  END eu0_instruction[29]
  PIN eu0_instruction[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 20.887199 ;
    PORT
      LAYER met2 ;
        RECT 1625.730 796.000 1626.010 800.000 ;
    END
  END eu0_instruction[2]
  PIN eu0_instruction[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1767.410 796.000 1767.690 800.000 ;
    END
  END eu0_instruction[30]
  PIN eu0_instruction[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1772.470 796.000 1772.750 800.000 ;
    END
  END eu0_instruction[31]
  PIN eu0_instruction[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1777.530 796.000 1777.810 800.000 ;
    END
  END eu0_instruction[32]
  PIN eu0_instruction[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1782.590 796.000 1782.870 800.000 ;
    END
  END eu0_instruction[33]
  PIN eu0_instruction[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1787.650 796.000 1787.930 800.000 ;
    END
  END eu0_instruction[34]
  PIN eu0_instruction[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1792.710 796.000 1792.990 800.000 ;
    END
  END eu0_instruction[35]
  PIN eu0_instruction[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1797.770 796.000 1798.050 800.000 ;
    END
  END eu0_instruction[36]
  PIN eu0_instruction[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1802.830 796.000 1803.110 800.000 ;
    END
  END eu0_instruction[37]
  PIN eu0_instruction[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1807.890 796.000 1808.170 800.000 ;
    END
  END eu0_instruction[38]
  PIN eu0_instruction[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1812.950 796.000 1813.230 800.000 ;
    END
  END eu0_instruction[39]
  PIN eu0_instruction[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 10.454400 ;
    PORT
      LAYER met2 ;
        RECT 1630.790 796.000 1631.070 800.000 ;
    END
  END eu0_instruction[3]
  PIN eu0_instruction[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1818.010 796.000 1818.290 800.000 ;
    END
  END eu0_instruction[40]
  PIN eu0_instruction[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1823.070 796.000 1823.350 800.000 ;
    END
  END eu0_instruction[41]
  PIN eu0_instruction[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 10.454400 ;
    PORT
      LAYER met2 ;
        RECT 1635.850 796.000 1636.130 800.000 ;
    END
  END eu0_instruction[4]
  PIN eu0_instruction[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 10.454400 ;
    PORT
      LAYER met2 ;
        RECT 1640.910 796.000 1641.190 800.000 ;
    END
  END eu0_instruction[5]
  PIN eu0_instruction[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 10.454400 ;
    PORT
      LAYER met2 ;
        RECT 1645.970 796.000 1646.250 800.000 ;
    END
  END eu0_instruction[6]
  PIN eu0_instruction[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 10.454400 ;
    PORT
      LAYER met2 ;
        RECT 1651.030 796.000 1651.310 800.000 ;
    END
  END eu0_instruction[7]
  PIN eu0_instruction[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 10.454400 ;
    PORT
      LAYER met2 ;
        RECT 1656.090 796.000 1656.370 800.000 ;
    END
  END eu0_instruction[8]
  PIN eu0_instruction[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 31.320000 ;
    PORT
      LAYER met2 ;
        RECT 1661.150 796.000 1661.430 800.000 ;
    END
  END eu0_instruction[9]
  PIN eu1_busy
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.621000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 427.080 2200.000 427.680 ;
    END
  END eu1_busy
  PIN eu1_instruction[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 429.800 2200.000 430.400 ;
    END
  END eu1_instruction[0]
  PIN eu1_instruction[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 457.000 2200.000 457.600 ;
    END
  END eu1_instruction[10]
  PIN eu1_instruction[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 459.720 2200.000 460.320 ;
    END
  END eu1_instruction[11]
  PIN eu1_instruction[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 462.440 2200.000 463.040 ;
    END
  END eu1_instruction[12]
  PIN eu1_instruction[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 465.160 2200.000 465.760 ;
    END
  END eu1_instruction[13]
  PIN eu1_instruction[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 467.880 2200.000 468.480 ;
    END
  END eu1_instruction[14]
  PIN eu1_instruction[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 470.600 2200.000 471.200 ;
    END
  END eu1_instruction[15]
  PIN eu1_instruction[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 473.320 2200.000 473.920 ;
    END
  END eu1_instruction[16]
  PIN eu1_instruction[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 476.040 2200.000 476.640 ;
    END
  END eu1_instruction[17]
  PIN eu1_instruction[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 478.760 2200.000 479.360 ;
    END
  END eu1_instruction[18]
  PIN eu1_instruction[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 481.480 2200.000 482.080 ;
    END
  END eu1_instruction[19]
  PIN eu1_instruction[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 432.520 2200.000 433.120 ;
    END
  END eu1_instruction[1]
  PIN eu1_instruction[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 484.200 2200.000 484.800 ;
    END
  END eu1_instruction[20]
  PIN eu1_instruction[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 486.920 2200.000 487.520 ;
    END
  END eu1_instruction[21]
  PIN eu1_instruction[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 489.640 2200.000 490.240 ;
    END
  END eu1_instruction[22]
  PIN eu1_instruction[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 492.360 2200.000 492.960 ;
    END
  END eu1_instruction[23]
  PIN eu1_instruction[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 495.080 2200.000 495.680 ;
    END
  END eu1_instruction[24]
  PIN eu1_instruction[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 497.800 2200.000 498.400 ;
    END
  END eu1_instruction[25]
  PIN eu1_instruction[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 500.520 2200.000 501.120 ;
    END
  END eu1_instruction[26]
  PIN eu1_instruction[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 503.240 2200.000 503.840 ;
    END
  END eu1_instruction[27]
  PIN eu1_instruction[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 505.960 2200.000 506.560 ;
    END
  END eu1_instruction[28]
  PIN eu1_instruction[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 508.680 2200.000 509.280 ;
    END
  END eu1_instruction[29]
  PIN eu1_instruction[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 435.240 2200.000 435.840 ;
    END
  END eu1_instruction[2]
  PIN eu1_instruction[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 511.400 2200.000 512.000 ;
    END
  END eu1_instruction[30]
  PIN eu1_instruction[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 514.120 2200.000 514.720 ;
    END
  END eu1_instruction[31]
  PIN eu1_instruction[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 516.840 2200.000 517.440 ;
    END
  END eu1_instruction[32]
  PIN eu1_instruction[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 519.560 2200.000 520.160 ;
    END
  END eu1_instruction[33]
  PIN eu1_instruction[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 522.280 2200.000 522.880 ;
    END
  END eu1_instruction[34]
  PIN eu1_instruction[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 525.000 2200.000 525.600 ;
    END
  END eu1_instruction[35]
  PIN eu1_instruction[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 527.720 2200.000 528.320 ;
    END
  END eu1_instruction[36]
  PIN eu1_instruction[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 530.440 2200.000 531.040 ;
    END
  END eu1_instruction[37]
  PIN eu1_instruction[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 533.160 2200.000 533.760 ;
    END
  END eu1_instruction[38]
  PIN eu1_instruction[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 535.880 2200.000 536.480 ;
    END
  END eu1_instruction[39]
  PIN eu1_instruction[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 437.960 2200.000 438.560 ;
    END
  END eu1_instruction[3]
  PIN eu1_instruction[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 538.600 2200.000 539.200 ;
    END
  END eu1_instruction[40]
  PIN eu1_instruction[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 541.320 2200.000 541.920 ;
    END
  END eu1_instruction[41]
  PIN eu1_instruction[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 440.680 2200.000 441.280 ;
    END
  END eu1_instruction[4]
  PIN eu1_instruction[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 443.400 2200.000 444.000 ;
    END
  END eu1_instruction[5]
  PIN eu1_instruction[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 446.120 2200.000 446.720 ;
    END
  END eu1_instruction[6]
  PIN eu1_instruction[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 448.840 2200.000 449.440 ;
    END
  END eu1_instruction[7]
  PIN eu1_instruction[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 451.560 2200.000 452.160 ;
    END
  END eu1_instruction[8]
  PIN eu1_instruction[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 454.280 2200.000 454.880 ;
    END
  END eu1_instruction[9]
  PIN eu2_busy
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.621000 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 421.640 4.000 422.240 ;
    END
  END eu2_busy
  PIN eu2_instruction[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 424.360 4.000 424.960 ;
    END
  END eu2_instruction[0]
  PIN eu2_instruction[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 451.560 4.000 452.160 ;
    END
  END eu2_instruction[10]
  PIN eu2_instruction[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 454.280 4.000 454.880 ;
    END
  END eu2_instruction[11]
  PIN eu2_instruction[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 457.000 4.000 457.600 ;
    END
  END eu2_instruction[12]
  PIN eu2_instruction[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 459.720 4.000 460.320 ;
    END
  END eu2_instruction[13]
  PIN eu2_instruction[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 462.440 4.000 463.040 ;
    END
  END eu2_instruction[14]
  PIN eu2_instruction[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 465.160 4.000 465.760 ;
    END
  END eu2_instruction[15]
  PIN eu2_instruction[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 467.880 4.000 468.480 ;
    END
  END eu2_instruction[16]
  PIN eu2_instruction[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 470.600 4.000 471.200 ;
    END
  END eu2_instruction[17]
  PIN eu2_instruction[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 473.320 4.000 473.920 ;
    END
  END eu2_instruction[18]
  PIN eu2_instruction[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 476.040 4.000 476.640 ;
    END
  END eu2_instruction[19]
  PIN eu2_instruction[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 427.080 4.000 427.680 ;
    END
  END eu2_instruction[1]
  PIN eu2_instruction[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 478.760 4.000 479.360 ;
    END
  END eu2_instruction[20]
  PIN eu2_instruction[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 481.480 4.000 482.080 ;
    END
  END eu2_instruction[21]
  PIN eu2_instruction[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 484.200 4.000 484.800 ;
    END
  END eu2_instruction[22]
  PIN eu2_instruction[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 486.920 4.000 487.520 ;
    END
  END eu2_instruction[23]
  PIN eu2_instruction[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 489.640 4.000 490.240 ;
    END
  END eu2_instruction[24]
  PIN eu2_instruction[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 492.360 4.000 492.960 ;
    END
  END eu2_instruction[25]
  PIN eu2_instruction[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 495.080 4.000 495.680 ;
    END
  END eu2_instruction[26]
  PIN eu2_instruction[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 497.800 4.000 498.400 ;
    END
  END eu2_instruction[27]
  PIN eu2_instruction[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 500.520 4.000 501.120 ;
    END
  END eu2_instruction[28]
  PIN eu2_instruction[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 503.240 4.000 503.840 ;
    END
  END eu2_instruction[29]
  PIN eu2_instruction[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 429.800 4.000 430.400 ;
    END
  END eu2_instruction[2]
  PIN eu2_instruction[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 505.960 4.000 506.560 ;
    END
  END eu2_instruction[30]
  PIN eu2_instruction[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 508.680 4.000 509.280 ;
    END
  END eu2_instruction[31]
  PIN eu2_instruction[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 511.400 4.000 512.000 ;
    END
  END eu2_instruction[32]
  PIN eu2_instruction[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 514.120 4.000 514.720 ;
    END
  END eu2_instruction[33]
  PIN eu2_instruction[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 516.840 4.000 517.440 ;
    END
  END eu2_instruction[34]
  PIN eu2_instruction[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 519.560 4.000 520.160 ;
    END
  END eu2_instruction[35]
  PIN eu2_instruction[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 522.280 4.000 522.880 ;
    END
  END eu2_instruction[36]
  PIN eu2_instruction[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 525.000 4.000 525.600 ;
    END
  END eu2_instruction[37]
  PIN eu2_instruction[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 527.720 4.000 528.320 ;
    END
  END eu2_instruction[38]
  PIN eu2_instruction[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 530.440 4.000 531.040 ;
    END
  END eu2_instruction[39]
  PIN eu2_instruction[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 432.520 4.000 433.120 ;
    END
  END eu2_instruction[3]
  PIN eu2_instruction[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 533.160 4.000 533.760 ;
    END
  END eu2_instruction[40]
  PIN eu2_instruction[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 535.880 4.000 536.480 ;
    END
  END eu2_instruction[41]
  PIN eu2_instruction[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.240 4.000 435.840 ;
    END
  END eu2_instruction[4]
  PIN eu2_instruction[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 437.960 4.000 438.560 ;
    END
  END eu2_instruction[5]
  PIN eu2_instruction[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 440.680 4.000 441.280 ;
    END
  END eu2_instruction[6]
  PIN eu2_instruction[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 443.400 4.000 444.000 ;
    END
  END eu2_instruction[7]
  PIN eu2_instruction[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 446.120 4.000 446.720 ;
    END
  END eu2_instruction[8]
  PIN eu2_instruction[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 448.840 4.000 449.440 ;
    END
  END eu2_instruction[9]
  PIN int_return0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 2157.030 796.000 2157.310 800.000 ;
    END
  END int_return0
  PIN int_return1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 720.840 2200.000 721.440 ;
    END
  END int_return1
  PIN int_return2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 715.400 4.000 716.000 ;
    END
  END int_return2
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 1160.670 0.000 1160.950 4.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.984500 ;
    PORT
      LAYER met2 ;
        RECT 1248.070 0.000 1248.350 4.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.858500 ;
    PORT
      LAYER met2 ;
        RECT 1256.810 0.000 1257.090 4.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.106000 ;
    PORT
      LAYER met2 ;
        RECT 1265.550 0.000 1265.830 4.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.858500 ;
    PORT
      LAYER met2 ;
        RECT 1274.290 0.000 1274.570 4.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.858500 ;
    PORT
      LAYER met2 ;
        RECT 1283.030 0.000 1283.310 4.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.106000 ;
    PORT
      LAYER met2 ;
        RECT 1291.770 0.000 1292.050 4.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.106000 ;
    PORT
      LAYER met2 ;
        RECT 1300.510 0.000 1300.790 4.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.358000 ;
    PORT
      LAYER met2 ;
        RECT 1309.250 0.000 1309.530 4.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.601000 ;
    PORT
      LAYER met2 ;
        RECT 1317.990 0.000 1318.270 4.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1326.730 0.000 1327.010 4.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1169.410 0.000 1169.690 4.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1335.470 0.000 1335.750 4.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1344.210 0.000 1344.490 4.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1352.950 0.000 1353.230 4.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1361.690 0.000 1361.970 4.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1370.430 0.000 1370.710 4.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1379.170 0.000 1379.450 4.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116000 ;
    PORT
      LAYER met2 ;
        RECT 1387.910 0.000 1388.190 4.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1396.650 0.000 1396.930 4.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1405.390 0.000 1405.670 4.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 1414.130 0.000 1414.410 4.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 1178.150 0.000 1178.430 4.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 1422.870 0.000 1423.150 4.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.621000 ;
    PORT
      LAYER met2 ;
        RECT 1431.610 0.000 1431.890 4.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1440.350 0.000 1440.630 4.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 1449.090 0.000 1449.370 4.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 1457.830 0.000 1458.110 4.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 1466.570 0.000 1466.850 4.000 ;
    END
  END io_in[35]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.106000 ;
    PORT
      LAYER met2 ;
        RECT 1186.890 0.000 1187.170 4.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.106000 ;
    PORT
      LAYER met2 ;
        RECT 1195.630 0.000 1195.910 4.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.106000 ;
    PORT
      LAYER met2 ;
        RECT 1204.370 0.000 1204.650 4.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.106000 ;
    PORT
      LAYER met2 ;
        RECT 1213.110 0.000 1213.390 4.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.984500 ;
    PORT
      LAYER met2 ;
        RECT 1221.850 0.000 1222.130 4.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.984500 ;
    PORT
      LAYER met2 ;
        RECT 1230.590 0.000 1230.870 4.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.984500 ;
    PORT
      LAYER met2 ;
        RECT 1239.330 0.000 1239.610 4.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.484000 ;
    PORT
      LAYER met2 ;
        RECT 1475.310 0.000 1475.590 4.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1562.710 0.000 1562.990 4.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1571.450 0.000 1571.730 4.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1580.190 0.000 1580.470 4.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1588.930 0.000 1589.210 4.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1597.670 0.000 1597.950 4.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1606.410 0.000 1606.690 4.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1615.150 0.000 1615.430 4.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1623.890 0.000 1624.170 4.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 14.849999 ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1632.630 0.000 1632.910 4.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1641.370 0.000 1641.650 4.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1484.050 0.000 1484.330 4.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1650.110 0.000 1650.390 4.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1658.850 0.000 1659.130 4.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1667.590 0.000 1667.870 4.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1676.330 0.000 1676.610 4.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1685.070 0.000 1685.350 4.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1693.810 0.000 1694.090 4.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1702.550 0.000 1702.830 4.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1711.290 0.000 1711.570 4.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1720.030 0.000 1720.310 4.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1728.770 0.000 1729.050 4.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.484000 ;
    PORT
      LAYER met2 ;
        RECT 1492.790 0.000 1493.070 4.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1737.510 0.000 1737.790 4.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1746.250 0.000 1746.530 4.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1754.990 0.000 1755.270 4.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1763.730 0.000 1764.010 4.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1772.470 0.000 1772.750 4.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met2 ;
        RECT 1781.210 0.000 1781.490 4.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1501.530 0.000 1501.810 4.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1510.270 0.000 1510.550 4.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1519.010 0.000 1519.290 4.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1527.750 0.000 1528.030 4.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1536.490 0.000 1536.770 4.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1545.230 0.000 1545.510 4.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1553.970 0.000 1554.250 4.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1789.950 0.000 1790.230 4.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1877.350 0.000 1877.630 4.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1886.090 0.000 1886.370 4.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1894.830 0.000 1895.110 4.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1903.570 0.000 1903.850 4.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1912.310 0.000 1912.590 4.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1921.050 0.000 1921.330 4.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1929.790 0.000 1930.070 4.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1938.530 0.000 1938.810 4.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1947.270 0.000 1947.550 4.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1956.010 0.000 1956.290 4.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1798.690 0.000 1798.970 4.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1964.750 0.000 1965.030 4.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1973.490 0.000 1973.770 4.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 1982.230 0.000 1982.510 4.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 1990.970 0.000 1991.250 4.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.715500 ;
    PORT
      LAYER met2 ;
        RECT 1999.710 0.000 1999.990 4.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 2008.450 0.000 2008.730 4.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2017.190 0.000 2017.470 4.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 2025.930 0.000 2026.210 4.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 2034.670 0.000 2034.950 4.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2043.410 0.000 2043.690 4.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1807.430 0.000 1807.710 4.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 2052.150 0.000 2052.430 4.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 4.803300 ;
    PORT
      LAYER met2 ;
        RECT 2060.890 0.000 2061.170 4.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 2.195100 ;
    PORT
      LAYER met2 ;
        RECT 2069.630 0.000 2069.910 4.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 6.107400 ;
    PORT
      LAYER met2 ;
        RECT 2078.370 0.000 2078.650 4.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.621000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 2087.110 0.000 2087.390 4.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.621000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 2095.850 0.000 2096.130 4.000 ;
    END
  END io_out[35]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1816.170 0.000 1816.450 4.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1824.910 0.000 1825.190 4.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1833.650 0.000 1833.930 4.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1842.390 0.000 1842.670 4.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1851.130 0.000 1851.410 4.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1859.870 0.000 1860.150 4.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 1868.610 0.000 1868.890 4.000 ;
    END
  END io_out[9]
  PIN is_load0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.980000 ;
    PORT
      LAYER met2 ;
        RECT 1438.510 796.000 1438.790 800.000 ;
    END
  END is_load0
  PIN is_load1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.489500 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 334.600 2200.000 335.200 ;
    END
  END is_load1
  PIN is_load2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.227500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.160 4.000 329.760 ;
    END
  END is_load2
  PIN is_store0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.858500 ;
    PORT
      LAYER met2 ;
        RECT 1443.570 796.000 1443.850 800.000 ;
    END
  END is_store0
  PIN is_store1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.363500 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 337.320 2200.000 337.920 ;
    END
  END is_store1
  PIN is_store2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.980000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 331.880 4.000 332.480 ;
    END
  END is_store2
  PIN loadstore_address0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 2.173500 ;
    PORT
      LAYER met2 ;
        RECT 1276.590 796.000 1276.870 800.000 ;
    END
  END loadstore_address0[0]
  PIN loadstore_address0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met2 ;
        RECT 1327.190 796.000 1327.470 800.000 ;
    END
  END loadstore_address0[10]
  PIN loadstore_address0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1332.250 796.000 1332.530 800.000 ;
    END
  END loadstore_address0[11]
  PIN loadstore_address0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 2.173500 ;
    PORT
      LAYER met2 ;
        RECT 1337.310 796.000 1337.590 800.000 ;
    END
  END loadstore_address0[12]
  PIN loadstore_address0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 2.173500 ;
    PORT
      LAYER met2 ;
        RECT 1342.370 796.000 1342.650 800.000 ;
    END
  END loadstore_address0[13]
  PIN loadstore_address0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met2 ;
        RECT 1347.430 796.000 1347.710 800.000 ;
    END
  END loadstore_address0[14]
  PIN loadstore_address0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1352.490 796.000 1352.770 800.000 ;
    END
  END loadstore_address0[15]
  PIN loadstore_address0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1357.550 796.000 1357.830 800.000 ;
    END
  END loadstore_address0[16]
  PIN loadstore_address0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1362.610 796.000 1362.890 800.000 ;
    END
  END loadstore_address0[17]
  PIN loadstore_address0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1367.670 796.000 1367.950 800.000 ;
    END
  END loadstore_address0[18]
  PIN loadstore_address0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met2 ;
        RECT 1372.730 796.000 1373.010 800.000 ;
    END
  END loadstore_address0[19]
  PIN loadstore_address0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 2.608200 ;
    PORT
      LAYER met2 ;
        RECT 1281.650 796.000 1281.930 800.000 ;
    END
  END loadstore_address0[1]
  PIN loadstore_address0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1377.790 796.000 1378.070 800.000 ;
    END
  END loadstore_address0[20]
  PIN loadstore_address0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met2 ;
        RECT 1382.850 796.000 1383.130 800.000 ;
    END
  END loadstore_address0[21]
  PIN loadstore_address0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met2 ;
        RECT 1387.910 796.000 1388.190 800.000 ;
    END
  END loadstore_address0[22]
  PIN loadstore_address0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1392.970 796.000 1393.250 800.000 ;
    END
  END loadstore_address0[23]
  PIN loadstore_address0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 2.608200 ;
    PORT
      LAYER met2 ;
        RECT 1398.030 796.000 1398.310 800.000 ;
    END
  END loadstore_address0[24]
  PIN loadstore_address0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1403.090 796.000 1403.370 800.000 ;
    END
  END loadstore_address0[25]
  PIN loadstore_address0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met2 ;
        RECT 1408.150 796.000 1408.430 800.000 ;
    END
  END loadstore_address0[26]
  PIN loadstore_address0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met2 ;
        RECT 1413.210 796.000 1413.490 800.000 ;
    END
  END loadstore_address0[27]
  PIN loadstore_address0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1418.270 796.000 1418.550 800.000 ;
    END
  END loadstore_address0[28]
  PIN loadstore_address0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1423.330 796.000 1423.610 800.000 ;
    END
  END loadstore_address0[29]
  PIN loadstore_address0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met2 ;
        RECT 1286.710 796.000 1286.990 800.000 ;
    END
  END loadstore_address0[2]
  PIN loadstore_address0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met2 ;
        RECT 1428.390 796.000 1428.670 800.000 ;
    END
  END loadstore_address0[30]
  PIN loadstore_address0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1433.450 796.000 1433.730 800.000 ;
    END
  END loadstore_address0[31]
  PIN loadstore_address0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met2 ;
        RECT 1291.770 796.000 1292.050 800.000 ;
    END
  END loadstore_address0[3]
  PIN loadstore_address0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1296.830 796.000 1297.110 800.000 ;
    END
  END loadstore_address0[4]
  PIN loadstore_address0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 3.042900 ;
    PORT
      LAYER met2 ;
        RECT 1301.890 796.000 1302.170 800.000 ;
    END
  END loadstore_address0[5]
  PIN loadstore_address0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 2.608200 ;
    PORT
      LAYER met2 ;
        RECT 1306.950 796.000 1307.230 800.000 ;
    END
  END loadstore_address0[6]
  PIN loadstore_address0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 5.216400 ;
    PORT
      LAYER met2 ;
        RECT 1312.010 796.000 1312.290 800.000 ;
    END
  END loadstore_address0[7]
  PIN loadstore_address0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 2.173500 ;
    PORT
      LAYER met2 ;
        RECT 1317.070 796.000 1317.350 800.000 ;
    END
  END loadstore_address0[8]
  PIN loadstore_address0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 3.042900 ;
    PORT
      LAYER met2 ;
        RECT 1322.130 796.000 1322.410 800.000 ;
    END
  END loadstore_address0[9]
  PIN loadstore_address1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 9.998099 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 247.560 2200.000 248.160 ;
    END
  END loadstore_address1[0]
  PIN loadstore_address1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 274.760 2200.000 275.360 ;
    END
  END loadstore_address1[10]
  PIN loadstore_address1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 9.998099 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 277.480 2200.000 278.080 ;
    END
  END loadstore_address1[11]
  PIN loadstore_address1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 280.200 2200.000 280.800 ;
    END
  END loadstore_address1[12]
  PIN loadstore_address1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 9.128699 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 282.920 2200.000 283.520 ;
    END
  END loadstore_address1[13]
  PIN loadstore_address1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 7.389900 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 285.640 2200.000 286.240 ;
    END
  END loadstore_address1[14]
  PIN loadstore_address1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 288.360 2200.000 288.960 ;
    END
  END loadstore_address1[15]
  PIN loadstore_address1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 9.998099 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 291.080 2200.000 291.680 ;
    END
  END loadstore_address1[16]
  PIN loadstore_address1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 9.128699 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 293.800 2200.000 294.400 ;
    END
  END loadstore_address1[17]
  PIN loadstore_address1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 9.563399 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 296.520 2200.000 297.120 ;
    END
  END loadstore_address1[18]
  PIN loadstore_address1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 299.240 2200.000 299.840 ;
    END
  END loadstore_address1[19]
  PIN loadstore_address1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 250.280 2200.000 250.880 ;
    END
  END loadstore_address1[1]
  PIN loadstore_address1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 9.563399 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 301.960 2200.000 302.560 ;
    END
  END loadstore_address1[20]
  PIN loadstore_address1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 9.998099 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 304.680 2200.000 305.280 ;
    END
  END loadstore_address1[21]
  PIN loadstore_address1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 307.400 2200.000 308.000 ;
    END
  END loadstore_address1[22]
  PIN loadstore_address1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 310.120 2200.000 310.720 ;
    END
  END loadstore_address1[23]
  PIN loadstore_address1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 9.998099 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 312.840 2200.000 313.440 ;
    END
  END loadstore_address1[24]
  PIN loadstore_address1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 8.694000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 315.560 2200.000 316.160 ;
    END
  END loadstore_address1[25]
  PIN loadstore_address1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 5.216400 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 318.280 2200.000 318.880 ;
    END
  END loadstore_address1[26]
  PIN loadstore_address1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 321.000 2200.000 321.600 ;
    END
  END loadstore_address1[27]
  PIN loadstore_address1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 323.720 2200.000 324.320 ;
    END
  END loadstore_address1[28]
  PIN loadstore_address1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 326.440 2200.000 327.040 ;
    END
  END loadstore_address1[29]
  PIN loadstore_address1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 9.998099 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 253.000 2200.000 253.600 ;
    END
  END loadstore_address1[2]
  PIN loadstore_address1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 329.160 2200.000 329.760 ;
    END
  END loadstore_address1[30]
  PIN loadstore_address1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 331.880 2200.000 332.480 ;
    END
  END loadstore_address1[31]
  PIN loadstore_address1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 255.720 2200.000 256.320 ;
    END
  END loadstore_address1[3]
  PIN loadstore_address1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 258.440 2200.000 259.040 ;
    END
  END loadstore_address1[4]
  PIN loadstore_address1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 261.160 2200.000 261.760 ;
    END
  END loadstore_address1[5]
  PIN loadstore_address1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 263.880 2200.000 264.480 ;
    END
  END loadstore_address1[6]
  PIN loadstore_address1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 9.563399 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 266.600 2200.000 267.200 ;
    END
  END loadstore_address1[7]
  PIN loadstore_address1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 269.320 2200.000 269.920 ;
    END
  END loadstore_address1[8]
  PIN loadstore_address1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 272.040 2200.000 272.640 ;
    END
  END loadstore_address1[9]
  PIN loadstore_address2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 16.518600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 242.120 4.000 242.720 ;
    END
  END loadstore_address2[0]
  PIN loadstore_address2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 14.779799 ;
    PORT
      LAYER met3 ;
        RECT 0.000 269.320 4.000 269.920 ;
    END
  END loadstore_address2[10]
  PIN loadstore_address2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 9.563399 ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.040 4.000 272.640 ;
    END
  END loadstore_address2[11]
  PIN loadstore_address2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 15.214499 ;
    PORT
      LAYER met3 ;
        RECT 0.000 274.760 4.000 275.360 ;
    END
  END loadstore_address2[12]
  PIN loadstore_address2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 2.608200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 277.480 4.000 278.080 ;
    END
  END loadstore_address2[13]
  PIN loadstore_address2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 280.200 4.000 280.800 ;
    END
  END loadstore_address2[14]
  PIN loadstore_address2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 18.692099 ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.920 4.000 283.520 ;
    END
  END loadstore_address2[15]
  PIN loadstore_address2[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 9.998099 ;
    PORT
      LAYER met3 ;
        RECT 0.000 285.640 4.000 286.240 ;
    END
  END loadstore_address2[16]
  PIN loadstore_address2[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 11.736899 ;
    PORT
      LAYER met3 ;
        RECT 0.000 288.360 4.000 288.960 ;
    END
  END loadstore_address2[17]
  PIN loadstore_address2[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 9.998099 ;
    PORT
      LAYER met3 ;
        RECT 0.000 291.080 4.000 291.680 ;
    END
  END loadstore_address2[18]
  PIN loadstore_address2[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 293.800 4.000 294.400 ;
    END
  END loadstore_address2[19]
  PIN loadstore_address2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 9.563399 ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.840 4.000 245.440 ;
    END
  END loadstore_address2[1]
  PIN loadstore_address2[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 13.475699 ;
    PORT
      LAYER met3 ;
        RECT 0.000 296.520 4.000 297.120 ;
    END
  END loadstore_address2[20]
  PIN loadstore_address2[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 5.216400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.240 4.000 299.840 ;
    END
  END loadstore_address2[21]
  PIN loadstore_address2[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 15.214499 ;
    PORT
      LAYER met3 ;
        RECT 0.000 301.960 4.000 302.560 ;
    END
  END loadstore_address2[22]
  PIN loadstore_address2[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 304.680 4.000 305.280 ;
    END
  END loadstore_address2[23]
  PIN loadstore_address2[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 19.561499 ;
    PORT
      LAYER met3 ;
        RECT 0.000 307.400 4.000 308.000 ;
    END
  END loadstore_address2[24]
  PIN loadstore_address2[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 11.736899 ;
    PORT
      LAYER met3 ;
        RECT 0.000 310.120 4.000 310.720 ;
    END
  END loadstore_address2[25]
  PIN loadstore_address2[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 9.998099 ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.840 4.000 313.440 ;
    END
  END loadstore_address2[26]
  PIN loadstore_address2[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 7.389900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 315.560 4.000 316.160 ;
    END
  END loadstore_address2[27]
  PIN loadstore_address2[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 13.475699 ;
    PORT
      LAYER met3 ;
        RECT 0.000 318.280 4.000 318.880 ;
    END
  END loadstore_address2[28]
  PIN loadstore_address2[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 321.000 4.000 321.600 ;
    END
  END loadstore_address2[29]
  PIN loadstore_address2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 9.998099 ;
    PORT
      LAYER met3 ;
        RECT 0.000 247.560 4.000 248.160 ;
    END
  END loadstore_address2[2]
  PIN loadstore_address2[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 10.432799 ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.720 4.000 324.320 ;
    END
  END loadstore_address2[30]
  PIN loadstore_address2[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 326.440 4.000 327.040 ;
    END
  END loadstore_address2[31]
  PIN loadstore_address2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 250.280 4.000 250.880 ;
    END
  END loadstore_address2[3]
  PIN loadstore_address2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 9.128699 ;
    PORT
      LAYER met3 ;
        RECT 0.000 253.000 4.000 253.600 ;
    END
  END loadstore_address2[4]
  PIN loadstore_address2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.720 4.000 256.320 ;
    END
  END loadstore_address2[5]
  PIN loadstore_address2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 14.345099 ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END loadstore_address2[6]
  PIN loadstore_address2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 15.214499 ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.160 4.000 261.760 ;
    END
  END loadstore_address2[7]
  PIN loadstore_address2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 9.998099 ;
    PORT
      LAYER met3 ;
        RECT 0.000 263.880 4.000 264.480 ;
    END
  END loadstore_address2[8]
  PIN loadstore_address2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 9.998099 ;
    PORT
      LAYER met3 ;
        RECT 0.000 266.600 4.000 267.200 ;
    END
  END loadstore_address2[9]
  PIN loadstore_size0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met2 ;
        RECT 1453.690 796.000 1453.970 800.000 ;
    END
  END loadstore_size0[0]
  PIN loadstore_size0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1458.750 796.000 1459.030 800.000 ;
    END
  END loadstore_size0[1]
  PIN loadstore_size1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 342.760 2200.000 343.360 ;
    END
  END loadstore_size1[0]
  PIN loadstore_size1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 345.480 2200.000 346.080 ;
    END
  END loadstore_size1[1]
  PIN loadstore_size2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 337.320 4.000 337.920 ;
    END
  END loadstore_size2[0]
  PIN loadstore_size2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.040 4.000 340.640 ;
    END
  END loadstore_size2[1]
  PIN new_PC0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met2 ;
        RECT 1468.870 796.000 1469.150 800.000 ;
    END
  END new_PC0[0]
  PIN new_PC0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1519.470 796.000 1519.750 800.000 ;
    END
  END new_PC0[10]
  PIN new_PC0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1524.530 796.000 1524.810 800.000 ;
    END
  END new_PC0[11]
  PIN new_PC0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1529.590 796.000 1529.870 800.000 ;
    END
  END new_PC0[12]
  PIN new_PC0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 1534.650 796.000 1534.930 800.000 ;
    END
  END new_PC0[13]
  PIN new_PC0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met2 ;
        RECT 1539.710 796.000 1539.990 800.000 ;
    END
  END new_PC0[14]
  PIN new_PC0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met2 ;
        RECT 1544.770 796.000 1545.050 800.000 ;
    END
  END new_PC0[15]
  PIN new_PC0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 1549.830 796.000 1550.110 800.000 ;
    END
  END new_PC0[16]
  PIN new_PC0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1554.890 796.000 1555.170 800.000 ;
    END
  END new_PC0[17]
  PIN new_PC0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met2 ;
        RECT 1559.950 796.000 1560.230 800.000 ;
    END
  END new_PC0[18]
  PIN new_PC0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1565.010 796.000 1565.290 800.000 ;
    END
  END new_PC0[19]
  PIN new_PC0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1473.930 796.000 1474.210 800.000 ;
    END
  END new_PC0[1]
  PIN new_PC0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.152000 ;
    PORT
      LAYER met2 ;
        RECT 1570.070 796.000 1570.350 800.000 ;
    END
  END new_PC0[20]
  PIN new_PC0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1575.130 796.000 1575.410 800.000 ;
    END
  END new_PC0[21]
  PIN new_PC0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 5.216400 ;
    PORT
      LAYER met2 ;
        RECT 1580.190 796.000 1580.470 800.000 ;
    END
  END new_PC0[22]
  PIN new_PC0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met2 ;
        RECT 1585.250 796.000 1585.530 800.000 ;
    END
  END new_PC0[23]
  PIN new_PC0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met2 ;
        RECT 1590.310 796.000 1590.590 800.000 ;
    END
  END new_PC0[24]
  PIN new_PC0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 3.912300 ;
    PORT
      LAYER met2 ;
        RECT 1595.370 796.000 1595.650 800.000 ;
    END
  END new_PC0[25]
  PIN new_PC0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 3.912300 ;
    PORT
      LAYER met2 ;
        RECT 1600.430 796.000 1600.710 800.000 ;
    END
  END new_PC0[26]
  PIN new_PC0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met2 ;
        RECT 1605.490 796.000 1605.770 800.000 ;
    END
  END new_PC0[27]
  PIN new_PC0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 3.477600 ;
    PORT
      LAYER met2 ;
        RECT 1478.990 796.000 1479.270 800.000 ;
    END
  END new_PC0[2]
  PIN new_PC0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1484.050 796.000 1484.330 800.000 ;
    END
  END new_PC0[3]
  PIN new_PC0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 1489.110 796.000 1489.390 800.000 ;
    END
  END new_PC0[4]
  PIN new_PC0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met2 ;
        RECT 1494.170 796.000 1494.450 800.000 ;
    END
  END new_PC0[5]
  PIN new_PC0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.152000 ;
    PORT
      LAYER met2 ;
        RECT 1499.230 796.000 1499.510 800.000 ;
    END
  END new_PC0[6]
  PIN new_PC0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1504.290 796.000 1504.570 800.000 ;
    END
  END new_PC0[7]
  PIN new_PC0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 2.608200 ;
    PORT
      LAYER met2 ;
        RECT 1509.350 796.000 1509.630 800.000 ;
    END
  END new_PC0[8]
  PIN new_PC0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 2.173500 ;
    PORT
      LAYER met2 ;
        RECT 1514.410 796.000 1514.690 800.000 ;
    END
  END new_PC0[9]
  PIN new_PC1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 350.920 2200.000 351.520 ;
    END
  END new_PC1[0]
  PIN new_PC1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 378.120 2200.000 378.720 ;
    END
  END new_PC1[10]
  PIN new_PC1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 20.430899 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 380.840 2200.000 381.440 ;
    END
  END new_PC1[11]
  PIN new_PC1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 383.560 2200.000 384.160 ;
    END
  END new_PC1[12]
  PIN new_PC1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 386.280 2200.000 386.880 ;
    END
  END new_PC1[13]
  PIN new_PC1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 389.000 2200.000 389.600 ;
    END
  END new_PC1[14]
  PIN new_PC1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 391.720 2200.000 392.320 ;
    END
  END new_PC1[15]
  PIN new_PC1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 9.998099 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 394.440 2200.000 395.040 ;
    END
  END new_PC1[16]
  PIN new_PC1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 9.998099 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 397.160 2200.000 397.760 ;
    END
  END new_PC1[17]
  PIN new_PC1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 399.880 2200.000 400.480 ;
    END
  END new_PC1[18]
  PIN new_PC1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 402.600 2200.000 403.200 ;
    END
  END new_PC1[19]
  PIN new_PC1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 9.998099 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 353.640 2200.000 354.240 ;
    END
  END new_PC1[1]
  PIN new_PC1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 405.320 2200.000 405.920 ;
    END
  END new_PC1[20]
  PIN new_PC1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 408.040 2200.000 408.640 ;
    END
  END new_PC1[21]
  PIN new_PC1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 3.477600 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 410.760 2200.000 411.360 ;
    END
  END new_PC1[22]
  PIN new_PC1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 2.173500 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 413.480 2200.000 414.080 ;
    END
  END new_PC1[23]
  PIN new_PC1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 30.863699 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 416.200 2200.000 416.800 ;
    END
  END new_PC1[24]
  PIN new_PC1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 418.920 2200.000 419.520 ;
    END
  END new_PC1[25]
  PIN new_PC1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 20.430899 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 421.640 2200.000 422.240 ;
    END
  END new_PC1[26]
  PIN new_PC1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 424.360 2200.000 424.960 ;
    END
  END new_PC1[27]
  PIN new_PC1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 3.912300 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 356.360 2200.000 356.960 ;
    END
  END new_PC1[2]
  PIN new_PC1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.304000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 359.080 2200.000 359.680 ;
    END
  END new_PC1[3]
  PIN new_PC1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 25.647299 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 361.800 2200.000 362.400 ;
    END
  END new_PC1[4]
  PIN new_PC1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 364.520 2200.000 365.120 ;
    END
  END new_PC1[5]
  PIN new_PC1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 367.240 2200.000 367.840 ;
    END
  END new_PC1[6]
  PIN new_PC1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 369.960 2200.000 370.560 ;
    END
  END new_PC1[7]
  PIN new_PC1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 9.998099 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 372.680 2200.000 373.280 ;
    END
  END new_PC1[8]
  PIN new_PC1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 375.400 2200.000 376.000 ;
    END
  END new_PC1[9]
  PIN new_PC2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 345.480 4.000 346.080 ;
    END
  END new_PC2[0]
  PIN new_PC2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 372.680 4.000 373.280 ;
    END
  END new_PC2[10]
  PIN new_PC2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 375.400 4.000 376.000 ;
    END
  END new_PC2[11]
  PIN new_PC2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 378.120 4.000 378.720 ;
    END
  END new_PC2[12]
  PIN new_PC2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.840 4.000 381.440 ;
    END
  END new_PC2[13]
  PIN new_PC2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 383.560 4.000 384.160 ;
    END
  END new_PC2[14]
  PIN new_PC2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 386.280 4.000 386.880 ;
    END
  END new_PC2[15]
  PIN new_PC2[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 389.000 4.000 389.600 ;
    END
  END new_PC2[16]
  PIN new_PC2[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.720 4.000 392.320 ;
    END
  END new_PC2[17]
  PIN new_PC2[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 394.440 4.000 395.040 ;
    END
  END new_PC2[18]
  PIN new_PC2[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.160 4.000 397.760 ;
    END
  END new_PC2[19]
  PIN new_PC2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 348.200 4.000 348.800 ;
    END
  END new_PC2[1]
  PIN new_PC2[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 399.880 4.000 400.480 ;
    END
  END new_PC2[20]
  PIN new_PC2[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 402.600 4.000 403.200 ;
    END
  END new_PC2[21]
  PIN new_PC2[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 405.320 4.000 405.920 ;
    END
  END new_PC2[22]
  PIN new_PC2[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 0.000 408.040 4.000 408.640 ;
    END
  END new_PC2[23]
  PIN new_PC2[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 410.760 4.000 411.360 ;
    END
  END new_PC2[24]
  PIN new_PC2[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 0.000 413.480 4.000 414.080 ;
    END
  END new_PC2[25]
  PIN new_PC2[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 416.200 4.000 416.800 ;
    END
  END new_PC2[26]
  PIN new_PC2[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 418.920 4.000 419.520 ;
    END
  END new_PC2[27]
  PIN new_PC2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.920 4.000 351.520 ;
    END
  END new_PC2[2]
  PIN new_PC2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 353.640 4.000 354.240 ;
    END
  END new_PC2[3]
  PIN new_PC2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 356.360 4.000 356.960 ;
    END
  END new_PC2[4]
  PIN new_PC2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 359.080 4.000 359.680 ;
    END
  END new_PC2[5]
  PIN new_PC2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 361.800 4.000 362.400 ;
    END
  END new_PC2[6]
  PIN new_PC2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 364.520 4.000 365.120 ;
    END
  END new_PC2[7]
  PIN new_PC2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 367.240 4.000 367.840 ;
    END
  END new_PC2[8]
  PIN new_PC2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 369.960 4.000 370.560 ;
    END
  END new_PC2[9]
  PIN pred_idx0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.630000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1241.170 796.000 1241.450 800.000 ;
    END
  END pred_idx0[0]
  PIN pred_idx0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.630000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1246.230 796.000 1246.510 800.000 ;
    END
  END pred_idx0[1]
  PIN pred_idx0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 1251.290 796.000 1251.570 800.000 ;
    END
  END pred_idx0[2]
  PIN pred_idx1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.630000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 228.520 2200.000 229.120 ;
    END
  END pred_idx1[0]
  PIN pred_idx1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.630000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 231.240 2200.000 231.840 ;
    END
  END pred_idx1[1]
  PIN pred_idx1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 233.960 2200.000 234.560 ;
    END
  END pred_idx1[2]
  PIN pred_idx2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.696000 ;
    ANTENNADIFFAREA 5.216400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.080 4.000 223.680 ;
    END
  END pred_idx2[0]
  PIN pred_idx2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.696000 ;
    ANTENNADIFFAREA 9.998099 ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.800 4.000 226.400 ;
    END
  END pred_idx2[1]
  PIN pred_idx2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 228.520 4.000 229.120 ;
    END
  END pred_idx2[2]
  PIN pred_val0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.962500 ;
    PORT
      LAYER met2 ;
        RECT 2151.970 796.000 2152.250 800.000 ;
    END
  END pred_val0
  PIN pred_val1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.962500 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 718.120 2200.000 718.720 ;
    END
  END pred_val1
  PIN pred_val2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.962500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 712.680 4.000 713.280 ;
    END
  END pred_val2
  PIN reg1_idx0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 978.050 796.000 978.330 800.000 ;
    END
  END reg1_idx0[0]
  PIN reg1_idx0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.148500 ;
    PORT
      LAYER met2 ;
        RECT 983.110 796.000 983.390 800.000 ;
    END
  END reg1_idx0[1]
  PIN reg1_idx0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 988.170 796.000 988.450 800.000 ;
    END
  END reg1_idx0[2]
  PIN reg1_idx0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.822000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 993.230 796.000 993.510 800.000 ;
    END
  END reg1_idx0[3]
  PIN reg1_idx0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.980000 ;
    PORT
      LAYER met2 ;
        RECT 998.290 796.000 998.570 800.000 ;
    END
  END reg1_idx0[4]
  PIN reg1_idx0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.812000 ;
    PORT
      LAYER met2 ;
        RECT 1003.350 796.000 1003.630 800.000 ;
    END
  END reg1_idx0[5]
  PIN reg1_idx1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.674000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 87.080 2200.000 87.680 ;
    END
  END reg1_idx1[0]
  PIN reg1_idx1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 89.800 2200.000 90.400 ;
    END
  END reg1_idx1[1]
  PIN reg1_idx1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 92.520 2200.000 93.120 ;
    END
  END reg1_idx1[2]
  PIN reg1_idx1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.684000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 95.240 2200.000 95.840 ;
    END
  END reg1_idx1[3]
  PIN reg1_idx1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 97.960 2200.000 98.560 ;
    END
  END reg1_idx1[4]
  PIN reg1_idx1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.327000 ;
    ANTENNADIFFAREA 3.477600 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 100.680 2200.000 101.280 ;
    END
  END reg1_idx1[5]
  PIN reg1_idx2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.980000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END reg1_idx2[0]
  PIN reg1_idx2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.360 4.000 84.960 ;
    END
  END reg1_idx2[1]
  PIN reg1_idx2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.080 4.000 87.680 ;
    END
  END reg1_idx2[2]
  PIN reg1_idx2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.822000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 4.000 90.400 ;
    END
  END reg1_idx2[3]
  PIN reg1_idx2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.475000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.520 4.000 93.120 ;
    END
  END reg1_idx2[4]
  PIN reg1_idx2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END reg1_idx2[5]
  PIN reg1_val0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1828.130 796.000 1828.410 800.000 ;
    END
  END reg1_val0[0]
  PIN reg1_val0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1878.730 796.000 1879.010 800.000 ;
    END
  END reg1_val0[10]
  PIN reg1_val0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1883.790 796.000 1884.070 800.000 ;
    END
  END reg1_val0[11]
  PIN reg1_val0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1888.850 796.000 1889.130 800.000 ;
    END
  END reg1_val0[12]
  PIN reg1_val0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1893.910 796.000 1894.190 800.000 ;
    END
  END reg1_val0[13]
  PIN reg1_val0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1898.970 796.000 1899.250 800.000 ;
    END
  END reg1_val0[14]
  PIN reg1_val0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1904.030 796.000 1904.310 800.000 ;
    END
  END reg1_val0[15]
  PIN reg1_val0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1909.090 796.000 1909.370 800.000 ;
    END
  END reg1_val0[16]
  PIN reg1_val0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1914.150 796.000 1914.430 800.000 ;
    END
  END reg1_val0[17]
  PIN reg1_val0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1919.210 796.000 1919.490 800.000 ;
    END
  END reg1_val0[18]
  PIN reg1_val0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1924.270 796.000 1924.550 800.000 ;
    END
  END reg1_val0[19]
  PIN reg1_val0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1833.190 796.000 1833.470 800.000 ;
    END
  END reg1_val0[1]
  PIN reg1_val0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1929.330 796.000 1929.610 800.000 ;
    END
  END reg1_val0[20]
  PIN reg1_val0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1934.390 796.000 1934.670 800.000 ;
    END
  END reg1_val0[21]
  PIN reg1_val0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1939.450 796.000 1939.730 800.000 ;
    END
  END reg1_val0[22]
  PIN reg1_val0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1944.510 796.000 1944.790 800.000 ;
    END
  END reg1_val0[23]
  PIN reg1_val0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1949.570 796.000 1949.850 800.000 ;
    END
  END reg1_val0[24]
  PIN reg1_val0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1954.630 796.000 1954.910 800.000 ;
    END
  END reg1_val0[25]
  PIN reg1_val0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1959.690 796.000 1959.970 800.000 ;
    END
  END reg1_val0[26]
  PIN reg1_val0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1964.750 796.000 1965.030 800.000 ;
    END
  END reg1_val0[27]
  PIN reg1_val0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1969.810 796.000 1970.090 800.000 ;
    END
  END reg1_val0[28]
  PIN reg1_val0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1974.870 796.000 1975.150 800.000 ;
    END
  END reg1_val0[29]
  PIN reg1_val0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1838.250 796.000 1838.530 800.000 ;
    END
  END reg1_val0[2]
  PIN reg1_val0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1979.930 796.000 1980.210 800.000 ;
    END
  END reg1_val0[30]
  PIN reg1_val0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1984.990 796.000 1985.270 800.000 ;
    END
  END reg1_val0[31]
  PIN reg1_val0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1843.310 796.000 1843.590 800.000 ;
    END
  END reg1_val0[3]
  PIN reg1_val0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1848.370 796.000 1848.650 800.000 ;
    END
  END reg1_val0[4]
  PIN reg1_val0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1853.430 796.000 1853.710 800.000 ;
    END
  END reg1_val0[5]
  PIN reg1_val0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1858.490 796.000 1858.770 800.000 ;
    END
  END reg1_val0[6]
  PIN reg1_val0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1863.550 796.000 1863.830 800.000 ;
    END
  END reg1_val0[7]
  PIN reg1_val0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1868.610 796.000 1868.890 800.000 ;
    END
  END reg1_val0[8]
  PIN reg1_val0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1873.670 796.000 1873.950 800.000 ;
    END
  END reg1_val0[9]
  PIN reg1_val1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 544.040 2200.000 544.640 ;
    END
  END reg1_val1[0]
  PIN reg1_val1[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 571.240 2200.000 571.840 ;
    END
  END reg1_val1[10]
  PIN reg1_val1[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 573.960 2200.000 574.560 ;
    END
  END reg1_val1[11]
  PIN reg1_val1[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 576.680 2200.000 577.280 ;
    END
  END reg1_val1[12]
  PIN reg1_val1[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 579.400 2200.000 580.000 ;
    END
  END reg1_val1[13]
  PIN reg1_val1[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 582.120 2200.000 582.720 ;
    END
  END reg1_val1[14]
  PIN reg1_val1[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 584.840 2200.000 585.440 ;
    END
  END reg1_val1[15]
  PIN reg1_val1[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 587.560 2200.000 588.160 ;
    END
  END reg1_val1[16]
  PIN reg1_val1[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 590.280 2200.000 590.880 ;
    END
  END reg1_val1[17]
  PIN reg1_val1[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 593.000 2200.000 593.600 ;
    END
  END reg1_val1[18]
  PIN reg1_val1[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 595.720 2200.000 596.320 ;
    END
  END reg1_val1[19]
  PIN reg1_val1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 546.760 2200.000 547.360 ;
    END
  END reg1_val1[1]
  PIN reg1_val1[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 598.440 2200.000 599.040 ;
    END
  END reg1_val1[20]
  PIN reg1_val1[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 601.160 2200.000 601.760 ;
    END
  END reg1_val1[21]
  PIN reg1_val1[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 603.880 2200.000 604.480 ;
    END
  END reg1_val1[22]
  PIN reg1_val1[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 606.600 2200.000 607.200 ;
    END
  END reg1_val1[23]
  PIN reg1_val1[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 609.320 2200.000 609.920 ;
    END
  END reg1_val1[24]
  PIN reg1_val1[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 612.040 2200.000 612.640 ;
    END
  END reg1_val1[25]
  PIN reg1_val1[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 614.760 2200.000 615.360 ;
    END
  END reg1_val1[26]
  PIN reg1_val1[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 617.480 2200.000 618.080 ;
    END
  END reg1_val1[27]
  PIN reg1_val1[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 620.200 2200.000 620.800 ;
    END
  END reg1_val1[28]
  PIN reg1_val1[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 622.920 2200.000 623.520 ;
    END
  END reg1_val1[29]
  PIN reg1_val1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 549.480 2200.000 550.080 ;
    END
  END reg1_val1[2]
  PIN reg1_val1[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 625.640 2200.000 626.240 ;
    END
  END reg1_val1[30]
  PIN reg1_val1[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 628.360 2200.000 628.960 ;
    END
  END reg1_val1[31]
  PIN reg1_val1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 552.200 2200.000 552.800 ;
    END
  END reg1_val1[3]
  PIN reg1_val1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 554.920 2200.000 555.520 ;
    END
  END reg1_val1[4]
  PIN reg1_val1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 557.640 2200.000 558.240 ;
    END
  END reg1_val1[5]
  PIN reg1_val1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 560.360 2200.000 560.960 ;
    END
  END reg1_val1[6]
  PIN reg1_val1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 563.080 2200.000 563.680 ;
    END
  END reg1_val1[7]
  PIN reg1_val1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 565.800 2200.000 566.400 ;
    END
  END reg1_val1[8]
  PIN reg1_val1[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 568.520 2200.000 569.120 ;
    END
  END reg1_val1[9]
  PIN reg1_val2[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 538.600 4.000 539.200 ;
    END
  END reg1_val2[0]
  PIN reg1_val2[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 565.800 4.000 566.400 ;
    END
  END reg1_val2[10]
  PIN reg1_val2[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 568.520 4.000 569.120 ;
    END
  END reg1_val2[11]
  PIN reg1_val2[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 571.240 4.000 571.840 ;
    END
  END reg1_val2[12]
  PIN reg1_val2[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 573.960 4.000 574.560 ;
    END
  END reg1_val2[13]
  PIN reg1_val2[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 576.680 4.000 577.280 ;
    END
  END reg1_val2[14]
  PIN reg1_val2[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 579.400 4.000 580.000 ;
    END
  END reg1_val2[15]
  PIN reg1_val2[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 582.120 4.000 582.720 ;
    END
  END reg1_val2[16]
  PIN reg1_val2[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 584.840 4.000 585.440 ;
    END
  END reg1_val2[17]
  PIN reg1_val2[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 587.560 4.000 588.160 ;
    END
  END reg1_val2[18]
  PIN reg1_val2[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 590.280 4.000 590.880 ;
    END
  END reg1_val2[19]
  PIN reg1_val2[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 541.320 4.000 541.920 ;
    END
  END reg1_val2[1]
  PIN reg1_val2[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 593.000 4.000 593.600 ;
    END
  END reg1_val2[20]
  PIN reg1_val2[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 595.720 4.000 596.320 ;
    END
  END reg1_val2[21]
  PIN reg1_val2[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 598.440 4.000 599.040 ;
    END
  END reg1_val2[22]
  PIN reg1_val2[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 601.160 4.000 601.760 ;
    END
  END reg1_val2[23]
  PIN reg1_val2[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 603.880 4.000 604.480 ;
    END
  END reg1_val2[24]
  PIN reg1_val2[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 606.600 4.000 607.200 ;
    END
  END reg1_val2[25]
  PIN reg1_val2[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 609.320 4.000 609.920 ;
    END
  END reg1_val2[26]
  PIN reg1_val2[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 612.040 4.000 612.640 ;
    END
  END reg1_val2[27]
  PIN reg1_val2[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 614.760 4.000 615.360 ;
    END
  END reg1_val2[28]
  PIN reg1_val2[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 617.480 4.000 618.080 ;
    END
  END reg1_val2[29]
  PIN reg1_val2[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 544.040 4.000 544.640 ;
    END
  END reg1_val2[2]
  PIN reg1_val2[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 620.200 4.000 620.800 ;
    END
  END reg1_val2[30]
  PIN reg1_val2[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 622.920 4.000 623.520 ;
    END
  END reg1_val2[31]
  PIN reg1_val2[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 546.760 4.000 547.360 ;
    END
  END reg1_val2[3]
  PIN reg1_val2[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 549.480 4.000 550.080 ;
    END
  END reg1_val2[4]
  PIN reg1_val2[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 552.200 4.000 552.800 ;
    END
  END reg1_val2[5]
  PIN reg1_val2[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 554.920 4.000 555.520 ;
    END
  END reg1_val2[6]
  PIN reg1_val2[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 557.640 4.000 558.240 ;
    END
  END reg1_val2[7]
  PIN reg1_val2[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 560.360 4.000 560.960 ;
    END
  END reg1_val2[8]
  PIN reg1_val2[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 563.080 4.000 563.680 ;
    END
  END reg1_val2[9]
  PIN reg2_idx0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.822000 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met2 ;
        RECT 1008.410 796.000 1008.690 800.000 ;
    END
  END reg2_idx0[0]
  PIN reg2_idx0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 1013.470 796.000 1013.750 800.000 ;
    END
  END reg2_idx0[1]
  PIN reg2_idx0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 1018.530 796.000 1018.810 800.000 ;
    END
  END reg2_idx0[2]
  PIN reg2_idx0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.684000 ;
    PORT
      LAYER met2 ;
        RECT 1023.590 796.000 1023.870 800.000 ;
    END
  END reg2_idx0[3]
  PIN reg2_idx0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.094000 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met2 ;
        RECT 1028.650 796.000 1028.930 800.000 ;
    END
  END reg2_idx0[4]
  PIN reg2_idx0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 1033.710 796.000 1033.990 800.000 ;
    END
  END reg2_idx0[5]
  PIN reg2_idx1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 103.400 2200.000 104.000 ;
    END
  END reg2_idx1[0]
  PIN reg2_idx1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.465000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 106.120 2200.000 106.720 ;
    END
  END reg2_idx1[1]
  PIN reg2_idx1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 108.840 2200.000 109.440 ;
    END
  END reg2_idx1[2]
  PIN reg2_idx1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.179000 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 111.560 2200.000 112.160 ;
    END
  END reg2_idx1[3]
  PIN reg2_idx1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.484000 ;
    ANTENNADIFFAREA 9.128699 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 114.280 2200.000 114.880 ;
    END
  END reg2_idx1[4]
  PIN reg2_idx1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.227500 ;
    ANTENNADIFFAREA 2.173500 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 117.000 2200.000 117.600 ;
    END
  END reg2_idx1[5]
  PIN reg2_idx2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.455000 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.960 4.000 98.560 ;
    END
  END reg2_idx2[0]
  PIN reg2_idx2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 4.000 101.280 ;
    END
  END reg2_idx2[1]
  PIN reg2_idx2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.400 4.000 104.000 ;
    END
  END reg2_idx2[2]
  PIN reg2_idx2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.822000 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.120 4.000 106.720 ;
    END
  END reg2_idx2[3]
  PIN reg2_idx2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.475000 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END reg2_idx2[4]
  PIN reg2_idx2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.832000 ;
    ANTENNADIFFAREA 2.173500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 111.560 4.000 112.160 ;
    END
  END reg2_idx2[5]
  PIN reg2_val0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1990.050 796.000 1990.330 800.000 ;
    END
  END reg2_val0[0]
  PIN reg2_val0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 2040.650 796.000 2040.930 800.000 ;
    END
  END reg2_val0[10]
  PIN reg2_val0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 2045.710 796.000 2045.990 800.000 ;
    END
  END reg2_val0[11]
  PIN reg2_val0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 2050.770 796.000 2051.050 800.000 ;
    END
  END reg2_val0[12]
  PIN reg2_val0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 2055.830 796.000 2056.110 800.000 ;
    END
  END reg2_val0[13]
  PIN reg2_val0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 2060.890 796.000 2061.170 800.000 ;
    END
  END reg2_val0[14]
  PIN reg2_val0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 2065.950 796.000 2066.230 800.000 ;
    END
  END reg2_val0[15]
  PIN reg2_val0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 2071.010 796.000 2071.290 800.000 ;
    END
  END reg2_val0[16]
  PIN reg2_val0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 2076.070 796.000 2076.350 800.000 ;
    END
  END reg2_val0[17]
  PIN reg2_val0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 2081.130 796.000 2081.410 800.000 ;
    END
  END reg2_val0[18]
  PIN reg2_val0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 2086.190 796.000 2086.470 800.000 ;
    END
  END reg2_val0[19]
  PIN reg2_val0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 1995.110 796.000 1995.390 800.000 ;
    END
  END reg2_val0[1]
  PIN reg2_val0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 2091.250 796.000 2091.530 800.000 ;
    END
  END reg2_val0[20]
  PIN reg2_val0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 2096.310 796.000 2096.590 800.000 ;
    END
  END reg2_val0[21]
  PIN reg2_val0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 2101.370 796.000 2101.650 800.000 ;
    END
  END reg2_val0[22]
  PIN reg2_val0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 2106.430 796.000 2106.710 800.000 ;
    END
  END reg2_val0[23]
  PIN reg2_val0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 2111.490 796.000 2111.770 800.000 ;
    END
  END reg2_val0[24]
  PIN reg2_val0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 2116.550 796.000 2116.830 800.000 ;
    END
  END reg2_val0[25]
  PIN reg2_val0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 2121.610 796.000 2121.890 800.000 ;
    END
  END reg2_val0[26]
  PIN reg2_val0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 2126.670 796.000 2126.950 800.000 ;
    END
  END reg2_val0[27]
  PIN reg2_val0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 2131.730 796.000 2132.010 800.000 ;
    END
  END reg2_val0[28]
  PIN reg2_val0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 2136.790 796.000 2137.070 800.000 ;
    END
  END reg2_val0[29]
  PIN reg2_val0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 2000.170 796.000 2000.450 800.000 ;
    END
  END reg2_val0[2]
  PIN reg2_val0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 2141.850 796.000 2142.130 800.000 ;
    END
  END reg2_val0[30]
  PIN reg2_val0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 2146.910 796.000 2147.190 800.000 ;
    END
  END reg2_val0[31]
  PIN reg2_val0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 2005.230 796.000 2005.510 800.000 ;
    END
  END reg2_val0[3]
  PIN reg2_val0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 2010.290 796.000 2010.570 800.000 ;
    END
  END reg2_val0[4]
  PIN reg2_val0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 2015.350 796.000 2015.630 800.000 ;
    END
  END reg2_val0[5]
  PIN reg2_val0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 2020.410 796.000 2020.690 800.000 ;
    END
  END reg2_val0[6]
  PIN reg2_val0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 2025.470 796.000 2025.750 800.000 ;
    END
  END reg2_val0[7]
  PIN reg2_val0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 2030.530 796.000 2030.810 800.000 ;
    END
  END reg2_val0[8]
  PIN reg2_val0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 2035.590 796.000 2035.870 800.000 ;
    END
  END reg2_val0[9]
  PIN reg2_val1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 631.080 2200.000 631.680 ;
    END
  END reg2_val1[0]
  PIN reg2_val1[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 658.280 2200.000 658.880 ;
    END
  END reg2_val1[10]
  PIN reg2_val1[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 661.000 2200.000 661.600 ;
    END
  END reg2_val1[11]
  PIN reg2_val1[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 663.720 2200.000 664.320 ;
    END
  END reg2_val1[12]
  PIN reg2_val1[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 666.440 2200.000 667.040 ;
    END
  END reg2_val1[13]
  PIN reg2_val1[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 669.160 2200.000 669.760 ;
    END
  END reg2_val1[14]
  PIN reg2_val1[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 671.880 2200.000 672.480 ;
    END
  END reg2_val1[15]
  PIN reg2_val1[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 674.600 2200.000 675.200 ;
    END
  END reg2_val1[16]
  PIN reg2_val1[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 677.320 2200.000 677.920 ;
    END
  END reg2_val1[17]
  PIN reg2_val1[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 680.040 2200.000 680.640 ;
    END
  END reg2_val1[18]
  PIN reg2_val1[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 682.760 2200.000 683.360 ;
    END
  END reg2_val1[19]
  PIN reg2_val1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 633.800 2200.000 634.400 ;
    END
  END reg2_val1[1]
  PIN reg2_val1[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 685.480 2200.000 686.080 ;
    END
  END reg2_val1[20]
  PIN reg2_val1[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 688.200 2200.000 688.800 ;
    END
  END reg2_val1[21]
  PIN reg2_val1[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 690.920 2200.000 691.520 ;
    END
  END reg2_val1[22]
  PIN reg2_val1[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 693.640 2200.000 694.240 ;
    END
  END reg2_val1[23]
  PIN reg2_val1[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 696.360 2200.000 696.960 ;
    END
  END reg2_val1[24]
  PIN reg2_val1[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 699.080 2200.000 699.680 ;
    END
  END reg2_val1[25]
  PIN reg2_val1[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 701.800 2200.000 702.400 ;
    END
  END reg2_val1[26]
  PIN reg2_val1[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 704.520 2200.000 705.120 ;
    END
  END reg2_val1[27]
  PIN reg2_val1[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 707.240 2200.000 707.840 ;
    END
  END reg2_val1[28]
  PIN reg2_val1[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 709.960 2200.000 710.560 ;
    END
  END reg2_val1[29]
  PIN reg2_val1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 636.520 2200.000 637.120 ;
    END
  END reg2_val1[2]
  PIN reg2_val1[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 712.680 2200.000 713.280 ;
    END
  END reg2_val1[30]
  PIN reg2_val1[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 715.400 2200.000 716.000 ;
    END
  END reg2_val1[31]
  PIN reg2_val1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 639.240 2200.000 639.840 ;
    END
  END reg2_val1[3]
  PIN reg2_val1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 641.960 2200.000 642.560 ;
    END
  END reg2_val1[4]
  PIN reg2_val1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 644.680 2200.000 645.280 ;
    END
  END reg2_val1[5]
  PIN reg2_val1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 647.400 2200.000 648.000 ;
    END
  END reg2_val1[6]
  PIN reg2_val1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 650.120 2200.000 650.720 ;
    END
  END reg2_val1[7]
  PIN reg2_val1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 652.840 2200.000 653.440 ;
    END
  END reg2_val1[8]
  PIN reg2_val1[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 655.560 2200.000 656.160 ;
    END
  END reg2_val1[9]
  PIN reg2_val2[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 625.640 4.000 626.240 ;
    END
  END reg2_val2[0]
  PIN reg2_val2[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 652.840 4.000 653.440 ;
    END
  END reg2_val2[10]
  PIN reg2_val2[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 655.560 4.000 656.160 ;
    END
  END reg2_val2[11]
  PIN reg2_val2[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 658.280 4.000 658.880 ;
    END
  END reg2_val2[12]
  PIN reg2_val2[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 661.000 4.000 661.600 ;
    END
  END reg2_val2[13]
  PIN reg2_val2[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 663.720 4.000 664.320 ;
    END
  END reg2_val2[14]
  PIN reg2_val2[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 666.440 4.000 667.040 ;
    END
  END reg2_val2[15]
  PIN reg2_val2[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 669.160 4.000 669.760 ;
    END
  END reg2_val2[16]
  PIN reg2_val2[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 671.880 4.000 672.480 ;
    END
  END reg2_val2[17]
  PIN reg2_val2[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 674.600 4.000 675.200 ;
    END
  END reg2_val2[18]
  PIN reg2_val2[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 677.320 4.000 677.920 ;
    END
  END reg2_val2[19]
  PIN reg2_val2[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 628.360 4.000 628.960 ;
    END
  END reg2_val2[1]
  PIN reg2_val2[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 680.040 4.000 680.640 ;
    END
  END reg2_val2[20]
  PIN reg2_val2[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 682.760 4.000 683.360 ;
    END
  END reg2_val2[21]
  PIN reg2_val2[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 685.480 4.000 686.080 ;
    END
  END reg2_val2[22]
  PIN reg2_val2[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 688.200 4.000 688.800 ;
    END
  END reg2_val2[23]
  PIN reg2_val2[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 690.920 4.000 691.520 ;
    END
  END reg2_val2[24]
  PIN reg2_val2[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 693.640 4.000 694.240 ;
    END
  END reg2_val2[25]
  PIN reg2_val2[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 696.360 4.000 696.960 ;
    END
  END reg2_val2[26]
  PIN reg2_val2[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 699.080 4.000 699.680 ;
    END
  END reg2_val2[27]
  PIN reg2_val2[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 701.800 4.000 702.400 ;
    END
  END reg2_val2[28]
  PIN reg2_val2[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 704.520 4.000 705.120 ;
    END
  END reg2_val2[29]
  PIN reg2_val2[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 631.080 4.000 631.680 ;
    END
  END reg2_val2[2]
  PIN reg2_val2[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 707.240 4.000 707.840 ;
    END
  END reg2_val2[30]
  PIN reg2_val2[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 709.960 4.000 710.560 ;
    END
  END reg2_val2[31]
  PIN reg2_val2[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 633.800 4.000 634.400 ;
    END
  END reg2_val2[3]
  PIN reg2_val2[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 636.520 4.000 637.120 ;
    END
  END reg2_val2[4]
  PIN reg2_val2[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 639.240 4.000 639.840 ;
    END
  END reg2_val2[5]
  PIN reg2_val2[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 641.960 4.000 642.560 ;
    END
  END reg2_val2[6]
  PIN reg2_val2[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 644.680 4.000 645.280 ;
    END
  END reg2_val2[7]
  PIN reg2_val2[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 647.400 4.000 648.000 ;
    END
  END reg2_val2[8]
  PIN reg2_val2[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 650.120 4.000 650.720 ;
    END
  END reg2_val2[9]
  PIN rst_eu
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.862000 ;
    PORT
      LAYER met2 ;
        RECT 831.310 796.000 831.590 800.000 ;
    END
  END rst_eu
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.086000 ;
    PORT
      LAYER met2 ;
        RECT 2113.330 0.000 2113.610 4.000 ;
    END
  END rst_n
  PIN sign_extend0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1448.630 796.000 1448.910 800.000 ;
    END
  END sign_extend0
  PIN sign_extend1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 340.040 2200.000 340.640 ;
    END
  END sign_extend1
  PIN sign_extend2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 334.600 4.000 335.200 ;
    END
  END sign_extend2
  PIN take_branch0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.415500 ;
    PORT
      LAYER met2 ;
        RECT 1463.810 796.000 1464.090 800.000 ;
    END
  END take_branch0
  PIN take_branch1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.710500 ;
    ANTENNADIFFAREA 2.608200 ;
    PORT
      LAYER met3 ;
        RECT 2196.000 348.200 2200.000 348.800 ;
    END
  END take_branch1
  PIN take_branch2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 342.760 4.000 343.360 ;
    END
  END take_branch2
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.040 10.640 1558.640 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1710.640 10.640 1712.240 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1864.240 10.640 1865.840 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2017.840 10.640 2019.440 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2171.440 10.640 2173.040 789.040 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1633.840 10.640 1635.440 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1787.440 10.640 1789.040 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1941.040 10.640 1942.640 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2094.640 10.640 2096.240 789.040 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 2104.590 0.000 2104.870 4.000 ;
    END
  END wb_clk_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2194.200 788.885 ;
      LAYER met1 ;
        RECT 5.520 0.380 2196.890 798.620 ;
      LAYER met2 ;
        RECT 6.530 795.720 41.670 798.650 ;
        RECT 42.510 795.720 46.730 798.650 ;
        RECT 47.570 795.720 51.790 798.650 ;
        RECT 52.630 795.720 56.850 798.650 ;
        RECT 57.690 795.720 61.910 798.650 ;
        RECT 62.750 795.720 66.970 798.650 ;
        RECT 67.810 795.720 72.030 798.650 ;
        RECT 72.870 795.720 77.090 798.650 ;
        RECT 77.930 795.720 82.150 798.650 ;
        RECT 82.990 795.720 87.210 798.650 ;
        RECT 88.050 795.720 92.270 798.650 ;
        RECT 93.110 795.720 97.330 798.650 ;
        RECT 98.170 795.720 102.390 798.650 ;
        RECT 103.230 795.720 107.450 798.650 ;
        RECT 108.290 795.720 112.510 798.650 ;
        RECT 113.350 795.720 117.570 798.650 ;
        RECT 118.410 795.720 122.630 798.650 ;
        RECT 123.470 795.720 127.690 798.650 ;
        RECT 128.530 795.720 132.750 798.650 ;
        RECT 133.590 795.720 137.810 798.650 ;
        RECT 138.650 795.720 142.870 798.650 ;
        RECT 143.710 795.720 147.930 798.650 ;
        RECT 148.770 795.720 152.990 798.650 ;
        RECT 153.830 795.720 158.050 798.650 ;
        RECT 158.890 795.720 163.110 798.650 ;
        RECT 163.950 795.720 168.170 798.650 ;
        RECT 169.010 795.720 173.230 798.650 ;
        RECT 174.070 795.720 178.290 798.650 ;
        RECT 179.130 795.720 183.350 798.650 ;
        RECT 184.190 795.720 188.410 798.650 ;
        RECT 189.250 795.720 193.470 798.650 ;
        RECT 194.310 795.720 198.530 798.650 ;
        RECT 199.370 795.720 203.590 798.650 ;
        RECT 204.430 795.720 208.650 798.650 ;
        RECT 209.490 795.720 213.710 798.650 ;
        RECT 214.550 795.720 218.770 798.650 ;
        RECT 219.610 795.720 223.830 798.650 ;
        RECT 224.670 795.720 228.890 798.650 ;
        RECT 229.730 795.720 233.950 798.650 ;
        RECT 234.790 795.720 239.010 798.650 ;
        RECT 239.850 795.720 244.070 798.650 ;
        RECT 244.910 795.720 249.130 798.650 ;
        RECT 249.970 795.720 254.190 798.650 ;
        RECT 255.030 795.720 259.250 798.650 ;
        RECT 260.090 795.720 264.310 798.650 ;
        RECT 265.150 795.720 269.370 798.650 ;
        RECT 270.210 795.720 274.430 798.650 ;
        RECT 275.270 795.720 279.490 798.650 ;
        RECT 280.330 795.720 284.550 798.650 ;
        RECT 285.390 795.720 289.610 798.650 ;
        RECT 290.450 795.720 294.670 798.650 ;
        RECT 295.510 795.720 299.730 798.650 ;
        RECT 300.570 795.720 304.790 798.650 ;
        RECT 305.630 795.720 309.850 798.650 ;
        RECT 310.690 795.720 314.910 798.650 ;
        RECT 315.750 795.720 319.970 798.650 ;
        RECT 320.810 795.720 325.030 798.650 ;
        RECT 325.870 795.720 330.090 798.650 ;
        RECT 330.930 795.720 335.150 798.650 ;
        RECT 335.990 795.720 340.210 798.650 ;
        RECT 341.050 795.720 345.270 798.650 ;
        RECT 346.110 795.720 350.330 798.650 ;
        RECT 351.170 795.720 355.390 798.650 ;
        RECT 356.230 795.720 360.450 798.650 ;
        RECT 361.290 795.720 365.510 798.650 ;
        RECT 366.350 795.720 370.570 798.650 ;
        RECT 371.410 795.720 375.630 798.650 ;
        RECT 376.470 795.720 380.690 798.650 ;
        RECT 381.530 795.720 385.750 798.650 ;
        RECT 386.590 795.720 390.810 798.650 ;
        RECT 391.650 795.720 395.870 798.650 ;
        RECT 396.710 795.720 400.930 798.650 ;
        RECT 401.770 795.720 405.990 798.650 ;
        RECT 406.830 795.720 411.050 798.650 ;
        RECT 411.890 795.720 416.110 798.650 ;
        RECT 416.950 795.720 421.170 798.650 ;
        RECT 422.010 795.720 426.230 798.650 ;
        RECT 427.070 795.720 431.290 798.650 ;
        RECT 432.130 795.720 436.350 798.650 ;
        RECT 437.190 795.720 441.410 798.650 ;
        RECT 442.250 795.720 446.470 798.650 ;
        RECT 447.310 795.720 451.530 798.650 ;
        RECT 452.370 795.720 456.590 798.650 ;
        RECT 457.430 795.720 461.650 798.650 ;
        RECT 462.490 795.720 466.710 798.650 ;
        RECT 467.550 795.720 471.770 798.650 ;
        RECT 472.610 795.720 476.830 798.650 ;
        RECT 477.670 795.720 481.890 798.650 ;
        RECT 482.730 795.720 486.950 798.650 ;
        RECT 487.790 795.720 492.010 798.650 ;
        RECT 492.850 795.720 497.070 798.650 ;
        RECT 497.910 795.720 502.130 798.650 ;
        RECT 502.970 795.720 507.190 798.650 ;
        RECT 508.030 795.720 512.250 798.650 ;
        RECT 513.090 795.720 517.310 798.650 ;
        RECT 518.150 795.720 522.370 798.650 ;
        RECT 523.210 795.720 527.430 798.650 ;
        RECT 528.270 795.720 532.490 798.650 ;
        RECT 533.330 795.720 537.550 798.650 ;
        RECT 538.390 795.720 542.610 798.650 ;
        RECT 543.450 795.720 547.670 798.650 ;
        RECT 548.510 795.720 552.730 798.650 ;
        RECT 553.570 795.720 557.790 798.650 ;
        RECT 558.630 795.720 562.850 798.650 ;
        RECT 563.690 795.720 567.910 798.650 ;
        RECT 568.750 795.720 572.970 798.650 ;
        RECT 573.810 795.720 578.030 798.650 ;
        RECT 578.870 795.720 583.090 798.650 ;
        RECT 583.930 795.720 588.150 798.650 ;
        RECT 588.990 795.720 593.210 798.650 ;
        RECT 594.050 795.720 598.270 798.650 ;
        RECT 599.110 795.720 603.330 798.650 ;
        RECT 604.170 795.720 608.390 798.650 ;
        RECT 609.230 795.720 613.450 798.650 ;
        RECT 614.290 795.720 618.510 798.650 ;
        RECT 619.350 795.720 623.570 798.650 ;
        RECT 624.410 795.720 628.630 798.650 ;
        RECT 629.470 795.720 633.690 798.650 ;
        RECT 634.530 795.720 638.750 798.650 ;
        RECT 639.590 795.720 643.810 798.650 ;
        RECT 644.650 795.720 648.870 798.650 ;
        RECT 649.710 795.720 653.930 798.650 ;
        RECT 654.770 795.720 658.990 798.650 ;
        RECT 659.830 795.720 664.050 798.650 ;
        RECT 664.890 795.720 669.110 798.650 ;
        RECT 669.950 795.720 674.170 798.650 ;
        RECT 675.010 795.720 679.230 798.650 ;
        RECT 680.070 795.720 684.290 798.650 ;
        RECT 685.130 795.720 689.350 798.650 ;
        RECT 690.190 795.720 694.410 798.650 ;
        RECT 695.250 795.720 699.470 798.650 ;
        RECT 700.310 795.720 704.530 798.650 ;
        RECT 705.370 795.720 709.590 798.650 ;
        RECT 710.430 795.720 714.650 798.650 ;
        RECT 715.490 795.720 719.710 798.650 ;
        RECT 720.550 795.720 724.770 798.650 ;
        RECT 725.610 795.720 729.830 798.650 ;
        RECT 730.670 795.720 734.890 798.650 ;
        RECT 735.730 795.720 739.950 798.650 ;
        RECT 740.790 795.720 745.010 798.650 ;
        RECT 745.850 795.720 750.070 798.650 ;
        RECT 750.910 795.720 755.130 798.650 ;
        RECT 755.970 795.720 760.190 798.650 ;
        RECT 761.030 795.720 765.250 798.650 ;
        RECT 766.090 795.720 770.310 798.650 ;
        RECT 771.150 795.720 775.370 798.650 ;
        RECT 776.210 795.720 780.430 798.650 ;
        RECT 781.270 795.720 785.490 798.650 ;
        RECT 786.330 795.720 790.550 798.650 ;
        RECT 791.390 795.720 795.610 798.650 ;
        RECT 796.450 795.720 800.670 798.650 ;
        RECT 801.510 795.720 805.730 798.650 ;
        RECT 806.570 795.720 810.790 798.650 ;
        RECT 811.630 795.720 815.850 798.650 ;
        RECT 816.690 795.720 820.910 798.650 ;
        RECT 821.750 795.720 825.970 798.650 ;
        RECT 826.810 795.720 831.030 798.650 ;
        RECT 831.870 795.720 836.090 798.650 ;
        RECT 836.930 795.720 841.150 798.650 ;
        RECT 841.990 795.720 846.210 798.650 ;
        RECT 847.050 795.720 851.270 798.650 ;
        RECT 852.110 795.720 856.330 798.650 ;
        RECT 857.170 795.720 861.390 798.650 ;
        RECT 862.230 795.720 866.450 798.650 ;
        RECT 867.290 795.720 871.510 798.650 ;
        RECT 872.350 795.720 876.570 798.650 ;
        RECT 877.410 795.720 881.630 798.650 ;
        RECT 882.470 795.720 886.690 798.650 ;
        RECT 887.530 795.720 891.750 798.650 ;
        RECT 892.590 795.720 896.810 798.650 ;
        RECT 897.650 795.720 901.870 798.650 ;
        RECT 902.710 795.720 906.930 798.650 ;
        RECT 907.770 795.720 911.990 798.650 ;
        RECT 912.830 795.720 917.050 798.650 ;
        RECT 917.890 795.720 922.110 798.650 ;
        RECT 922.950 795.720 927.170 798.650 ;
        RECT 928.010 795.720 932.230 798.650 ;
        RECT 933.070 795.720 937.290 798.650 ;
        RECT 938.130 795.720 942.350 798.650 ;
        RECT 943.190 795.720 947.410 798.650 ;
        RECT 948.250 795.720 952.470 798.650 ;
        RECT 953.310 795.720 957.530 798.650 ;
        RECT 958.370 795.720 962.590 798.650 ;
        RECT 963.430 795.720 967.650 798.650 ;
        RECT 968.490 795.720 972.710 798.650 ;
        RECT 973.550 795.720 977.770 798.650 ;
        RECT 978.610 795.720 982.830 798.650 ;
        RECT 983.670 795.720 987.890 798.650 ;
        RECT 988.730 795.720 992.950 798.650 ;
        RECT 993.790 795.720 998.010 798.650 ;
        RECT 998.850 795.720 1003.070 798.650 ;
        RECT 1003.910 795.720 1008.130 798.650 ;
        RECT 1008.970 795.720 1013.190 798.650 ;
        RECT 1014.030 795.720 1018.250 798.650 ;
        RECT 1019.090 795.720 1023.310 798.650 ;
        RECT 1024.150 795.720 1028.370 798.650 ;
        RECT 1029.210 795.720 1033.430 798.650 ;
        RECT 1034.270 795.720 1038.490 798.650 ;
        RECT 1039.330 795.720 1043.550 798.650 ;
        RECT 1044.390 795.720 1048.610 798.650 ;
        RECT 1049.450 795.720 1053.670 798.650 ;
        RECT 1054.510 795.720 1058.730 798.650 ;
        RECT 1059.570 795.720 1063.790 798.650 ;
        RECT 1064.630 795.720 1068.850 798.650 ;
        RECT 1069.690 795.720 1073.910 798.650 ;
        RECT 1074.750 795.720 1078.970 798.650 ;
        RECT 1079.810 795.720 1084.030 798.650 ;
        RECT 1084.870 795.720 1089.090 798.650 ;
        RECT 1089.930 795.720 1094.150 798.650 ;
        RECT 1094.990 795.720 1099.210 798.650 ;
        RECT 1100.050 795.720 1104.270 798.650 ;
        RECT 1105.110 795.720 1109.330 798.650 ;
        RECT 1110.170 795.720 1114.390 798.650 ;
        RECT 1115.230 795.720 1119.450 798.650 ;
        RECT 1120.290 795.720 1124.510 798.650 ;
        RECT 1125.350 795.720 1129.570 798.650 ;
        RECT 1130.410 795.720 1134.630 798.650 ;
        RECT 1135.470 795.720 1139.690 798.650 ;
        RECT 1140.530 795.720 1144.750 798.650 ;
        RECT 1145.590 795.720 1149.810 798.650 ;
        RECT 1150.650 795.720 1154.870 798.650 ;
        RECT 1155.710 795.720 1159.930 798.650 ;
        RECT 1160.770 795.720 1164.990 798.650 ;
        RECT 1165.830 795.720 1170.050 798.650 ;
        RECT 1170.890 795.720 1175.110 798.650 ;
        RECT 1175.950 795.720 1180.170 798.650 ;
        RECT 1181.010 795.720 1185.230 798.650 ;
        RECT 1186.070 795.720 1190.290 798.650 ;
        RECT 1191.130 795.720 1195.350 798.650 ;
        RECT 1196.190 795.720 1200.410 798.650 ;
        RECT 1201.250 795.720 1205.470 798.650 ;
        RECT 1206.310 795.720 1210.530 798.650 ;
        RECT 1211.370 795.720 1215.590 798.650 ;
        RECT 1216.430 795.720 1220.650 798.650 ;
        RECT 1221.490 795.720 1225.710 798.650 ;
        RECT 1226.550 795.720 1230.770 798.650 ;
        RECT 1231.610 795.720 1235.830 798.650 ;
        RECT 1236.670 795.720 1240.890 798.650 ;
        RECT 1241.730 795.720 1245.950 798.650 ;
        RECT 1246.790 795.720 1251.010 798.650 ;
        RECT 1251.850 795.720 1256.070 798.650 ;
        RECT 1256.910 795.720 1261.130 798.650 ;
        RECT 1261.970 795.720 1266.190 798.650 ;
        RECT 1267.030 795.720 1271.250 798.650 ;
        RECT 1272.090 795.720 1276.310 798.650 ;
        RECT 1277.150 795.720 1281.370 798.650 ;
        RECT 1282.210 795.720 1286.430 798.650 ;
        RECT 1287.270 795.720 1291.490 798.650 ;
        RECT 1292.330 795.720 1296.550 798.650 ;
        RECT 1297.390 795.720 1301.610 798.650 ;
        RECT 1302.450 795.720 1306.670 798.650 ;
        RECT 1307.510 795.720 1311.730 798.650 ;
        RECT 1312.570 795.720 1316.790 798.650 ;
        RECT 1317.630 795.720 1321.850 798.650 ;
        RECT 1322.690 795.720 1326.910 798.650 ;
        RECT 1327.750 795.720 1331.970 798.650 ;
        RECT 1332.810 795.720 1337.030 798.650 ;
        RECT 1337.870 795.720 1342.090 798.650 ;
        RECT 1342.930 795.720 1347.150 798.650 ;
        RECT 1347.990 795.720 1352.210 798.650 ;
        RECT 1353.050 795.720 1357.270 798.650 ;
        RECT 1358.110 795.720 1362.330 798.650 ;
        RECT 1363.170 795.720 1367.390 798.650 ;
        RECT 1368.230 795.720 1372.450 798.650 ;
        RECT 1373.290 795.720 1377.510 798.650 ;
        RECT 1378.350 795.720 1382.570 798.650 ;
        RECT 1383.410 795.720 1387.630 798.650 ;
        RECT 1388.470 795.720 1392.690 798.650 ;
        RECT 1393.530 795.720 1397.750 798.650 ;
        RECT 1398.590 795.720 1402.810 798.650 ;
        RECT 1403.650 795.720 1407.870 798.650 ;
        RECT 1408.710 795.720 1412.930 798.650 ;
        RECT 1413.770 795.720 1417.990 798.650 ;
        RECT 1418.830 795.720 1423.050 798.650 ;
        RECT 1423.890 795.720 1428.110 798.650 ;
        RECT 1428.950 795.720 1433.170 798.650 ;
        RECT 1434.010 795.720 1438.230 798.650 ;
        RECT 1439.070 795.720 1443.290 798.650 ;
        RECT 1444.130 795.720 1448.350 798.650 ;
        RECT 1449.190 795.720 1453.410 798.650 ;
        RECT 1454.250 795.720 1458.470 798.650 ;
        RECT 1459.310 795.720 1463.530 798.650 ;
        RECT 1464.370 795.720 1468.590 798.650 ;
        RECT 1469.430 795.720 1473.650 798.650 ;
        RECT 1474.490 795.720 1478.710 798.650 ;
        RECT 1479.550 795.720 1483.770 798.650 ;
        RECT 1484.610 795.720 1488.830 798.650 ;
        RECT 1489.670 795.720 1493.890 798.650 ;
        RECT 1494.730 795.720 1498.950 798.650 ;
        RECT 1499.790 795.720 1504.010 798.650 ;
        RECT 1504.850 795.720 1509.070 798.650 ;
        RECT 1509.910 795.720 1514.130 798.650 ;
        RECT 1514.970 795.720 1519.190 798.650 ;
        RECT 1520.030 795.720 1524.250 798.650 ;
        RECT 1525.090 795.720 1529.310 798.650 ;
        RECT 1530.150 795.720 1534.370 798.650 ;
        RECT 1535.210 795.720 1539.430 798.650 ;
        RECT 1540.270 795.720 1544.490 798.650 ;
        RECT 1545.330 795.720 1549.550 798.650 ;
        RECT 1550.390 795.720 1554.610 798.650 ;
        RECT 1555.450 795.720 1559.670 798.650 ;
        RECT 1560.510 795.720 1564.730 798.650 ;
        RECT 1565.570 795.720 1569.790 798.650 ;
        RECT 1570.630 795.720 1574.850 798.650 ;
        RECT 1575.690 795.720 1579.910 798.650 ;
        RECT 1580.750 795.720 1584.970 798.650 ;
        RECT 1585.810 795.720 1590.030 798.650 ;
        RECT 1590.870 795.720 1595.090 798.650 ;
        RECT 1595.930 795.720 1600.150 798.650 ;
        RECT 1600.990 795.720 1605.210 798.650 ;
        RECT 1606.050 795.720 1610.270 798.650 ;
        RECT 1611.110 795.720 1615.330 798.650 ;
        RECT 1616.170 795.720 1620.390 798.650 ;
        RECT 1621.230 795.720 1625.450 798.650 ;
        RECT 1626.290 795.720 1630.510 798.650 ;
        RECT 1631.350 795.720 1635.570 798.650 ;
        RECT 1636.410 795.720 1640.630 798.650 ;
        RECT 1641.470 795.720 1645.690 798.650 ;
        RECT 1646.530 795.720 1650.750 798.650 ;
        RECT 1651.590 795.720 1655.810 798.650 ;
        RECT 1656.650 795.720 1660.870 798.650 ;
        RECT 1661.710 795.720 1665.930 798.650 ;
        RECT 1666.770 795.720 1670.990 798.650 ;
        RECT 1671.830 795.720 1676.050 798.650 ;
        RECT 1676.890 795.720 1681.110 798.650 ;
        RECT 1681.950 795.720 1686.170 798.650 ;
        RECT 1687.010 795.720 1691.230 798.650 ;
        RECT 1692.070 795.720 1696.290 798.650 ;
        RECT 1697.130 795.720 1701.350 798.650 ;
        RECT 1702.190 795.720 1706.410 798.650 ;
        RECT 1707.250 795.720 1711.470 798.650 ;
        RECT 1712.310 795.720 1716.530 798.650 ;
        RECT 1717.370 795.720 1721.590 798.650 ;
        RECT 1722.430 795.720 1726.650 798.650 ;
        RECT 1727.490 795.720 1731.710 798.650 ;
        RECT 1732.550 795.720 1736.770 798.650 ;
        RECT 1737.610 795.720 1741.830 798.650 ;
        RECT 1742.670 795.720 1746.890 798.650 ;
        RECT 1747.730 795.720 1751.950 798.650 ;
        RECT 1752.790 795.720 1757.010 798.650 ;
        RECT 1757.850 795.720 1762.070 798.650 ;
        RECT 1762.910 795.720 1767.130 798.650 ;
        RECT 1767.970 795.720 1772.190 798.650 ;
        RECT 1773.030 795.720 1777.250 798.650 ;
        RECT 1778.090 795.720 1782.310 798.650 ;
        RECT 1783.150 795.720 1787.370 798.650 ;
        RECT 1788.210 795.720 1792.430 798.650 ;
        RECT 1793.270 795.720 1797.490 798.650 ;
        RECT 1798.330 795.720 1802.550 798.650 ;
        RECT 1803.390 795.720 1807.610 798.650 ;
        RECT 1808.450 795.720 1812.670 798.650 ;
        RECT 1813.510 795.720 1817.730 798.650 ;
        RECT 1818.570 795.720 1822.790 798.650 ;
        RECT 1823.630 795.720 1827.850 798.650 ;
        RECT 1828.690 795.720 1832.910 798.650 ;
        RECT 1833.750 795.720 1837.970 798.650 ;
        RECT 1838.810 795.720 1843.030 798.650 ;
        RECT 1843.870 795.720 1848.090 798.650 ;
        RECT 1848.930 795.720 1853.150 798.650 ;
        RECT 1853.990 795.720 1858.210 798.650 ;
        RECT 1859.050 795.720 1863.270 798.650 ;
        RECT 1864.110 795.720 1868.330 798.650 ;
        RECT 1869.170 795.720 1873.390 798.650 ;
        RECT 1874.230 795.720 1878.450 798.650 ;
        RECT 1879.290 795.720 1883.510 798.650 ;
        RECT 1884.350 795.720 1888.570 798.650 ;
        RECT 1889.410 795.720 1893.630 798.650 ;
        RECT 1894.470 795.720 1898.690 798.650 ;
        RECT 1899.530 795.720 1903.750 798.650 ;
        RECT 1904.590 795.720 1908.810 798.650 ;
        RECT 1909.650 795.720 1913.870 798.650 ;
        RECT 1914.710 795.720 1918.930 798.650 ;
        RECT 1919.770 795.720 1923.990 798.650 ;
        RECT 1924.830 795.720 1929.050 798.650 ;
        RECT 1929.890 795.720 1934.110 798.650 ;
        RECT 1934.950 795.720 1939.170 798.650 ;
        RECT 1940.010 795.720 1944.230 798.650 ;
        RECT 1945.070 795.720 1949.290 798.650 ;
        RECT 1950.130 795.720 1954.350 798.650 ;
        RECT 1955.190 795.720 1959.410 798.650 ;
        RECT 1960.250 795.720 1964.470 798.650 ;
        RECT 1965.310 795.720 1969.530 798.650 ;
        RECT 1970.370 795.720 1974.590 798.650 ;
        RECT 1975.430 795.720 1979.650 798.650 ;
        RECT 1980.490 795.720 1984.710 798.650 ;
        RECT 1985.550 795.720 1989.770 798.650 ;
        RECT 1990.610 795.720 1994.830 798.650 ;
        RECT 1995.670 795.720 1999.890 798.650 ;
        RECT 2000.730 795.720 2004.950 798.650 ;
        RECT 2005.790 795.720 2010.010 798.650 ;
        RECT 2010.850 795.720 2015.070 798.650 ;
        RECT 2015.910 795.720 2020.130 798.650 ;
        RECT 2020.970 795.720 2025.190 798.650 ;
        RECT 2026.030 795.720 2030.250 798.650 ;
        RECT 2031.090 795.720 2035.310 798.650 ;
        RECT 2036.150 795.720 2040.370 798.650 ;
        RECT 2041.210 795.720 2045.430 798.650 ;
        RECT 2046.270 795.720 2050.490 798.650 ;
        RECT 2051.330 795.720 2055.550 798.650 ;
        RECT 2056.390 795.720 2060.610 798.650 ;
        RECT 2061.450 795.720 2065.670 798.650 ;
        RECT 2066.510 795.720 2070.730 798.650 ;
        RECT 2071.570 795.720 2075.790 798.650 ;
        RECT 2076.630 795.720 2080.850 798.650 ;
        RECT 2081.690 795.720 2085.910 798.650 ;
        RECT 2086.750 795.720 2090.970 798.650 ;
        RECT 2091.810 795.720 2096.030 798.650 ;
        RECT 2096.870 795.720 2101.090 798.650 ;
        RECT 2101.930 795.720 2106.150 798.650 ;
        RECT 2106.990 795.720 2111.210 798.650 ;
        RECT 2112.050 795.720 2116.270 798.650 ;
        RECT 2117.110 795.720 2121.330 798.650 ;
        RECT 2122.170 795.720 2126.390 798.650 ;
        RECT 2127.230 795.720 2131.450 798.650 ;
        RECT 2132.290 795.720 2136.510 798.650 ;
        RECT 2137.350 795.720 2141.570 798.650 ;
        RECT 2142.410 795.720 2146.630 798.650 ;
        RECT 2147.470 795.720 2151.690 798.650 ;
        RECT 2152.530 795.720 2156.750 798.650 ;
        RECT 2157.590 795.720 2196.860 798.650 ;
        RECT 6.530 4.280 2196.860 795.720 ;
        RECT 6.530 0.350 41.670 4.280 ;
        RECT 42.510 0.350 50.410 4.280 ;
        RECT 51.250 0.350 59.150 4.280 ;
        RECT 59.990 0.350 67.890 4.280 ;
        RECT 68.730 0.350 76.630 4.280 ;
        RECT 77.470 0.350 85.370 4.280 ;
        RECT 86.210 0.350 94.110 4.280 ;
        RECT 94.950 0.350 102.850 4.280 ;
        RECT 103.690 0.350 111.590 4.280 ;
        RECT 112.430 0.350 120.330 4.280 ;
        RECT 121.170 0.350 129.070 4.280 ;
        RECT 129.910 0.350 137.810 4.280 ;
        RECT 138.650 0.350 146.550 4.280 ;
        RECT 147.390 0.350 155.290 4.280 ;
        RECT 156.130 0.350 164.030 4.280 ;
        RECT 164.870 0.350 172.770 4.280 ;
        RECT 173.610 0.350 181.510 4.280 ;
        RECT 182.350 0.350 190.250 4.280 ;
        RECT 191.090 0.350 198.990 4.280 ;
        RECT 199.830 0.350 207.730 4.280 ;
        RECT 208.570 0.350 216.470 4.280 ;
        RECT 217.310 0.350 225.210 4.280 ;
        RECT 226.050 0.350 233.950 4.280 ;
        RECT 234.790 0.350 242.690 4.280 ;
        RECT 243.530 0.350 251.430 4.280 ;
        RECT 252.270 0.350 260.170 4.280 ;
        RECT 261.010 0.350 268.910 4.280 ;
        RECT 269.750 0.350 277.650 4.280 ;
        RECT 278.490 0.350 286.390 4.280 ;
        RECT 287.230 0.350 295.130 4.280 ;
        RECT 295.970 0.350 303.870 4.280 ;
        RECT 304.710 0.350 312.610 4.280 ;
        RECT 313.450 0.350 321.350 4.280 ;
        RECT 322.190 0.350 330.090 4.280 ;
        RECT 330.930 0.350 338.830 4.280 ;
        RECT 339.670 0.350 347.570 4.280 ;
        RECT 348.410 0.350 356.310 4.280 ;
        RECT 357.150 0.350 365.050 4.280 ;
        RECT 365.890 0.350 373.790 4.280 ;
        RECT 374.630 0.350 382.530 4.280 ;
        RECT 383.370 0.350 391.270 4.280 ;
        RECT 392.110 0.350 400.010 4.280 ;
        RECT 400.850 0.350 408.750 4.280 ;
        RECT 409.590 0.350 417.490 4.280 ;
        RECT 418.330 0.350 426.230 4.280 ;
        RECT 427.070 0.350 434.970 4.280 ;
        RECT 435.810 0.350 443.710 4.280 ;
        RECT 444.550 0.350 452.450 4.280 ;
        RECT 453.290 0.350 461.190 4.280 ;
        RECT 462.030 0.350 469.930 4.280 ;
        RECT 470.770 0.350 478.670 4.280 ;
        RECT 479.510 0.350 487.410 4.280 ;
        RECT 488.250 0.350 496.150 4.280 ;
        RECT 496.990 0.350 504.890 4.280 ;
        RECT 505.730 0.350 513.630 4.280 ;
        RECT 514.470 0.350 522.370 4.280 ;
        RECT 523.210 0.350 531.110 4.280 ;
        RECT 531.950 0.350 539.850 4.280 ;
        RECT 540.690 0.350 548.590 4.280 ;
        RECT 549.430 0.350 557.330 4.280 ;
        RECT 558.170 0.350 566.070 4.280 ;
        RECT 566.910 0.350 574.810 4.280 ;
        RECT 575.650 0.350 583.550 4.280 ;
        RECT 584.390 0.350 592.290 4.280 ;
        RECT 593.130 0.350 601.030 4.280 ;
        RECT 601.870 0.350 609.770 4.280 ;
        RECT 610.610 0.350 618.510 4.280 ;
        RECT 619.350 0.350 627.250 4.280 ;
        RECT 628.090 0.350 635.990 4.280 ;
        RECT 636.830 0.350 644.730 4.280 ;
        RECT 645.570 0.350 653.470 4.280 ;
        RECT 654.310 0.350 662.210 4.280 ;
        RECT 663.050 0.350 670.950 4.280 ;
        RECT 671.790 0.350 679.690 4.280 ;
        RECT 680.530 0.350 688.430 4.280 ;
        RECT 689.270 0.350 697.170 4.280 ;
        RECT 698.010 0.350 705.910 4.280 ;
        RECT 706.750 0.350 714.650 4.280 ;
        RECT 715.490 0.350 723.390 4.280 ;
        RECT 724.230 0.350 732.130 4.280 ;
        RECT 732.970 0.350 740.870 4.280 ;
        RECT 741.710 0.350 749.610 4.280 ;
        RECT 750.450 0.350 758.350 4.280 ;
        RECT 759.190 0.350 767.090 4.280 ;
        RECT 767.930 0.350 775.830 4.280 ;
        RECT 776.670 0.350 784.570 4.280 ;
        RECT 785.410 0.350 793.310 4.280 ;
        RECT 794.150 0.350 802.050 4.280 ;
        RECT 802.890 0.350 810.790 4.280 ;
        RECT 811.630 0.350 819.530 4.280 ;
        RECT 820.370 0.350 828.270 4.280 ;
        RECT 829.110 0.350 837.010 4.280 ;
        RECT 837.850 0.350 845.750 4.280 ;
        RECT 846.590 0.350 854.490 4.280 ;
        RECT 855.330 0.350 863.230 4.280 ;
        RECT 864.070 0.350 871.970 4.280 ;
        RECT 872.810 0.350 880.710 4.280 ;
        RECT 881.550 0.350 889.450 4.280 ;
        RECT 890.290 0.350 898.190 4.280 ;
        RECT 899.030 0.350 906.930 4.280 ;
        RECT 907.770 0.350 915.670 4.280 ;
        RECT 916.510 0.350 924.410 4.280 ;
        RECT 925.250 0.350 933.150 4.280 ;
        RECT 933.990 0.350 941.890 4.280 ;
        RECT 942.730 0.350 950.630 4.280 ;
        RECT 951.470 0.350 959.370 4.280 ;
        RECT 960.210 0.350 968.110 4.280 ;
        RECT 968.950 0.350 976.850 4.280 ;
        RECT 977.690 0.350 985.590 4.280 ;
        RECT 986.430 0.350 994.330 4.280 ;
        RECT 995.170 0.350 1003.070 4.280 ;
        RECT 1003.910 0.350 1011.810 4.280 ;
        RECT 1012.650 0.350 1020.550 4.280 ;
        RECT 1021.390 0.350 1029.290 4.280 ;
        RECT 1030.130 0.350 1038.030 4.280 ;
        RECT 1038.870 0.350 1046.770 4.280 ;
        RECT 1047.610 0.350 1055.510 4.280 ;
        RECT 1056.350 0.350 1064.250 4.280 ;
        RECT 1065.090 0.350 1072.990 4.280 ;
        RECT 1073.830 0.350 1081.730 4.280 ;
        RECT 1082.570 0.350 1090.470 4.280 ;
        RECT 1091.310 0.350 1099.210 4.280 ;
        RECT 1100.050 0.350 1107.950 4.280 ;
        RECT 1108.790 0.350 1116.690 4.280 ;
        RECT 1117.530 0.350 1125.430 4.280 ;
        RECT 1126.270 0.350 1134.170 4.280 ;
        RECT 1135.010 0.350 1142.910 4.280 ;
        RECT 1143.750 0.350 1151.650 4.280 ;
        RECT 1152.490 0.350 1160.390 4.280 ;
        RECT 1161.230 0.350 1169.130 4.280 ;
        RECT 1169.970 0.350 1177.870 4.280 ;
        RECT 1178.710 0.350 1186.610 4.280 ;
        RECT 1187.450 0.350 1195.350 4.280 ;
        RECT 1196.190 0.350 1204.090 4.280 ;
        RECT 1204.930 0.350 1212.830 4.280 ;
        RECT 1213.670 0.350 1221.570 4.280 ;
        RECT 1222.410 0.350 1230.310 4.280 ;
        RECT 1231.150 0.350 1239.050 4.280 ;
        RECT 1239.890 0.350 1247.790 4.280 ;
        RECT 1248.630 0.350 1256.530 4.280 ;
        RECT 1257.370 0.350 1265.270 4.280 ;
        RECT 1266.110 0.350 1274.010 4.280 ;
        RECT 1274.850 0.350 1282.750 4.280 ;
        RECT 1283.590 0.350 1291.490 4.280 ;
        RECT 1292.330 0.350 1300.230 4.280 ;
        RECT 1301.070 0.350 1308.970 4.280 ;
        RECT 1309.810 0.350 1317.710 4.280 ;
        RECT 1318.550 0.350 1326.450 4.280 ;
        RECT 1327.290 0.350 1335.190 4.280 ;
        RECT 1336.030 0.350 1343.930 4.280 ;
        RECT 1344.770 0.350 1352.670 4.280 ;
        RECT 1353.510 0.350 1361.410 4.280 ;
        RECT 1362.250 0.350 1370.150 4.280 ;
        RECT 1370.990 0.350 1378.890 4.280 ;
        RECT 1379.730 0.350 1387.630 4.280 ;
        RECT 1388.470 0.350 1396.370 4.280 ;
        RECT 1397.210 0.350 1405.110 4.280 ;
        RECT 1405.950 0.350 1413.850 4.280 ;
        RECT 1414.690 0.350 1422.590 4.280 ;
        RECT 1423.430 0.350 1431.330 4.280 ;
        RECT 1432.170 0.350 1440.070 4.280 ;
        RECT 1440.910 0.350 1448.810 4.280 ;
        RECT 1449.650 0.350 1457.550 4.280 ;
        RECT 1458.390 0.350 1466.290 4.280 ;
        RECT 1467.130 0.350 1475.030 4.280 ;
        RECT 1475.870 0.350 1483.770 4.280 ;
        RECT 1484.610 0.350 1492.510 4.280 ;
        RECT 1493.350 0.350 1501.250 4.280 ;
        RECT 1502.090 0.350 1509.990 4.280 ;
        RECT 1510.830 0.350 1518.730 4.280 ;
        RECT 1519.570 0.350 1527.470 4.280 ;
        RECT 1528.310 0.350 1536.210 4.280 ;
        RECT 1537.050 0.350 1544.950 4.280 ;
        RECT 1545.790 0.350 1553.690 4.280 ;
        RECT 1554.530 0.350 1562.430 4.280 ;
        RECT 1563.270 0.350 1571.170 4.280 ;
        RECT 1572.010 0.350 1579.910 4.280 ;
        RECT 1580.750 0.350 1588.650 4.280 ;
        RECT 1589.490 0.350 1597.390 4.280 ;
        RECT 1598.230 0.350 1606.130 4.280 ;
        RECT 1606.970 0.350 1614.870 4.280 ;
        RECT 1615.710 0.350 1623.610 4.280 ;
        RECT 1624.450 0.350 1632.350 4.280 ;
        RECT 1633.190 0.350 1641.090 4.280 ;
        RECT 1641.930 0.350 1649.830 4.280 ;
        RECT 1650.670 0.350 1658.570 4.280 ;
        RECT 1659.410 0.350 1667.310 4.280 ;
        RECT 1668.150 0.350 1676.050 4.280 ;
        RECT 1676.890 0.350 1684.790 4.280 ;
        RECT 1685.630 0.350 1693.530 4.280 ;
        RECT 1694.370 0.350 1702.270 4.280 ;
        RECT 1703.110 0.350 1711.010 4.280 ;
        RECT 1711.850 0.350 1719.750 4.280 ;
        RECT 1720.590 0.350 1728.490 4.280 ;
        RECT 1729.330 0.350 1737.230 4.280 ;
        RECT 1738.070 0.350 1745.970 4.280 ;
        RECT 1746.810 0.350 1754.710 4.280 ;
        RECT 1755.550 0.350 1763.450 4.280 ;
        RECT 1764.290 0.350 1772.190 4.280 ;
        RECT 1773.030 0.350 1780.930 4.280 ;
        RECT 1781.770 0.350 1789.670 4.280 ;
        RECT 1790.510 0.350 1798.410 4.280 ;
        RECT 1799.250 0.350 1807.150 4.280 ;
        RECT 1807.990 0.350 1815.890 4.280 ;
        RECT 1816.730 0.350 1824.630 4.280 ;
        RECT 1825.470 0.350 1833.370 4.280 ;
        RECT 1834.210 0.350 1842.110 4.280 ;
        RECT 1842.950 0.350 1850.850 4.280 ;
        RECT 1851.690 0.350 1859.590 4.280 ;
        RECT 1860.430 0.350 1868.330 4.280 ;
        RECT 1869.170 0.350 1877.070 4.280 ;
        RECT 1877.910 0.350 1885.810 4.280 ;
        RECT 1886.650 0.350 1894.550 4.280 ;
        RECT 1895.390 0.350 1903.290 4.280 ;
        RECT 1904.130 0.350 1912.030 4.280 ;
        RECT 1912.870 0.350 1920.770 4.280 ;
        RECT 1921.610 0.350 1929.510 4.280 ;
        RECT 1930.350 0.350 1938.250 4.280 ;
        RECT 1939.090 0.350 1946.990 4.280 ;
        RECT 1947.830 0.350 1955.730 4.280 ;
        RECT 1956.570 0.350 1964.470 4.280 ;
        RECT 1965.310 0.350 1973.210 4.280 ;
        RECT 1974.050 0.350 1981.950 4.280 ;
        RECT 1982.790 0.350 1990.690 4.280 ;
        RECT 1991.530 0.350 1999.430 4.280 ;
        RECT 2000.270 0.350 2008.170 4.280 ;
        RECT 2009.010 0.350 2016.910 4.280 ;
        RECT 2017.750 0.350 2025.650 4.280 ;
        RECT 2026.490 0.350 2034.390 4.280 ;
        RECT 2035.230 0.350 2043.130 4.280 ;
        RECT 2043.970 0.350 2051.870 4.280 ;
        RECT 2052.710 0.350 2060.610 4.280 ;
        RECT 2061.450 0.350 2069.350 4.280 ;
        RECT 2070.190 0.350 2078.090 4.280 ;
        RECT 2078.930 0.350 2086.830 4.280 ;
        RECT 2087.670 0.350 2095.570 4.280 ;
        RECT 2096.410 0.350 2104.310 4.280 ;
        RECT 2105.150 0.350 2113.050 4.280 ;
        RECT 2113.890 0.350 2121.790 4.280 ;
        RECT 2122.630 0.350 2130.530 4.280 ;
        RECT 2131.370 0.350 2139.270 4.280 ;
        RECT 2140.110 0.350 2148.010 4.280 ;
        RECT 2148.850 0.350 2156.750 4.280 ;
        RECT 2157.590 0.350 2196.860 4.280 ;
      LAYER met3 ;
        RECT 4.000 721.840 2196.000 796.785 ;
        RECT 4.000 720.440 2195.600 721.840 ;
        RECT 4.000 719.120 2196.000 720.440 ;
        RECT 4.000 717.720 2195.600 719.120 ;
        RECT 4.000 716.400 2196.000 717.720 ;
        RECT 4.400 715.000 2195.600 716.400 ;
        RECT 4.000 713.680 2196.000 715.000 ;
        RECT 4.400 712.280 2195.600 713.680 ;
        RECT 4.000 710.960 2196.000 712.280 ;
        RECT 4.400 709.560 2195.600 710.960 ;
        RECT 4.000 708.240 2196.000 709.560 ;
        RECT 4.400 706.840 2195.600 708.240 ;
        RECT 4.000 705.520 2196.000 706.840 ;
        RECT 4.400 704.120 2195.600 705.520 ;
        RECT 4.000 702.800 2196.000 704.120 ;
        RECT 4.400 701.400 2195.600 702.800 ;
        RECT 4.000 700.080 2196.000 701.400 ;
        RECT 4.400 698.680 2195.600 700.080 ;
        RECT 4.000 697.360 2196.000 698.680 ;
        RECT 4.400 695.960 2195.600 697.360 ;
        RECT 4.000 694.640 2196.000 695.960 ;
        RECT 4.400 693.240 2195.600 694.640 ;
        RECT 4.000 691.920 2196.000 693.240 ;
        RECT 4.400 690.520 2195.600 691.920 ;
        RECT 4.000 689.200 2196.000 690.520 ;
        RECT 4.400 687.800 2195.600 689.200 ;
        RECT 4.000 686.480 2196.000 687.800 ;
        RECT 4.400 685.080 2195.600 686.480 ;
        RECT 4.000 683.760 2196.000 685.080 ;
        RECT 4.400 682.360 2195.600 683.760 ;
        RECT 4.000 681.040 2196.000 682.360 ;
        RECT 4.400 679.640 2195.600 681.040 ;
        RECT 4.000 678.320 2196.000 679.640 ;
        RECT 4.400 676.920 2195.600 678.320 ;
        RECT 4.000 675.600 2196.000 676.920 ;
        RECT 4.400 674.200 2195.600 675.600 ;
        RECT 4.000 672.880 2196.000 674.200 ;
        RECT 4.400 671.480 2195.600 672.880 ;
        RECT 4.000 670.160 2196.000 671.480 ;
        RECT 4.400 668.760 2195.600 670.160 ;
        RECT 4.000 667.440 2196.000 668.760 ;
        RECT 4.400 666.040 2195.600 667.440 ;
        RECT 4.000 664.720 2196.000 666.040 ;
        RECT 4.400 663.320 2195.600 664.720 ;
        RECT 4.000 662.000 2196.000 663.320 ;
        RECT 4.400 660.600 2195.600 662.000 ;
        RECT 4.000 659.280 2196.000 660.600 ;
        RECT 4.400 657.880 2195.600 659.280 ;
        RECT 4.000 656.560 2196.000 657.880 ;
        RECT 4.400 655.160 2195.600 656.560 ;
        RECT 4.000 653.840 2196.000 655.160 ;
        RECT 4.400 652.440 2195.600 653.840 ;
        RECT 4.000 651.120 2196.000 652.440 ;
        RECT 4.400 649.720 2195.600 651.120 ;
        RECT 4.000 648.400 2196.000 649.720 ;
        RECT 4.400 647.000 2195.600 648.400 ;
        RECT 4.000 645.680 2196.000 647.000 ;
        RECT 4.400 644.280 2195.600 645.680 ;
        RECT 4.000 642.960 2196.000 644.280 ;
        RECT 4.400 641.560 2195.600 642.960 ;
        RECT 4.000 640.240 2196.000 641.560 ;
        RECT 4.400 638.840 2195.600 640.240 ;
        RECT 4.000 637.520 2196.000 638.840 ;
        RECT 4.400 636.120 2195.600 637.520 ;
        RECT 4.000 634.800 2196.000 636.120 ;
        RECT 4.400 633.400 2195.600 634.800 ;
        RECT 4.000 632.080 2196.000 633.400 ;
        RECT 4.400 630.680 2195.600 632.080 ;
        RECT 4.000 629.360 2196.000 630.680 ;
        RECT 4.400 627.960 2195.600 629.360 ;
        RECT 4.000 626.640 2196.000 627.960 ;
        RECT 4.400 625.240 2195.600 626.640 ;
        RECT 4.000 623.920 2196.000 625.240 ;
        RECT 4.400 622.520 2195.600 623.920 ;
        RECT 4.000 621.200 2196.000 622.520 ;
        RECT 4.400 619.800 2195.600 621.200 ;
        RECT 4.000 618.480 2196.000 619.800 ;
        RECT 4.400 617.080 2195.600 618.480 ;
        RECT 4.000 615.760 2196.000 617.080 ;
        RECT 4.400 614.360 2195.600 615.760 ;
        RECT 4.000 613.040 2196.000 614.360 ;
        RECT 4.400 611.640 2195.600 613.040 ;
        RECT 4.000 610.320 2196.000 611.640 ;
        RECT 4.400 608.920 2195.600 610.320 ;
        RECT 4.000 607.600 2196.000 608.920 ;
        RECT 4.400 606.200 2195.600 607.600 ;
        RECT 4.000 604.880 2196.000 606.200 ;
        RECT 4.400 603.480 2195.600 604.880 ;
        RECT 4.000 602.160 2196.000 603.480 ;
        RECT 4.400 600.760 2195.600 602.160 ;
        RECT 4.000 599.440 2196.000 600.760 ;
        RECT 4.400 598.040 2195.600 599.440 ;
        RECT 4.000 596.720 2196.000 598.040 ;
        RECT 4.400 595.320 2195.600 596.720 ;
        RECT 4.000 594.000 2196.000 595.320 ;
        RECT 4.400 592.600 2195.600 594.000 ;
        RECT 4.000 591.280 2196.000 592.600 ;
        RECT 4.400 589.880 2195.600 591.280 ;
        RECT 4.000 588.560 2196.000 589.880 ;
        RECT 4.400 587.160 2195.600 588.560 ;
        RECT 4.000 585.840 2196.000 587.160 ;
        RECT 4.400 584.440 2195.600 585.840 ;
        RECT 4.000 583.120 2196.000 584.440 ;
        RECT 4.400 581.720 2195.600 583.120 ;
        RECT 4.000 580.400 2196.000 581.720 ;
        RECT 4.400 579.000 2195.600 580.400 ;
        RECT 4.000 577.680 2196.000 579.000 ;
        RECT 4.400 576.280 2195.600 577.680 ;
        RECT 4.000 574.960 2196.000 576.280 ;
        RECT 4.400 573.560 2195.600 574.960 ;
        RECT 4.000 572.240 2196.000 573.560 ;
        RECT 4.400 570.840 2195.600 572.240 ;
        RECT 4.000 569.520 2196.000 570.840 ;
        RECT 4.400 568.120 2195.600 569.520 ;
        RECT 4.000 566.800 2196.000 568.120 ;
        RECT 4.400 565.400 2195.600 566.800 ;
        RECT 4.000 564.080 2196.000 565.400 ;
        RECT 4.400 562.680 2195.600 564.080 ;
        RECT 4.000 561.360 2196.000 562.680 ;
        RECT 4.400 559.960 2195.600 561.360 ;
        RECT 4.000 558.640 2196.000 559.960 ;
        RECT 4.400 557.240 2195.600 558.640 ;
        RECT 4.000 555.920 2196.000 557.240 ;
        RECT 4.400 554.520 2195.600 555.920 ;
        RECT 4.000 553.200 2196.000 554.520 ;
        RECT 4.400 551.800 2195.600 553.200 ;
        RECT 4.000 550.480 2196.000 551.800 ;
        RECT 4.400 549.080 2195.600 550.480 ;
        RECT 4.000 547.760 2196.000 549.080 ;
        RECT 4.400 546.360 2195.600 547.760 ;
        RECT 4.000 545.040 2196.000 546.360 ;
        RECT 4.400 543.640 2195.600 545.040 ;
        RECT 4.000 542.320 2196.000 543.640 ;
        RECT 4.400 540.920 2195.600 542.320 ;
        RECT 4.000 539.600 2196.000 540.920 ;
        RECT 4.400 538.200 2195.600 539.600 ;
        RECT 4.000 536.880 2196.000 538.200 ;
        RECT 4.400 535.480 2195.600 536.880 ;
        RECT 4.000 534.160 2196.000 535.480 ;
        RECT 4.400 532.760 2195.600 534.160 ;
        RECT 4.000 531.440 2196.000 532.760 ;
        RECT 4.400 530.040 2195.600 531.440 ;
        RECT 4.000 528.720 2196.000 530.040 ;
        RECT 4.400 527.320 2195.600 528.720 ;
        RECT 4.000 526.000 2196.000 527.320 ;
        RECT 4.400 524.600 2195.600 526.000 ;
        RECT 4.000 523.280 2196.000 524.600 ;
        RECT 4.400 521.880 2195.600 523.280 ;
        RECT 4.000 520.560 2196.000 521.880 ;
        RECT 4.400 519.160 2195.600 520.560 ;
        RECT 4.000 517.840 2196.000 519.160 ;
        RECT 4.400 516.440 2195.600 517.840 ;
        RECT 4.000 515.120 2196.000 516.440 ;
        RECT 4.400 513.720 2195.600 515.120 ;
        RECT 4.000 512.400 2196.000 513.720 ;
        RECT 4.400 511.000 2195.600 512.400 ;
        RECT 4.000 509.680 2196.000 511.000 ;
        RECT 4.400 508.280 2195.600 509.680 ;
        RECT 4.000 506.960 2196.000 508.280 ;
        RECT 4.400 505.560 2195.600 506.960 ;
        RECT 4.000 504.240 2196.000 505.560 ;
        RECT 4.400 502.840 2195.600 504.240 ;
        RECT 4.000 501.520 2196.000 502.840 ;
        RECT 4.400 500.120 2195.600 501.520 ;
        RECT 4.000 498.800 2196.000 500.120 ;
        RECT 4.400 497.400 2195.600 498.800 ;
        RECT 4.000 496.080 2196.000 497.400 ;
        RECT 4.400 494.680 2195.600 496.080 ;
        RECT 4.000 493.360 2196.000 494.680 ;
        RECT 4.400 491.960 2195.600 493.360 ;
        RECT 4.000 490.640 2196.000 491.960 ;
        RECT 4.400 489.240 2195.600 490.640 ;
        RECT 4.000 487.920 2196.000 489.240 ;
        RECT 4.400 486.520 2195.600 487.920 ;
        RECT 4.000 485.200 2196.000 486.520 ;
        RECT 4.400 483.800 2195.600 485.200 ;
        RECT 4.000 482.480 2196.000 483.800 ;
        RECT 4.400 481.080 2195.600 482.480 ;
        RECT 4.000 479.760 2196.000 481.080 ;
        RECT 4.400 478.360 2195.600 479.760 ;
        RECT 4.000 477.040 2196.000 478.360 ;
        RECT 4.400 475.640 2195.600 477.040 ;
        RECT 4.000 474.320 2196.000 475.640 ;
        RECT 4.400 472.920 2195.600 474.320 ;
        RECT 4.000 471.600 2196.000 472.920 ;
        RECT 4.400 470.200 2195.600 471.600 ;
        RECT 4.000 468.880 2196.000 470.200 ;
        RECT 4.400 467.480 2195.600 468.880 ;
        RECT 4.000 466.160 2196.000 467.480 ;
        RECT 4.400 464.760 2195.600 466.160 ;
        RECT 4.000 463.440 2196.000 464.760 ;
        RECT 4.400 462.040 2195.600 463.440 ;
        RECT 4.000 460.720 2196.000 462.040 ;
        RECT 4.400 459.320 2195.600 460.720 ;
        RECT 4.000 458.000 2196.000 459.320 ;
        RECT 4.400 456.600 2195.600 458.000 ;
        RECT 4.000 455.280 2196.000 456.600 ;
        RECT 4.400 453.880 2195.600 455.280 ;
        RECT 4.000 452.560 2196.000 453.880 ;
        RECT 4.400 451.160 2195.600 452.560 ;
        RECT 4.000 449.840 2196.000 451.160 ;
        RECT 4.400 448.440 2195.600 449.840 ;
        RECT 4.000 447.120 2196.000 448.440 ;
        RECT 4.400 445.720 2195.600 447.120 ;
        RECT 4.000 444.400 2196.000 445.720 ;
        RECT 4.400 443.000 2195.600 444.400 ;
        RECT 4.000 441.680 2196.000 443.000 ;
        RECT 4.400 440.280 2195.600 441.680 ;
        RECT 4.000 438.960 2196.000 440.280 ;
        RECT 4.400 437.560 2195.600 438.960 ;
        RECT 4.000 436.240 2196.000 437.560 ;
        RECT 4.400 434.840 2195.600 436.240 ;
        RECT 4.000 433.520 2196.000 434.840 ;
        RECT 4.400 432.120 2195.600 433.520 ;
        RECT 4.000 430.800 2196.000 432.120 ;
        RECT 4.400 429.400 2195.600 430.800 ;
        RECT 4.000 428.080 2196.000 429.400 ;
        RECT 4.400 426.680 2195.600 428.080 ;
        RECT 4.000 425.360 2196.000 426.680 ;
        RECT 4.400 423.960 2195.600 425.360 ;
        RECT 4.000 422.640 2196.000 423.960 ;
        RECT 4.400 421.240 2195.600 422.640 ;
        RECT 4.000 419.920 2196.000 421.240 ;
        RECT 4.400 418.520 2195.600 419.920 ;
        RECT 4.000 417.200 2196.000 418.520 ;
        RECT 4.400 415.800 2195.600 417.200 ;
        RECT 4.000 414.480 2196.000 415.800 ;
        RECT 4.400 413.080 2195.600 414.480 ;
        RECT 4.000 411.760 2196.000 413.080 ;
        RECT 4.400 410.360 2195.600 411.760 ;
        RECT 4.000 409.040 2196.000 410.360 ;
        RECT 4.400 407.640 2195.600 409.040 ;
        RECT 4.000 406.320 2196.000 407.640 ;
        RECT 4.400 404.920 2195.600 406.320 ;
        RECT 4.000 403.600 2196.000 404.920 ;
        RECT 4.400 402.200 2195.600 403.600 ;
        RECT 4.000 400.880 2196.000 402.200 ;
        RECT 4.400 399.480 2195.600 400.880 ;
        RECT 4.000 398.160 2196.000 399.480 ;
        RECT 4.400 396.760 2195.600 398.160 ;
        RECT 4.000 395.440 2196.000 396.760 ;
        RECT 4.400 394.040 2195.600 395.440 ;
        RECT 4.000 392.720 2196.000 394.040 ;
        RECT 4.400 391.320 2195.600 392.720 ;
        RECT 4.000 390.000 2196.000 391.320 ;
        RECT 4.400 388.600 2195.600 390.000 ;
        RECT 4.000 387.280 2196.000 388.600 ;
        RECT 4.400 385.880 2195.600 387.280 ;
        RECT 4.000 384.560 2196.000 385.880 ;
        RECT 4.400 383.160 2195.600 384.560 ;
        RECT 4.000 381.840 2196.000 383.160 ;
        RECT 4.400 380.440 2195.600 381.840 ;
        RECT 4.000 379.120 2196.000 380.440 ;
        RECT 4.400 377.720 2195.600 379.120 ;
        RECT 4.000 376.400 2196.000 377.720 ;
        RECT 4.400 375.000 2195.600 376.400 ;
        RECT 4.000 373.680 2196.000 375.000 ;
        RECT 4.400 372.280 2195.600 373.680 ;
        RECT 4.000 370.960 2196.000 372.280 ;
        RECT 4.400 369.560 2195.600 370.960 ;
        RECT 4.000 368.240 2196.000 369.560 ;
        RECT 4.400 366.840 2195.600 368.240 ;
        RECT 4.000 365.520 2196.000 366.840 ;
        RECT 4.400 364.120 2195.600 365.520 ;
        RECT 4.000 362.800 2196.000 364.120 ;
        RECT 4.400 361.400 2195.600 362.800 ;
        RECT 4.000 360.080 2196.000 361.400 ;
        RECT 4.400 358.680 2195.600 360.080 ;
        RECT 4.000 357.360 2196.000 358.680 ;
        RECT 4.400 355.960 2195.600 357.360 ;
        RECT 4.000 354.640 2196.000 355.960 ;
        RECT 4.400 353.240 2195.600 354.640 ;
        RECT 4.000 351.920 2196.000 353.240 ;
        RECT 4.400 350.520 2195.600 351.920 ;
        RECT 4.000 349.200 2196.000 350.520 ;
        RECT 4.400 347.800 2195.600 349.200 ;
        RECT 4.000 346.480 2196.000 347.800 ;
        RECT 4.400 345.080 2195.600 346.480 ;
        RECT 4.000 343.760 2196.000 345.080 ;
        RECT 4.400 342.360 2195.600 343.760 ;
        RECT 4.000 341.040 2196.000 342.360 ;
        RECT 4.400 339.640 2195.600 341.040 ;
        RECT 4.000 338.320 2196.000 339.640 ;
        RECT 4.400 336.920 2195.600 338.320 ;
        RECT 4.000 335.600 2196.000 336.920 ;
        RECT 4.400 334.200 2195.600 335.600 ;
        RECT 4.000 332.880 2196.000 334.200 ;
        RECT 4.400 331.480 2195.600 332.880 ;
        RECT 4.000 330.160 2196.000 331.480 ;
        RECT 4.400 328.760 2195.600 330.160 ;
        RECT 4.000 327.440 2196.000 328.760 ;
        RECT 4.400 326.040 2195.600 327.440 ;
        RECT 4.000 324.720 2196.000 326.040 ;
        RECT 4.400 323.320 2195.600 324.720 ;
        RECT 4.000 322.000 2196.000 323.320 ;
        RECT 4.400 320.600 2195.600 322.000 ;
        RECT 4.000 319.280 2196.000 320.600 ;
        RECT 4.400 317.880 2195.600 319.280 ;
        RECT 4.000 316.560 2196.000 317.880 ;
        RECT 4.400 315.160 2195.600 316.560 ;
        RECT 4.000 313.840 2196.000 315.160 ;
        RECT 4.400 312.440 2195.600 313.840 ;
        RECT 4.000 311.120 2196.000 312.440 ;
        RECT 4.400 309.720 2195.600 311.120 ;
        RECT 4.000 308.400 2196.000 309.720 ;
        RECT 4.400 307.000 2195.600 308.400 ;
        RECT 4.000 305.680 2196.000 307.000 ;
        RECT 4.400 304.280 2195.600 305.680 ;
        RECT 4.000 302.960 2196.000 304.280 ;
        RECT 4.400 301.560 2195.600 302.960 ;
        RECT 4.000 300.240 2196.000 301.560 ;
        RECT 4.400 298.840 2195.600 300.240 ;
        RECT 4.000 297.520 2196.000 298.840 ;
        RECT 4.400 296.120 2195.600 297.520 ;
        RECT 4.000 294.800 2196.000 296.120 ;
        RECT 4.400 293.400 2195.600 294.800 ;
        RECT 4.000 292.080 2196.000 293.400 ;
        RECT 4.400 290.680 2195.600 292.080 ;
        RECT 4.000 289.360 2196.000 290.680 ;
        RECT 4.400 287.960 2195.600 289.360 ;
        RECT 4.000 286.640 2196.000 287.960 ;
        RECT 4.400 285.240 2195.600 286.640 ;
        RECT 4.000 283.920 2196.000 285.240 ;
        RECT 4.400 282.520 2195.600 283.920 ;
        RECT 4.000 281.200 2196.000 282.520 ;
        RECT 4.400 279.800 2195.600 281.200 ;
        RECT 4.000 278.480 2196.000 279.800 ;
        RECT 4.400 277.080 2195.600 278.480 ;
        RECT 4.000 275.760 2196.000 277.080 ;
        RECT 4.400 274.360 2195.600 275.760 ;
        RECT 4.000 273.040 2196.000 274.360 ;
        RECT 4.400 271.640 2195.600 273.040 ;
        RECT 4.000 270.320 2196.000 271.640 ;
        RECT 4.400 268.920 2195.600 270.320 ;
        RECT 4.000 267.600 2196.000 268.920 ;
        RECT 4.400 266.200 2195.600 267.600 ;
        RECT 4.000 264.880 2196.000 266.200 ;
        RECT 4.400 263.480 2195.600 264.880 ;
        RECT 4.000 262.160 2196.000 263.480 ;
        RECT 4.400 260.760 2195.600 262.160 ;
        RECT 4.000 259.440 2196.000 260.760 ;
        RECT 4.400 258.040 2195.600 259.440 ;
        RECT 4.000 256.720 2196.000 258.040 ;
        RECT 4.400 255.320 2195.600 256.720 ;
        RECT 4.000 254.000 2196.000 255.320 ;
        RECT 4.400 252.600 2195.600 254.000 ;
        RECT 4.000 251.280 2196.000 252.600 ;
        RECT 4.400 249.880 2195.600 251.280 ;
        RECT 4.000 248.560 2196.000 249.880 ;
        RECT 4.400 247.160 2195.600 248.560 ;
        RECT 4.000 245.840 2196.000 247.160 ;
        RECT 4.400 244.440 2195.600 245.840 ;
        RECT 4.000 243.120 2196.000 244.440 ;
        RECT 4.400 241.720 2195.600 243.120 ;
        RECT 4.000 240.400 2196.000 241.720 ;
        RECT 4.400 239.000 2195.600 240.400 ;
        RECT 4.000 237.680 2196.000 239.000 ;
        RECT 4.400 236.280 2195.600 237.680 ;
        RECT 4.000 234.960 2196.000 236.280 ;
        RECT 4.400 233.560 2195.600 234.960 ;
        RECT 4.000 232.240 2196.000 233.560 ;
        RECT 4.400 230.840 2195.600 232.240 ;
        RECT 4.000 229.520 2196.000 230.840 ;
        RECT 4.400 228.120 2195.600 229.520 ;
        RECT 4.000 226.800 2196.000 228.120 ;
        RECT 4.400 225.400 2195.600 226.800 ;
        RECT 4.000 224.080 2196.000 225.400 ;
        RECT 4.400 222.680 2195.600 224.080 ;
        RECT 4.000 221.360 2196.000 222.680 ;
        RECT 4.400 219.960 2195.600 221.360 ;
        RECT 4.000 218.640 2196.000 219.960 ;
        RECT 4.400 217.240 2195.600 218.640 ;
        RECT 4.000 215.920 2196.000 217.240 ;
        RECT 4.400 214.520 2195.600 215.920 ;
        RECT 4.000 213.200 2196.000 214.520 ;
        RECT 4.400 211.800 2195.600 213.200 ;
        RECT 4.000 210.480 2196.000 211.800 ;
        RECT 4.400 209.080 2195.600 210.480 ;
        RECT 4.000 207.760 2196.000 209.080 ;
        RECT 4.400 206.360 2195.600 207.760 ;
        RECT 4.000 205.040 2196.000 206.360 ;
        RECT 4.400 203.640 2195.600 205.040 ;
        RECT 4.000 202.320 2196.000 203.640 ;
        RECT 4.400 200.920 2195.600 202.320 ;
        RECT 4.000 199.600 2196.000 200.920 ;
        RECT 4.400 198.200 2195.600 199.600 ;
        RECT 4.000 196.880 2196.000 198.200 ;
        RECT 4.400 195.480 2195.600 196.880 ;
        RECT 4.000 194.160 2196.000 195.480 ;
        RECT 4.400 192.760 2195.600 194.160 ;
        RECT 4.000 191.440 2196.000 192.760 ;
        RECT 4.400 190.040 2195.600 191.440 ;
        RECT 4.000 188.720 2196.000 190.040 ;
        RECT 4.400 187.320 2195.600 188.720 ;
        RECT 4.000 186.000 2196.000 187.320 ;
        RECT 4.400 184.600 2195.600 186.000 ;
        RECT 4.000 183.280 2196.000 184.600 ;
        RECT 4.400 181.880 2195.600 183.280 ;
        RECT 4.000 180.560 2196.000 181.880 ;
        RECT 4.400 179.160 2195.600 180.560 ;
        RECT 4.000 177.840 2196.000 179.160 ;
        RECT 4.400 176.440 2195.600 177.840 ;
        RECT 4.000 175.120 2196.000 176.440 ;
        RECT 4.400 173.720 2195.600 175.120 ;
        RECT 4.000 172.400 2196.000 173.720 ;
        RECT 4.400 171.000 2195.600 172.400 ;
        RECT 4.000 169.680 2196.000 171.000 ;
        RECT 4.400 168.280 2195.600 169.680 ;
        RECT 4.000 166.960 2196.000 168.280 ;
        RECT 4.400 165.560 2195.600 166.960 ;
        RECT 4.000 164.240 2196.000 165.560 ;
        RECT 4.400 162.840 2195.600 164.240 ;
        RECT 4.000 161.520 2196.000 162.840 ;
        RECT 4.400 160.120 2195.600 161.520 ;
        RECT 4.000 158.800 2196.000 160.120 ;
        RECT 4.400 157.400 2195.600 158.800 ;
        RECT 4.000 156.080 2196.000 157.400 ;
        RECT 4.400 154.680 2195.600 156.080 ;
        RECT 4.000 153.360 2196.000 154.680 ;
        RECT 4.400 151.960 2195.600 153.360 ;
        RECT 4.000 150.640 2196.000 151.960 ;
        RECT 4.400 149.240 2195.600 150.640 ;
        RECT 4.000 147.920 2196.000 149.240 ;
        RECT 4.400 146.520 2195.600 147.920 ;
        RECT 4.000 145.200 2196.000 146.520 ;
        RECT 4.400 143.800 2195.600 145.200 ;
        RECT 4.000 142.480 2196.000 143.800 ;
        RECT 4.400 141.080 2195.600 142.480 ;
        RECT 4.000 139.760 2196.000 141.080 ;
        RECT 4.400 138.360 2195.600 139.760 ;
        RECT 4.000 137.040 2196.000 138.360 ;
        RECT 4.400 135.640 2195.600 137.040 ;
        RECT 4.000 134.320 2196.000 135.640 ;
        RECT 4.400 132.920 2195.600 134.320 ;
        RECT 4.000 131.600 2196.000 132.920 ;
        RECT 4.400 130.200 2195.600 131.600 ;
        RECT 4.000 128.880 2196.000 130.200 ;
        RECT 4.400 127.480 2195.600 128.880 ;
        RECT 4.000 126.160 2196.000 127.480 ;
        RECT 4.400 124.760 2195.600 126.160 ;
        RECT 4.000 123.440 2196.000 124.760 ;
        RECT 4.400 122.040 2195.600 123.440 ;
        RECT 4.000 120.720 2196.000 122.040 ;
        RECT 4.400 119.320 2195.600 120.720 ;
        RECT 4.000 118.000 2196.000 119.320 ;
        RECT 4.400 116.600 2195.600 118.000 ;
        RECT 4.000 115.280 2196.000 116.600 ;
        RECT 4.400 113.880 2195.600 115.280 ;
        RECT 4.000 112.560 2196.000 113.880 ;
        RECT 4.400 111.160 2195.600 112.560 ;
        RECT 4.000 109.840 2196.000 111.160 ;
        RECT 4.400 108.440 2195.600 109.840 ;
        RECT 4.000 107.120 2196.000 108.440 ;
        RECT 4.400 105.720 2195.600 107.120 ;
        RECT 4.000 104.400 2196.000 105.720 ;
        RECT 4.400 103.000 2195.600 104.400 ;
        RECT 4.000 101.680 2196.000 103.000 ;
        RECT 4.400 100.280 2195.600 101.680 ;
        RECT 4.000 98.960 2196.000 100.280 ;
        RECT 4.400 97.560 2195.600 98.960 ;
        RECT 4.000 96.240 2196.000 97.560 ;
        RECT 4.400 94.840 2195.600 96.240 ;
        RECT 4.000 93.520 2196.000 94.840 ;
        RECT 4.400 92.120 2195.600 93.520 ;
        RECT 4.000 90.800 2196.000 92.120 ;
        RECT 4.400 89.400 2195.600 90.800 ;
        RECT 4.000 88.080 2196.000 89.400 ;
        RECT 4.400 86.680 2195.600 88.080 ;
        RECT 4.000 85.360 2196.000 86.680 ;
        RECT 4.400 83.960 2195.600 85.360 ;
        RECT 4.000 82.640 2196.000 83.960 ;
        RECT 4.400 81.240 2195.600 82.640 ;
        RECT 4.000 79.920 2196.000 81.240 ;
        RECT 4.000 78.520 2195.600 79.920 ;
        RECT 4.000 77.200 2196.000 78.520 ;
        RECT 4.000 75.800 2195.600 77.200 ;
        RECT 4.000 9.695 2196.000 75.800 ;
      LAYER met4 ;
        RECT 16.855 789.440 2186.545 796.785 ;
        RECT 16.855 15.135 20.640 789.440 ;
        RECT 23.040 15.135 97.440 789.440 ;
        RECT 99.840 15.135 174.240 789.440 ;
        RECT 176.640 15.135 251.040 789.440 ;
        RECT 253.440 15.135 327.840 789.440 ;
        RECT 330.240 15.135 404.640 789.440 ;
        RECT 407.040 15.135 481.440 789.440 ;
        RECT 483.840 15.135 558.240 789.440 ;
        RECT 560.640 15.135 635.040 789.440 ;
        RECT 637.440 15.135 711.840 789.440 ;
        RECT 714.240 15.135 788.640 789.440 ;
        RECT 791.040 15.135 865.440 789.440 ;
        RECT 867.840 15.135 942.240 789.440 ;
        RECT 944.640 15.135 1019.040 789.440 ;
        RECT 1021.440 15.135 1095.840 789.440 ;
        RECT 1098.240 15.135 1172.640 789.440 ;
        RECT 1175.040 15.135 1249.440 789.440 ;
        RECT 1251.840 15.135 1326.240 789.440 ;
        RECT 1328.640 15.135 1403.040 789.440 ;
        RECT 1405.440 15.135 1479.840 789.440 ;
        RECT 1482.240 15.135 1556.640 789.440 ;
        RECT 1559.040 15.135 1633.440 789.440 ;
        RECT 1635.840 15.135 1710.240 789.440 ;
        RECT 1712.640 15.135 1787.040 789.440 ;
        RECT 1789.440 15.135 1863.840 789.440 ;
        RECT 1866.240 15.135 1940.640 789.440 ;
        RECT 1943.040 15.135 2017.440 789.440 ;
        RECT 2019.840 15.135 2094.240 789.440 ;
        RECT 2096.640 15.135 2171.040 789.440 ;
        RECT 2173.440 15.135 2186.545 789.440 ;
  END
END vliw
END LIBRARY

