magic
tech sky130B
magscale 1 2
timestamp 1717251224
<< obsli1 >>
rect 1104 2159 418876 125681
<< obsm1 >>
rect 1104 1232 418876 127968
<< metal2 >>
rect 4250 127200 4306 128000
rect 5814 127200 5870 128000
rect 7378 127200 7434 128000
rect 8942 127200 8998 128000
rect 10506 127200 10562 128000
rect 12070 127200 12126 128000
rect 13634 127200 13690 128000
rect 15198 127200 15254 128000
rect 16762 127200 16818 128000
rect 18326 127200 18382 128000
rect 19890 127200 19946 128000
rect 21454 127200 21510 128000
rect 23018 127200 23074 128000
rect 24582 127200 24638 128000
rect 26146 127200 26202 128000
rect 27710 127200 27766 128000
rect 29274 127200 29330 128000
rect 30838 127200 30894 128000
rect 32402 127200 32458 128000
rect 33966 127200 34022 128000
rect 35530 127200 35586 128000
rect 37094 127200 37150 128000
rect 38658 127200 38714 128000
rect 40222 127200 40278 128000
rect 41786 127200 41842 128000
rect 43350 127200 43406 128000
rect 44914 127200 44970 128000
rect 46478 127200 46534 128000
rect 48042 127200 48098 128000
rect 49606 127200 49662 128000
rect 51170 127200 51226 128000
rect 52734 127200 52790 128000
rect 54298 127200 54354 128000
rect 55862 127200 55918 128000
rect 57426 127200 57482 128000
rect 58990 127200 59046 128000
rect 60554 127200 60610 128000
rect 62118 127200 62174 128000
rect 63682 127200 63738 128000
rect 65246 127200 65302 128000
rect 66810 127200 66866 128000
rect 68374 127200 68430 128000
rect 69938 127200 69994 128000
rect 71502 127200 71558 128000
rect 73066 127200 73122 128000
rect 74630 127200 74686 128000
rect 76194 127200 76250 128000
rect 77758 127200 77814 128000
rect 79322 127200 79378 128000
rect 80886 127200 80942 128000
rect 82450 127200 82506 128000
rect 84014 127200 84070 128000
rect 85578 127200 85634 128000
rect 87142 127200 87198 128000
rect 88706 127200 88762 128000
rect 90270 127200 90326 128000
rect 91834 127200 91890 128000
rect 93398 127200 93454 128000
rect 94962 127200 95018 128000
rect 96526 127200 96582 128000
rect 98090 127200 98146 128000
rect 99654 127200 99710 128000
rect 101218 127200 101274 128000
rect 102782 127200 102838 128000
rect 104346 127200 104402 128000
rect 105910 127200 105966 128000
rect 107474 127200 107530 128000
rect 109038 127200 109094 128000
rect 110602 127200 110658 128000
rect 112166 127200 112222 128000
rect 113730 127200 113786 128000
rect 115294 127200 115350 128000
rect 116858 127200 116914 128000
rect 118422 127200 118478 128000
rect 119986 127200 120042 128000
rect 121550 127200 121606 128000
rect 123114 127200 123170 128000
rect 124678 127200 124734 128000
rect 126242 127200 126298 128000
rect 127806 127200 127862 128000
rect 129370 127200 129426 128000
rect 130934 127200 130990 128000
rect 132498 127200 132554 128000
rect 134062 127200 134118 128000
rect 135626 127200 135682 128000
rect 137190 127200 137246 128000
rect 138754 127200 138810 128000
rect 140318 127200 140374 128000
rect 141882 127200 141938 128000
rect 143446 127200 143502 128000
rect 145010 127200 145066 128000
rect 146574 127200 146630 128000
rect 148138 127200 148194 128000
rect 149702 127200 149758 128000
rect 151266 127200 151322 128000
rect 152830 127200 152886 128000
rect 154394 127200 154450 128000
rect 155958 127200 156014 128000
rect 157522 127200 157578 128000
rect 159086 127200 159142 128000
rect 160650 127200 160706 128000
rect 162214 127200 162270 128000
rect 163778 127200 163834 128000
rect 165342 127200 165398 128000
rect 166906 127200 166962 128000
rect 168470 127200 168526 128000
rect 170034 127200 170090 128000
rect 171598 127200 171654 128000
rect 173162 127200 173218 128000
rect 174726 127200 174782 128000
rect 176290 127200 176346 128000
rect 177854 127200 177910 128000
rect 179418 127200 179474 128000
rect 180982 127200 181038 128000
rect 182546 127200 182602 128000
rect 184110 127200 184166 128000
rect 185674 127200 185730 128000
rect 187238 127200 187294 128000
rect 188802 127200 188858 128000
rect 190366 127200 190422 128000
rect 191930 127200 191986 128000
rect 193494 127200 193550 128000
rect 195058 127200 195114 128000
rect 196622 127200 196678 128000
rect 198186 127200 198242 128000
rect 199750 127200 199806 128000
rect 201314 127200 201370 128000
rect 202878 127200 202934 128000
rect 204442 127200 204498 128000
rect 206006 127200 206062 128000
rect 207570 127200 207626 128000
rect 209134 127200 209190 128000
rect 210698 127200 210754 128000
rect 212262 127200 212318 128000
rect 213826 127200 213882 128000
rect 215390 127200 215446 128000
rect 216954 127200 217010 128000
rect 218518 127200 218574 128000
rect 220082 127200 220138 128000
rect 221646 127200 221702 128000
rect 223210 127200 223266 128000
rect 224774 127200 224830 128000
rect 226338 127200 226394 128000
rect 227902 127200 227958 128000
rect 229466 127200 229522 128000
rect 231030 127200 231086 128000
rect 232594 127200 232650 128000
rect 234158 127200 234214 128000
rect 235722 127200 235778 128000
rect 237286 127200 237342 128000
rect 238850 127200 238906 128000
rect 240414 127200 240470 128000
rect 241978 127200 242034 128000
rect 243542 127200 243598 128000
rect 245106 127200 245162 128000
rect 246670 127200 246726 128000
rect 248234 127200 248290 128000
rect 249798 127200 249854 128000
rect 251362 127200 251418 128000
rect 252926 127200 252982 128000
rect 254490 127200 254546 128000
rect 256054 127200 256110 128000
rect 257618 127200 257674 128000
rect 259182 127200 259238 128000
rect 260746 127200 260802 128000
rect 262310 127200 262366 128000
rect 263874 127200 263930 128000
rect 265438 127200 265494 128000
rect 267002 127200 267058 128000
rect 268566 127200 268622 128000
rect 270130 127200 270186 128000
rect 271694 127200 271750 128000
rect 273258 127200 273314 128000
rect 274822 127200 274878 128000
rect 276386 127200 276442 128000
rect 277950 127200 278006 128000
rect 279514 127200 279570 128000
rect 281078 127200 281134 128000
rect 282642 127200 282698 128000
rect 284206 127200 284262 128000
rect 285770 127200 285826 128000
rect 287334 127200 287390 128000
rect 288898 127200 288954 128000
rect 290462 127200 290518 128000
rect 292026 127200 292082 128000
rect 293590 127200 293646 128000
rect 295154 127200 295210 128000
rect 296718 127200 296774 128000
rect 298282 127200 298338 128000
rect 299846 127200 299902 128000
rect 301410 127200 301466 128000
rect 302974 127200 303030 128000
rect 304538 127200 304594 128000
rect 306102 127200 306158 128000
rect 307666 127200 307722 128000
rect 309230 127200 309286 128000
rect 310794 127200 310850 128000
rect 312358 127200 312414 128000
rect 313922 127200 313978 128000
rect 315486 127200 315542 128000
rect 317050 127200 317106 128000
rect 318614 127200 318670 128000
rect 320178 127200 320234 128000
rect 321742 127200 321798 128000
rect 323306 127200 323362 128000
rect 324870 127200 324926 128000
rect 326434 127200 326490 128000
rect 327998 127200 328054 128000
rect 329562 127200 329618 128000
rect 331126 127200 331182 128000
rect 332690 127200 332746 128000
rect 334254 127200 334310 128000
rect 335818 127200 335874 128000
rect 337382 127200 337438 128000
rect 338946 127200 339002 128000
rect 340510 127200 340566 128000
rect 342074 127200 342130 128000
rect 343638 127200 343694 128000
rect 345202 127200 345258 128000
rect 346766 127200 346822 128000
rect 348330 127200 348386 128000
rect 349894 127200 349950 128000
rect 351458 127200 351514 128000
rect 353022 127200 353078 128000
rect 354586 127200 354642 128000
rect 356150 127200 356206 128000
rect 357714 127200 357770 128000
rect 359278 127200 359334 128000
rect 360842 127200 360898 128000
rect 362406 127200 362462 128000
rect 363970 127200 364026 128000
rect 365534 127200 365590 128000
rect 367098 127200 367154 128000
rect 368662 127200 368718 128000
rect 370226 127200 370282 128000
rect 371790 127200 371846 128000
rect 373354 127200 373410 128000
rect 374918 127200 374974 128000
rect 376482 127200 376538 128000
rect 378046 127200 378102 128000
rect 379610 127200 379666 128000
rect 381174 127200 381230 128000
rect 382738 127200 382794 128000
rect 384302 127200 384358 128000
rect 385866 127200 385922 128000
rect 387430 127200 387486 128000
rect 388994 127200 389050 128000
rect 390558 127200 390614 128000
rect 392122 127200 392178 128000
rect 393686 127200 393742 128000
rect 395250 127200 395306 128000
rect 396814 127200 396870 128000
rect 398378 127200 398434 128000
rect 399942 127200 399998 128000
rect 401506 127200 401562 128000
rect 403070 127200 403126 128000
rect 404634 127200 404690 128000
rect 406198 127200 406254 128000
rect 407762 127200 407818 128000
rect 409326 127200 409382 128000
rect 410890 127200 410946 128000
rect 412454 127200 412510 128000
rect 414018 127200 414074 128000
rect 415582 127200 415638 128000
rect 5446 0 5502 800
rect 9034 0 9090 800
rect 12622 0 12678 800
rect 16210 0 16266 800
rect 19798 0 19854 800
rect 23386 0 23442 800
rect 26974 0 27030 800
rect 30562 0 30618 800
rect 34150 0 34206 800
rect 37738 0 37794 800
rect 41326 0 41382 800
rect 44914 0 44970 800
rect 48502 0 48558 800
rect 52090 0 52146 800
rect 55678 0 55734 800
rect 59266 0 59322 800
rect 62854 0 62910 800
rect 66442 0 66498 800
rect 70030 0 70086 800
rect 73618 0 73674 800
rect 77206 0 77262 800
rect 80794 0 80850 800
rect 84382 0 84438 800
rect 87970 0 88026 800
rect 91558 0 91614 800
rect 95146 0 95202 800
rect 98734 0 98790 800
rect 102322 0 102378 800
rect 105910 0 105966 800
rect 109498 0 109554 800
rect 113086 0 113142 800
rect 116674 0 116730 800
rect 120262 0 120318 800
rect 123850 0 123906 800
rect 127438 0 127494 800
rect 131026 0 131082 800
rect 134614 0 134670 800
rect 138202 0 138258 800
rect 141790 0 141846 800
rect 145378 0 145434 800
rect 148966 0 149022 800
rect 152554 0 152610 800
rect 156142 0 156198 800
rect 159730 0 159786 800
rect 163318 0 163374 800
rect 166906 0 166962 800
rect 170494 0 170550 800
rect 174082 0 174138 800
rect 177670 0 177726 800
rect 181258 0 181314 800
rect 184846 0 184902 800
rect 188434 0 188490 800
rect 192022 0 192078 800
rect 195610 0 195666 800
rect 199198 0 199254 800
rect 202786 0 202842 800
rect 206374 0 206430 800
rect 209962 0 210018 800
rect 213550 0 213606 800
rect 217138 0 217194 800
rect 220726 0 220782 800
rect 224314 0 224370 800
rect 227902 0 227958 800
rect 231490 0 231546 800
rect 235078 0 235134 800
rect 238666 0 238722 800
rect 242254 0 242310 800
rect 245842 0 245898 800
rect 249430 0 249486 800
rect 253018 0 253074 800
rect 256606 0 256662 800
rect 260194 0 260250 800
rect 263782 0 263838 800
rect 267370 0 267426 800
rect 270958 0 271014 800
rect 274546 0 274602 800
rect 278134 0 278190 800
rect 281722 0 281778 800
rect 285310 0 285366 800
rect 288898 0 288954 800
rect 292486 0 292542 800
rect 296074 0 296130 800
rect 299662 0 299718 800
rect 303250 0 303306 800
rect 306838 0 306894 800
rect 310426 0 310482 800
rect 314014 0 314070 800
rect 317602 0 317658 800
rect 321190 0 321246 800
rect 324778 0 324834 800
rect 328366 0 328422 800
rect 331954 0 332010 800
rect 335542 0 335598 800
rect 339130 0 339186 800
rect 342718 0 342774 800
rect 346306 0 346362 800
rect 349894 0 349950 800
rect 353482 0 353538 800
rect 357070 0 357126 800
rect 360658 0 360714 800
rect 364246 0 364302 800
rect 367834 0 367890 800
rect 371422 0 371478 800
rect 375010 0 375066 800
rect 378598 0 378654 800
rect 382186 0 382242 800
rect 385774 0 385830 800
rect 389362 0 389418 800
rect 392950 0 393006 800
rect 396538 0 396594 800
rect 400126 0 400182 800
rect 403714 0 403770 800
rect 407302 0 407358 800
rect 410890 0 410946 800
rect 414478 0 414534 800
<< obsm2 >>
rect 2410 127144 4194 127974
rect 4362 127144 5758 127974
rect 5926 127144 7322 127974
rect 7490 127144 8886 127974
rect 9054 127144 10450 127974
rect 10618 127144 12014 127974
rect 12182 127144 13578 127974
rect 13746 127144 15142 127974
rect 15310 127144 16706 127974
rect 16874 127144 18270 127974
rect 18438 127144 19834 127974
rect 20002 127144 21398 127974
rect 21566 127144 22962 127974
rect 23130 127144 24526 127974
rect 24694 127144 26090 127974
rect 26258 127144 27654 127974
rect 27822 127144 29218 127974
rect 29386 127144 30782 127974
rect 30950 127144 32346 127974
rect 32514 127144 33910 127974
rect 34078 127144 35474 127974
rect 35642 127144 37038 127974
rect 37206 127144 38602 127974
rect 38770 127144 40166 127974
rect 40334 127144 41730 127974
rect 41898 127144 43294 127974
rect 43462 127144 44858 127974
rect 45026 127144 46422 127974
rect 46590 127144 47986 127974
rect 48154 127144 49550 127974
rect 49718 127144 51114 127974
rect 51282 127144 52678 127974
rect 52846 127144 54242 127974
rect 54410 127144 55806 127974
rect 55974 127144 57370 127974
rect 57538 127144 58934 127974
rect 59102 127144 60498 127974
rect 60666 127144 62062 127974
rect 62230 127144 63626 127974
rect 63794 127144 65190 127974
rect 65358 127144 66754 127974
rect 66922 127144 68318 127974
rect 68486 127144 69882 127974
rect 70050 127144 71446 127974
rect 71614 127144 73010 127974
rect 73178 127144 74574 127974
rect 74742 127144 76138 127974
rect 76306 127144 77702 127974
rect 77870 127144 79266 127974
rect 79434 127144 80830 127974
rect 80998 127144 82394 127974
rect 82562 127144 83958 127974
rect 84126 127144 85522 127974
rect 85690 127144 87086 127974
rect 87254 127144 88650 127974
rect 88818 127144 90214 127974
rect 90382 127144 91778 127974
rect 91946 127144 93342 127974
rect 93510 127144 94906 127974
rect 95074 127144 96470 127974
rect 96638 127144 98034 127974
rect 98202 127144 99598 127974
rect 99766 127144 101162 127974
rect 101330 127144 102726 127974
rect 102894 127144 104290 127974
rect 104458 127144 105854 127974
rect 106022 127144 107418 127974
rect 107586 127144 108982 127974
rect 109150 127144 110546 127974
rect 110714 127144 112110 127974
rect 112278 127144 113674 127974
rect 113842 127144 115238 127974
rect 115406 127144 116802 127974
rect 116970 127144 118366 127974
rect 118534 127144 119930 127974
rect 120098 127144 121494 127974
rect 121662 127144 123058 127974
rect 123226 127144 124622 127974
rect 124790 127144 126186 127974
rect 126354 127144 127750 127974
rect 127918 127144 129314 127974
rect 129482 127144 130878 127974
rect 131046 127144 132442 127974
rect 132610 127144 134006 127974
rect 134174 127144 135570 127974
rect 135738 127144 137134 127974
rect 137302 127144 138698 127974
rect 138866 127144 140262 127974
rect 140430 127144 141826 127974
rect 141994 127144 143390 127974
rect 143558 127144 144954 127974
rect 145122 127144 146518 127974
rect 146686 127144 148082 127974
rect 148250 127144 149646 127974
rect 149814 127144 151210 127974
rect 151378 127144 152774 127974
rect 152942 127144 154338 127974
rect 154506 127144 155902 127974
rect 156070 127144 157466 127974
rect 157634 127144 159030 127974
rect 159198 127144 160594 127974
rect 160762 127144 162158 127974
rect 162326 127144 163722 127974
rect 163890 127144 165286 127974
rect 165454 127144 166850 127974
rect 167018 127144 168414 127974
rect 168582 127144 169978 127974
rect 170146 127144 171542 127974
rect 171710 127144 173106 127974
rect 173274 127144 174670 127974
rect 174838 127144 176234 127974
rect 176402 127144 177798 127974
rect 177966 127144 179362 127974
rect 179530 127144 180926 127974
rect 181094 127144 182490 127974
rect 182658 127144 184054 127974
rect 184222 127144 185618 127974
rect 185786 127144 187182 127974
rect 187350 127144 188746 127974
rect 188914 127144 190310 127974
rect 190478 127144 191874 127974
rect 192042 127144 193438 127974
rect 193606 127144 195002 127974
rect 195170 127144 196566 127974
rect 196734 127144 198130 127974
rect 198298 127144 199694 127974
rect 199862 127144 201258 127974
rect 201426 127144 202822 127974
rect 202990 127144 204386 127974
rect 204554 127144 205950 127974
rect 206118 127144 207514 127974
rect 207682 127144 209078 127974
rect 209246 127144 210642 127974
rect 210810 127144 212206 127974
rect 212374 127144 213770 127974
rect 213938 127144 215334 127974
rect 215502 127144 216898 127974
rect 217066 127144 218462 127974
rect 218630 127144 220026 127974
rect 220194 127144 221590 127974
rect 221758 127144 223154 127974
rect 223322 127144 224718 127974
rect 224886 127144 226282 127974
rect 226450 127144 227846 127974
rect 228014 127144 229410 127974
rect 229578 127144 230974 127974
rect 231142 127144 232538 127974
rect 232706 127144 234102 127974
rect 234270 127144 235666 127974
rect 235834 127144 237230 127974
rect 237398 127144 238794 127974
rect 238962 127144 240358 127974
rect 240526 127144 241922 127974
rect 242090 127144 243486 127974
rect 243654 127144 245050 127974
rect 245218 127144 246614 127974
rect 246782 127144 248178 127974
rect 248346 127144 249742 127974
rect 249910 127144 251306 127974
rect 251474 127144 252870 127974
rect 253038 127144 254434 127974
rect 254602 127144 255998 127974
rect 256166 127144 257562 127974
rect 257730 127144 259126 127974
rect 259294 127144 260690 127974
rect 260858 127144 262254 127974
rect 262422 127144 263818 127974
rect 263986 127144 265382 127974
rect 265550 127144 266946 127974
rect 267114 127144 268510 127974
rect 268678 127144 270074 127974
rect 270242 127144 271638 127974
rect 271806 127144 273202 127974
rect 273370 127144 274766 127974
rect 274934 127144 276330 127974
rect 276498 127144 277894 127974
rect 278062 127144 279458 127974
rect 279626 127144 281022 127974
rect 281190 127144 282586 127974
rect 282754 127144 284150 127974
rect 284318 127144 285714 127974
rect 285882 127144 287278 127974
rect 287446 127144 288842 127974
rect 289010 127144 290406 127974
rect 290574 127144 291970 127974
rect 292138 127144 293534 127974
rect 293702 127144 295098 127974
rect 295266 127144 296662 127974
rect 296830 127144 298226 127974
rect 298394 127144 299790 127974
rect 299958 127144 301354 127974
rect 301522 127144 302918 127974
rect 303086 127144 304482 127974
rect 304650 127144 306046 127974
rect 306214 127144 307610 127974
rect 307778 127144 309174 127974
rect 309342 127144 310738 127974
rect 310906 127144 312302 127974
rect 312470 127144 313866 127974
rect 314034 127144 315430 127974
rect 315598 127144 316994 127974
rect 317162 127144 318558 127974
rect 318726 127144 320122 127974
rect 320290 127144 321686 127974
rect 321854 127144 323250 127974
rect 323418 127144 324814 127974
rect 324982 127144 326378 127974
rect 326546 127144 327942 127974
rect 328110 127144 329506 127974
rect 329674 127144 331070 127974
rect 331238 127144 332634 127974
rect 332802 127144 334198 127974
rect 334366 127144 335762 127974
rect 335930 127144 337326 127974
rect 337494 127144 338890 127974
rect 339058 127144 340454 127974
rect 340622 127144 342018 127974
rect 342186 127144 343582 127974
rect 343750 127144 345146 127974
rect 345314 127144 346710 127974
rect 346878 127144 348274 127974
rect 348442 127144 349838 127974
rect 350006 127144 351402 127974
rect 351570 127144 352966 127974
rect 353134 127144 354530 127974
rect 354698 127144 356094 127974
rect 356262 127144 357658 127974
rect 357826 127144 359222 127974
rect 359390 127144 360786 127974
rect 360954 127144 362350 127974
rect 362518 127144 363914 127974
rect 364082 127144 365478 127974
rect 365646 127144 367042 127974
rect 367210 127144 368606 127974
rect 368774 127144 370170 127974
rect 370338 127144 371734 127974
rect 371902 127144 373298 127974
rect 373466 127144 374862 127974
rect 375030 127144 376426 127974
rect 376594 127144 377990 127974
rect 378158 127144 379554 127974
rect 379722 127144 381118 127974
rect 381286 127144 382682 127974
rect 382850 127144 384246 127974
rect 384414 127144 385810 127974
rect 385978 127144 387374 127974
rect 387542 127144 388938 127974
rect 389106 127144 390502 127974
rect 390670 127144 392066 127974
rect 392234 127144 393630 127974
rect 393798 127144 395194 127974
rect 395362 127144 396758 127974
rect 396926 127144 398322 127974
rect 398490 127144 399886 127974
rect 400054 127144 401450 127974
rect 401618 127144 403014 127974
rect 403182 127144 404578 127974
rect 404746 127144 406142 127974
rect 406310 127144 407706 127974
rect 407874 127144 409270 127974
rect 409438 127144 410834 127974
rect 411002 127144 412398 127974
rect 412566 127144 413962 127974
rect 414130 127144 415526 127974
rect 415694 127144 418398 127974
rect 2410 856 418398 127144
rect 2410 303 5390 856
rect 5558 303 8978 856
rect 9146 303 12566 856
rect 12734 303 16154 856
rect 16322 303 19742 856
rect 19910 303 23330 856
rect 23498 303 26918 856
rect 27086 303 30506 856
rect 30674 303 34094 856
rect 34262 303 37682 856
rect 37850 303 41270 856
rect 41438 303 44858 856
rect 45026 303 48446 856
rect 48614 303 52034 856
rect 52202 303 55622 856
rect 55790 303 59210 856
rect 59378 303 62798 856
rect 62966 303 66386 856
rect 66554 303 69974 856
rect 70142 303 73562 856
rect 73730 303 77150 856
rect 77318 303 80738 856
rect 80906 303 84326 856
rect 84494 303 87914 856
rect 88082 303 91502 856
rect 91670 303 95090 856
rect 95258 303 98678 856
rect 98846 303 102266 856
rect 102434 303 105854 856
rect 106022 303 109442 856
rect 109610 303 113030 856
rect 113198 303 116618 856
rect 116786 303 120206 856
rect 120374 303 123794 856
rect 123962 303 127382 856
rect 127550 303 130970 856
rect 131138 303 134558 856
rect 134726 303 138146 856
rect 138314 303 141734 856
rect 141902 303 145322 856
rect 145490 303 148910 856
rect 149078 303 152498 856
rect 152666 303 156086 856
rect 156254 303 159674 856
rect 159842 303 163262 856
rect 163430 303 166850 856
rect 167018 303 170438 856
rect 170606 303 174026 856
rect 174194 303 177614 856
rect 177782 303 181202 856
rect 181370 303 184790 856
rect 184958 303 188378 856
rect 188546 303 191966 856
rect 192134 303 195554 856
rect 195722 303 199142 856
rect 199310 303 202730 856
rect 202898 303 206318 856
rect 206486 303 209906 856
rect 210074 303 213494 856
rect 213662 303 217082 856
rect 217250 303 220670 856
rect 220838 303 224258 856
rect 224426 303 227846 856
rect 228014 303 231434 856
rect 231602 303 235022 856
rect 235190 303 238610 856
rect 238778 303 242198 856
rect 242366 303 245786 856
rect 245954 303 249374 856
rect 249542 303 252962 856
rect 253130 303 256550 856
rect 256718 303 260138 856
rect 260306 303 263726 856
rect 263894 303 267314 856
rect 267482 303 270902 856
rect 271070 303 274490 856
rect 274658 303 278078 856
rect 278246 303 281666 856
rect 281834 303 285254 856
rect 285422 303 288842 856
rect 289010 303 292430 856
rect 292598 303 296018 856
rect 296186 303 299606 856
rect 299774 303 303194 856
rect 303362 303 306782 856
rect 306950 303 310370 856
rect 310538 303 313958 856
rect 314126 303 317546 856
rect 317714 303 321134 856
rect 321302 303 324722 856
rect 324890 303 328310 856
rect 328478 303 331898 856
rect 332066 303 335486 856
rect 335654 303 339074 856
rect 339242 303 342662 856
rect 342830 303 346250 856
rect 346418 303 349838 856
rect 350006 303 353426 856
rect 353594 303 357014 856
rect 357182 303 360602 856
rect 360770 303 364190 856
rect 364358 303 367778 856
rect 367946 303 371366 856
rect 371534 303 374954 856
rect 375122 303 378542 856
rect 378710 303 382130 856
rect 382298 303 385718 856
rect 385886 303 389306 856
rect 389474 303 392894 856
rect 393062 303 396482 856
rect 396650 303 400070 856
rect 400238 303 403658 856
rect 403826 303 407246 856
rect 407414 303 410834 856
rect 411002 303 414422 856
rect 414590 303 418398 856
<< metal3 >>
rect 0 127576 800 127696
rect 419200 127576 420000 127696
rect 0 127032 800 127152
rect 419200 127032 420000 127152
rect 0 126488 800 126608
rect 419200 126488 420000 126608
rect 0 125944 800 126064
rect 419200 125944 420000 126064
rect 0 125400 800 125520
rect 419200 125400 420000 125520
rect 0 124856 800 124976
rect 419200 124856 420000 124976
rect 0 124312 800 124432
rect 419200 124312 420000 124432
rect 0 123768 800 123888
rect 419200 123768 420000 123888
rect 0 123224 800 123344
rect 419200 123224 420000 123344
rect 0 122680 800 122800
rect 419200 122680 420000 122800
rect 0 122136 800 122256
rect 419200 122136 420000 122256
rect 0 121592 800 121712
rect 419200 121592 420000 121712
rect 0 121048 800 121168
rect 419200 121048 420000 121168
rect 0 120504 800 120624
rect 419200 120504 420000 120624
rect 0 119960 800 120080
rect 419200 119960 420000 120080
rect 0 119416 800 119536
rect 419200 119416 420000 119536
rect 0 118872 800 118992
rect 419200 118872 420000 118992
rect 0 118328 800 118448
rect 419200 118328 420000 118448
rect 0 117784 800 117904
rect 419200 117784 420000 117904
rect 0 117240 800 117360
rect 419200 117240 420000 117360
rect 0 116696 800 116816
rect 419200 116696 420000 116816
rect 0 116152 800 116272
rect 419200 116152 420000 116272
rect 0 115608 800 115728
rect 419200 115608 420000 115728
rect 0 115064 800 115184
rect 419200 115064 420000 115184
rect 0 114520 800 114640
rect 419200 114520 420000 114640
rect 0 113976 800 114096
rect 419200 113976 420000 114096
rect 0 113432 800 113552
rect 419200 113432 420000 113552
rect 0 112888 800 113008
rect 419200 112888 420000 113008
rect 0 112344 800 112464
rect 419200 112344 420000 112464
rect 0 111800 800 111920
rect 419200 111800 420000 111920
rect 0 111256 800 111376
rect 419200 111256 420000 111376
rect 0 110712 800 110832
rect 419200 110712 420000 110832
rect 0 110168 800 110288
rect 419200 110168 420000 110288
rect 0 109624 800 109744
rect 419200 109624 420000 109744
rect 0 109080 800 109200
rect 419200 109080 420000 109200
rect 0 108536 800 108656
rect 419200 108536 420000 108656
rect 0 107992 800 108112
rect 419200 107992 420000 108112
rect 0 107448 800 107568
rect 419200 107448 420000 107568
rect 0 106904 800 107024
rect 419200 106904 420000 107024
rect 0 106360 800 106480
rect 419200 106360 420000 106480
rect 0 105816 800 105936
rect 419200 105816 420000 105936
rect 0 105272 800 105392
rect 419200 105272 420000 105392
rect 0 104728 800 104848
rect 419200 104728 420000 104848
rect 0 104184 800 104304
rect 419200 104184 420000 104304
rect 0 103640 800 103760
rect 419200 103640 420000 103760
rect 0 103096 800 103216
rect 419200 103096 420000 103216
rect 0 102552 800 102672
rect 419200 102552 420000 102672
rect 0 102008 800 102128
rect 419200 102008 420000 102128
rect 0 101464 800 101584
rect 419200 101464 420000 101584
rect 0 100920 800 101040
rect 419200 100920 420000 101040
rect 0 100376 800 100496
rect 419200 100376 420000 100496
rect 0 99832 800 99952
rect 419200 99832 420000 99952
rect 0 99288 800 99408
rect 419200 99288 420000 99408
rect 0 98744 800 98864
rect 419200 98744 420000 98864
rect 0 98200 800 98320
rect 419200 98200 420000 98320
rect 0 97656 800 97776
rect 419200 97656 420000 97776
rect 0 97112 800 97232
rect 419200 97112 420000 97232
rect 0 96568 800 96688
rect 419200 96568 420000 96688
rect 0 96024 800 96144
rect 419200 96024 420000 96144
rect 0 95480 800 95600
rect 419200 95480 420000 95600
rect 0 94936 800 95056
rect 419200 94936 420000 95056
rect 0 94392 800 94512
rect 419200 94392 420000 94512
rect 0 93848 800 93968
rect 419200 93848 420000 93968
rect 0 93304 800 93424
rect 419200 93304 420000 93424
rect 0 92760 800 92880
rect 419200 92760 420000 92880
rect 0 92216 800 92336
rect 419200 92216 420000 92336
rect 0 91672 800 91792
rect 419200 91672 420000 91792
rect 0 91128 800 91248
rect 419200 91128 420000 91248
rect 0 90584 800 90704
rect 419200 90584 420000 90704
rect 0 90040 800 90160
rect 419200 90040 420000 90160
rect 0 89496 800 89616
rect 419200 89496 420000 89616
rect 0 88952 800 89072
rect 419200 88952 420000 89072
rect 0 88408 800 88528
rect 419200 88408 420000 88528
rect 0 87864 800 87984
rect 419200 87864 420000 87984
rect 0 87320 800 87440
rect 419200 87320 420000 87440
rect 0 86776 800 86896
rect 419200 86776 420000 86896
rect 0 86232 800 86352
rect 419200 86232 420000 86352
rect 0 85688 800 85808
rect 419200 85688 420000 85808
rect 0 85144 800 85264
rect 419200 85144 420000 85264
rect 0 84600 800 84720
rect 419200 84600 420000 84720
rect 0 84056 800 84176
rect 419200 84056 420000 84176
rect 0 83512 800 83632
rect 419200 83512 420000 83632
rect 0 82968 800 83088
rect 419200 82968 420000 83088
rect 0 82424 800 82544
rect 419200 82424 420000 82544
rect 0 81880 800 82000
rect 419200 81880 420000 82000
rect 0 81336 800 81456
rect 419200 81336 420000 81456
rect 0 80792 800 80912
rect 419200 80792 420000 80912
rect 0 80248 800 80368
rect 419200 80248 420000 80368
rect 0 79704 800 79824
rect 419200 79704 420000 79824
rect 0 79160 800 79280
rect 419200 79160 420000 79280
rect 0 78616 800 78736
rect 419200 78616 420000 78736
rect 0 78072 800 78192
rect 419200 78072 420000 78192
rect 0 77528 800 77648
rect 419200 77528 420000 77648
rect 0 76984 800 77104
rect 419200 76984 420000 77104
rect 0 76440 800 76560
rect 419200 76440 420000 76560
rect 0 75896 800 76016
rect 419200 75896 420000 76016
rect 0 75352 800 75472
rect 419200 75352 420000 75472
rect 0 74808 800 74928
rect 419200 74808 420000 74928
rect 0 74264 800 74384
rect 419200 74264 420000 74384
rect 0 73720 800 73840
rect 419200 73720 420000 73840
rect 0 73176 800 73296
rect 419200 73176 420000 73296
rect 0 72632 800 72752
rect 419200 72632 420000 72752
rect 0 72088 800 72208
rect 419200 72088 420000 72208
rect 0 71544 800 71664
rect 419200 71544 420000 71664
rect 0 71000 800 71120
rect 419200 71000 420000 71120
rect 0 70456 800 70576
rect 419200 70456 420000 70576
rect 0 69912 800 70032
rect 419200 69912 420000 70032
rect 0 69368 800 69488
rect 419200 69368 420000 69488
rect 0 68824 800 68944
rect 419200 68824 420000 68944
rect 0 68280 800 68400
rect 419200 68280 420000 68400
rect 0 67736 800 67856
rect 419200 67736 420000 67856
rect 0 67192 800 67312
rect 419200 67192 420000 67312
rect 0 66648 800 66768
rect 419200 66648 420000 66768
rect 0 66104 800 66224
rect 419200 66104 420000 66224
rect 0 65560 800 65680
rect 419200 65560 420000 65680
rect 0 65016 800 65136
rect 419200 65016 420000 65136
rect 0 64472 800 64592
rect 419200 64472 420000 64592
rect 0 63928 800 64048
rect 419200 63928 420000 64048
rect 0 63384 800 63504
rect 419200 63384 420000 63504
rect 0 62840 800 62960
rect 419200 62840 420000 62960
rect 0 62296 800 62416
rect 419200 62296 420000 62416
rect 0 61752 800 61872
rect 419200 61752 420000 61872
rect 0 61208 800 61328
rect 419200 61208 420000 61328
rect 0 60664 800 60784
rect 419200 60664 420000 60784
rect 0 60120 800 60240
rect 419200 60120 420000 60240
rect 0 59576 800 59696
rect 419200 59576 420000 59696
rect 0 59032 800 59152
rect 419200 59032 420000 59152
rect 0 58488 800 58608
rect 419200 58488 420000 58608
rect 0 57944 800 58064
rect 419200 57944 420000 58064
rect 0 57400 800 57520
rect 419200 57400 420000 57520
rect 0 56856 800 56976
rect 419200 56856 420000 56976
rect 0 56312 800 56432
rect 419200 56312 420000 56432
rect 0 55768 800 55888
rect 419200 55768 420000 55888
rect 0 55224 800 55344
rect 419200 55224 420000 55344
rect 0 54680 800 54800
rect 419200 54680 420000 54800
rect 0 54136 800 54256
rect 419200 54136 420000 54256
rect 0 53592 800 53712
rect 419200 53592 420000 53712
rect 0 53048 800 53168
rect 419200 53048 420000 53168
rect 0 52504 800 52624
rect 419200 52504 420000 52624
rect 0 51960 800 52080
rect 419200 51960 420000 52080
rect 0 51416 800 51536
rect 419200 51416 420000 51536
rect 0 50872 800 50992
rect 419200 50872 420000 50992
rect 0 50328 800 50448
rect 419200 50328 420000 50448
rect 0 49784 800 49904
rect 419200 49784 420000 49904
rect 0 49240 800 49360
rect 419200 49240 420000 49360
rect 0 48696 800 48816
rect 419200 48696 420000 48816
rect 0 48152 800 48272
rect 419200 48152 420000 48272
rect 0 47608 800 47728
rect 419200 47608 420000 47728
rect 0 47064 800 47184
rect 419200 47064 420000 47184
rect 0 46520 800 46640
rect 419200 46520 420000 46640
rect 0 45976 800 46096
rect 419200 45976 420000 46096
rect 0 45432 800 45552
rect 419200 45432 420000 45552
rect 0 44888 800 45008
rect 419200 44888 420000 45008
rect 0 44344 800 44464
rect 419200 44344 420000 44464
rect 0 43800 800 43920
rect 419200 43800 420000 43920
rect 0 43256 800 43376
rect 419200 43256 420000 43376
rect 0 42712 800 42832
rect 419200 42712 420000 42832
rect 0 42168 800 42288
rect 419200 42168 420000 42288
rect 0 41624 800 41744
rect 419200 41624 420000 41744
rect 0 41080 800 41200
rect 419200 41080 420000 41200
rect 0 40536 800 40656
rect 419200 40536 420000 40656
rect 0 39992 800 40112
rect 419200 39992 420000 40112
rect 0 39448 800 39568
rect 419200 39448 420000 39568
rect 0 38904 800 39024
rect 419200 38904 420000 39024
rect 0 38360 800 38480
rect 419200 38360 420000 38480
rect 0 37816 800 37936
rect 419200 37816 420000 37936
rect 0 37272 800 37392
rect 419200 37272 420000 37392
rect 0 36728 800 36848
rect 419200 36728 420000 36848
rect 0 36184 800 36304
rect 419200 36184 420000 36304
rect 0 35640 800 35760
rect 419200 35640 420000 35760
rect 0 35096 800 35216
rect 419200 35096 420000 35216
rect 0 34552 800 34672
rect 419200 34552 420000 34672
rect 0 34008 800 34128
rect 419200 34008 420000 34128
rect 0 33464 800 33584
rect 419200 33464 420000 33584
rect 0 32920 800 33040
rect 419200 32920 420000 33040
rect 0 32376 800 32496
rect 419200 32376 420000 32496
rect 0 31832 800 31952
rect 419200 31832 420000 31952
rect 0 31288 800 31408
rect 419200 31288 420000 31408
rect 0 30744 800 30864
rect 419200 30744 420000 30864
rect 0 30200 800 30320
rect 419200 30200 420000 30320
rect 0 29656 800 29776
rect 419200 29656 420000 29776
rect 0 29112 800 29232
rect 419200 29112 420000 29232
rect 0 28568 800 28688
rect 419200 28568 420000 28688
rect 0 28024 800 28144
rect 419200 28024 420000 28144
rect 0 27480 800 27600
rect 419200 27480 420000 27600
rect 0 26936 800 27056
rect 419200 26936 420000 27056
rect 0 26392 800 26512
rect 419200 26392 420000 26512
rect 0 25848 800 25968
rect 419200 25848 420000 25968
rect 0 25304 800 25424
rect 419200 25304 420000 25424
rect 0 24760 800 24880
rect 419200 24760 420000 24880
rect 0 24216 800 24336
rect 419200 24216 420000 24336
rect 0 23672 800 23792
rect 419200 23672 420000 23792
rect 0 23128 800 23248
rect 419200 23128 420000 23248
rect 0 22584 800 22704
rect 419200 22584 420000 22704
rect 0 22040 800 22160
rect 419200 22040 420000 22160
rect 0 21496 800 21616
rect 419200 21496 420000 21616
rect 0 20952 800 21072
rect 419200 20952 420000 21072
rect 0 20408 800 20528
rect 419200 20408 420000 20528
rect 0 19864 800 19984
rect 419200 19864 420000 19984
rect 0 19320 800 19440
rect 419200 19320 420000 19440
rect 0 18776 800 18896
rect 419200 18776 420000 18896
rect 0 18232 800 18352
rect 419200 18232 420000 18352
rect 0 17688 800 17808
rect 419200 17688 420000 17808
rect 0 17144 800 17264
rect 419200 17144 420000 17264
rect 0 16600 800 16720
rect 419200 16600 420000 16720
rect 0 16056 800 16176
rect 419200 16056 420000 16176
rect 0 15512 800 15632
rect 419200 15512 420000 15632
rect 0 14968 800 15088
rect 419200 14968 420000 15088
rect 0 14424 800 14544
rect 419200 14424 420000 14544
rect 0 13880 800 14000
rect 419200 13880 420000 14000
rect 0 13336 800 13456
rect 419200 13336 420000 13456
rect 0 12792 800 12912
rect 419200 12792 420000 12912
rect 0 12248 800 12368
rect 419200 12248 420000 12368
rect 0 11704 800 11824
rect 419200 11704 420000 11824
rect 0 11160 800 11280
rect 419200 11160 420000 11280
rect 0 10616 800 10736
rect 419200 10616 420000 10736
rect 0 10072 800 10192
rect 419200 10072 420000 10192
rect 0 9528 800 9648
rect 419200 9528 420000 9648
rect 0 8984 800 9104
rect 419200 8984 420000 9104
rect 0 8440 800 8560
rect 419200 8440 420000 8560
rect 0 7896 800 8016
rect 419200 7896 420000 8016
rect 0 7352 800 7472
rect 419200 7352 420000 7472
rect 0 6808 800 6928
rect 419200 6808 420000 6928
rect 0 6264 800 6384
rect 419200 6264 420000 6384
rect 0 5720 800 5840
rect 419200 5720 420000 5840
rect 0 5176 800 5296
rect 419200 5176 420000 5296
rect 0 4632 800 4752
rect 419200 4632 420000 4752
rect 0 4088 800 4208
rect 419200 4088 420000 4208
rect 0 3544 800 3664
rect 419200 3544 420000 3664
rect 0 3000 800 3120
rect 419200 3000 420000 3120
rect 0 2456 800 2576
rect 419200 2456 420000 2576
rect 0 1912 800 2032
rect 419200 1912 420000 2032
rect 0 1368 800 1488
rect 419200 1368 420000 1488
rect 0 824 800 944
rect 419200 824 420000 944
rect 0 280 800 400
rect 419200 280 420000 400
<< obsm3 >>
rect 880 127496 419120 127669
rect 800 127232 419200 127496
rect 880 126952 419120 127232
rect 800 126688 419200 126952
rect 880 126408 419120 126688
rect 800 126144 419200 126408
rect 880 125864 419120 126144
rect 800 125600 419200 125864
rect 880 125320 419120 125600
rect 800 125056 419200 125320
rect 880 124776 419120 125056
rect 800 124512 419200 124776
rect 880 124232 419120 124512
rect 800 123968 419200 124232
rect 880 123688 419120 123968
rect 800 123424 419200 123688
rect 880 123144 419120 123424
rect 800 122880 419200 123144
rect 880 122600 419120 122880
rect 800 122336 419200 122600
rect 880 122056 419120 122336
rect 800 121792 419200 122056
rect 880 121512 419120 121792
rect 800 121248 419200 121512
rect 880 120968 419120 121248
rect 800 120704 419200 120968
rect 880 120424 419120 120704
rect 800 120160 419200 120424
rect 880 119880 419120 120160
rect 800 119616 419200 119880
rect 880 119336 419120 119616
rect 800 119072 419200 119336
rect 880 118792 419120 119072
rect 800 118528 419200 118792
rect 880 118248 419120 118528
rect 800 117984 419200 118248
rect 880 117704 419120 117984
rect 800 117440 419200 117704
rect 880 117160 419120 117440
rect 800 116896 419200 117160
rect 880 116616 419120 116896
rect 800 116352 419200 116616
rect 880 116072 419120 116352
rect 800 115808 419200 116072
rect 880 115528 419120 115808
rect 800 115264 419200 115528
rect 880 114984 419120 115264
rect 800 114720 419200 114984
rect 880 114440 419120 114720
rect 800 114176 419200 114440
rect 880 113896 419120 114176
rect 800 113632 419200 113896
rect 880 113352 419120 113632
rect 800 113088 419200 113352
rect 880 112808 419120 113088
rect 800 112544 419200 112808
rect 880 112264 419120 112544
rect 800 112000 419200 112264
rect 880 111720 419120 112000
rect 800 111456 419200 111720
rect 880 111176 419120 111456
rect 800 110912 419200 111176
rect 880 110632 419120 110912
rect 800 110368 419200 110632
rect 880 110088 419120 110368
rect 800 109824 419200 110088
rect 880 109544 419120 109824
rect 800 109280 419200 109544
rect 880 109000 419120 109280
rect 800 108736 419200 109000
rect 880 108456 419120 108736
rect 800 108192 419200 108456
rect 880 107912 419120 108192
rect 800 107648 419200 107912
rect 880 107368 419120 107648
rect 800 107104 419200 107368
rect 880 106824 419120 107104
rect 800 106560 419200 106824
rect 880 106280 419120 106560
rect 800 106016 419200 106280
rect 880 105736 419120 106016
rect 800 105472 419200 105736
rect 880 105192 419120 105472
rect 800 104928 419200 105192
rect 880 104648 419120 104928
rect 800 104384 419200 104648
rect 880 104104 419120 104384
rect 800 103840 419200 104104
rect 880 103560 419120 103840
rect 800 103296 419200 103560
rect 880 103016 419120 103296
rect 800 102752 419200 103016
rect 880 102472 419120 102752
rect 800 102208 419200 102472
rect 880 101928 419120 102208
rect 800 101664 419200 101928
rect 880 101384 419120 101664
rect 800 101120 419200 101384
rect 880 100840 419120 101120
rect 800 100576 419200 100840
rect 880 100296 419120 100576
rect 800 100032 419200 100296
rect 880 99752 419120 100032
rect 800 99488 419200 99752
rect 880 99208 419120 99488
rect 800 98944 419200 99208
rect 880 98664 419120 98944
rect 800 98400 419200 98664
rect 880 98120 419120 98400
rect 800 97856 419200 98120
rect 880 97576 419120 97856
rect 800 97312 419200 97576
rect 880 97032 419120 97312
rect 800 96768 419200 97032
rect 880 96488 419120 96768
rect 800 96224 419200 96488
rect 880 95944 419120 96224
rect 800 95680 419200 95944
rect 880 95400 419120 95680
rect 800 95136 419200 95400
rect 880 94856 419120 95136
rect 800 94592 419200 94856
rect 880 94312 419120 94592
rect 800 94048 419200 94312
rect 880 93768 419120 94048
rect 800 93504 419200 93768
rect 880 93224 419120 93504
rect 800 92960 419200 93224
rect 880 92680 419120 92960
rect 800 92416 419200 92680
rect 880 92136 419120 92416
rect 800 91872 419200 92136
rect 880 91592 419120 91872
rect 800 91328 419200 91592
rect 880 91048 419120 91328
rect 800 90784 419200 91048
rect 880 90504 419120 90784
rect 800 90240 419200 90504
rect 880 89960 419120 90240
rect 800 89696 419200 89960
rect 880 89416 419120 89696
rect 800 89152 419200 89416
rect 880 88872 419120 89152
rect 800 88608 419200 88872
rect 880 88328 419120 88608
rect 800 88064 419200 88328
rect 880 87784 419120 88064
rect 800 87520 419200 87784
rect 880 87240 419120 87520
rect 800 86976 419200 87240
rect 880 86696 419120 86976
rect 800 86432 419200 86696
rect 880 86152 419120 86432
rect 800 85888 419200 86152
rect 880 85608 419120 85888
rect 800 85344 419200 85608
rect 880 85064 419120 85344
rect 800 84800 419200 85064
rect 880 84520 419120 84800
rect 800 84256 419200 84520
rect 880 83976 419120 84256
rect 800 83712 419200 83976
rect 880 83432 419120 83712
rect 800 83168 419200 83432
rect 880 82888 419120 83168
rect 800 82624 419200 82888
rect 880 82344 419120 82624
rect 800 82080 419200 82344
rect 880 81800 419120 82080
rect 800 81536 419200 81800
rect 880 81256 419120 81536
rect 800 80992 419200 81256
rect 880 80712 419120 80992
rect 800 80448 419200 80712
rect 880 80168 419120 80448
rect 800 79904 419200 80168
rect 880 79624 419120 79904
rect 800 79360 419200 79624
rect 880 79080 419120 79360
rect 800 78816 419200 79080
rect 880 78536 419120 78816
rect 800 78272 419200 78536
rect 880 77992 419120 78272
rect 800 77728 419200 77992
rect 880 77448 419120 77728
rect 800 77184 419200 77448
rect 880 76904 419120 77184
rect 800 76640 419200 76904
rect 880 76360 419120 76640
rect 800 76096 419200 76360
rect 880 75816 419120 76096
rect 800 75552 419200 75816
rect 880 75272 419120 75552
rect 800 75008 419200 75272
rect 880 74728 419120 75008
rect 800 74464 419200 74728
rect 880 74184 419120 74464
rect 800 73920 419200 74184
rect 880 73640 419120 73920
rect 800 73376 419200 73640
rect 880 73096 419120 73376
rect 800 72832 419200 73096
rect 880 72552 419120 72832
rect 800 72288 419200 72552
rect 880 72008 419120 72288
rect 800 71744 419200 72008
rect 880 71464 419120 71744
rect 800 71200 419200 71464
rect 880 70920 419120 71200
rect 800 70656 419200 70920
rect 880 70376 419120 70656
rect 800 70112 419200 70376
rect 880 69832 419120 70112
rect 800 69568 419200 69832
rect 880 69288 419120 69568
rect 800 69024 419200 69288
rect 880 68744 419120 69024
rect 800 68480 419200 68744
rect 880 68200 419120 68480
rect 800 67936 419200 68200
rect 880 67656 419120 67936
rect 800 67392 419200 67656
rect 880 67112 419120 67392
rect 800 66848 419200 67112
rect 880 66568 419120 66848
rect 800 66304 419200 66568
rect 880 66024 419120 66304
rect 800 65760 419200 66024
rect 880 65480 419120 65760
rect 800 65216 419200 65480
rect 880 64936 419120 65216
rect 800 64672 419200 64936
rect 880 64392 419120 64672
rect 800 64128 419200 64392
rect 880 63848 419120 64128
rect 800 63584 419200 63848
rect 880 63304 419120 63584
rect 800 63040 419200 63304
rect 880 62760 419120 63040
rect 800 62496 419200 62760
rect 880 62216 419120 62496
rect 800 61952 419200 62216
rect 880 61672 419120 61952
rect 800 61408 419200 61672
rect 880 61128 419120 61408
rect 800 60864 419200 61128
rect 880 60584 419120 60864
rect 800 60320 419200 60584
rect 880 60040 419120 60320
rect 800 59776 419200 60040
rect 880 59496 419120 59776
rect 800 59232 419200 59496
rect 880 58952 419120 59232
rect 800 58688 419200 58952
rect 880 58408 419120 58688
rect 800 58144 419200 58408
rect 880 57864 419120 58144
rect 800 57600 419200 57864
rect 880 57320 419120 57600
rect 800 57056 419200 57320
rect 880 56776 419120 57056
rect 800 56512 419200 56776
rect 880 56232 419120 56512
rect 800 55968 419200 56232
rect 880 55688 419120 55968
rect 800 55424 419200 55688
rect 880 55144 419120 55424
rect 800 54880 419200 55144
rect 880 54600 419120 54880
rect 800 54336 419200 54600
rect 880 54056 419120 54336
rect 800 53792 419200 54056
rect 880 53512 419120 53792
rect 800 53248 419200 53512
rect 880 52968 419120 53248
rect 800 52704 419200 52968
rect 880 52424 419120 52704
rect 800 52160 419200 52424
rect 880 51880 419120 52160
rect 800 51616 419200 51880
rect 880 51336 419120 51616
rect 800 51072 419200 51336
rect 880 50792 419120 51072
rect 800 50528 419200 50792
rect 880 50248 419120 50528
rect 800 49984 419200 50248
rect 880 49704 419120 49984
rect 800 49440 419200 49704
rect 880 49160 419120 49440
rect 800 48896 419200 49160
rect 880 48616 419120 48896
rect 800 48352 419200 48616
rect 880 48072 419120 48352
rect 800 47808 419200 48072
rect 880 47528 419120 47808
rect 800 47264 419200 47528
rect 880 46984 419120 47264
rect 800 46720 419200 46984
rect 880 46440 419120 46720
rect 800 46176 419200 46440
rect 880 45896 419120 46176
rect 800 45632 419200 45896
rect 880 45352 419120 45632
rect 800 45088 419200 45352
rect 880 44808 419120 45088
rect 800 44544 419200 44808
rect 880 44264 419120 44544
rect 800 44000 419200 44264
rect 880 43720 419120 44000
rect 800 43456 419200 43720
rect 880 43176 419120 43456
rect 800 42912 419200 43176
rect 880 42632 419120 42912
rect 800 42368 419200 42632
rect 880 42088 419120 42368
rect 800 41824 419200 42088
rect 880 41544 419120 41824
rect 800 41280 419200 41544
rect 880 41000 419120 41280
rect 800 40736 419200 41000
rect 880 40456 419120 40736
rect 800 40192 419200 40456
rect 880 39912 419120 40192
rect 800 39648 419200 39912
rect 880 39368 419120 39648
rect 800 39104 419200 39368
rect 880 38824 419120 39104
rect 800 38560 419200 38824
rect 880 38280 419120 38560
rect 800 38016 419200 38280
rect 880 37736 419120 38016
rect 800 37472 419200 37736
rect 880 37192 419120 37472
rect 800 36928 419200 37192
rect 880 36648 419120 36928
rect 800 36384 419200 36648
rect 880 36104 419120 36384
rect 800 35840 419200 36104
rect 880 35560 419120 35840
rect 800 35296 419200 35560
rect 880 35016 419120 35296
rect 800 34752 419200 35016
rect 880 34472 419120 34752
rect 800 34208 419200 34472
rect 880 33928 419120 34208
rect 800 33664 419200 33928
rect 880 33384 419120 33664
rect 800 33120 419200 33384
rect 880 32840 419120 33120
rect 800 32576 419200 32840
rect 880 32296 419120 32576
rect 800 32032 419200 32296
rect 880 31752 419120 32032
rect 800 31488 419200 31752
rect 880 31208 419120 31488
rect 800 30944 419200 31208
rect 880 30664 419120 30944
rect 800 30400 419200 30664
rect 880 30120 419120 30400
rect 800 29856 419200 30120
rect 880 29576 419120 29856
rect 800 29312 419200 29576
rect 880 29032 419120 29312
rect 800 28768 419200 29032
rect 880 28488 419120 28768
rect 800 28224 419200 28488
rect 880 27944 419120 28224
rect 800 27680 419200 27944
rect 880 27400 419120 27680
rect 800 27136 419200 27400
rect 880 26856 419120 27136
rect 800 26592 419200 26856
rect 880 26312 419120 26592
rect 800 26048 419200 26312
rect 880 25768 419120 26048
rect 800 25504 419200 25768
rect 880 25224 419120 25504
rect 800 24960 419200 25224
rect 880 24680 419120 24960
rect 800 24416 419200 24680
rect 880 24136 419120 24416
rect 800 23872 419200 24136
rect 880 23592 419120 23872
rect 800 23328 419200 23592
rect 880 23048 419120 23328
rect 800 22784 419200 23048
rect 880 22504 419120 22784
rect 800 22240 419200 22504
rect 880 21960 419120 22240
rect 800 21696 419200 21960
rect 880 21416 419120 21696
rect 800 21152 419200 21416
rect 880 20872 419120 21152
rect 800 20608 419200 20872
rect 880 20328 419120 20608
rect 800 20064 419200 20328
rect 880 19784 419120 20064
rect 800 19520 419200 19784
rect 880 19240 419120 19520
rect 800 18976 419200 19240
rect 880 18696 419120 18976
rect 800 18432 419200 18696
rect 880 18152 419120 18432
rect 800 17888 419200 18152
rect 880 17608 419120 17888
rect 800 17344 419200 17608
rect 880 17064 419120 17344
rect 800 16800 419200 17064
rect 880 16520 419120 16800
rect 800 16256 419200 16520
rect 880 15976 419120 16256
rect 800 15712 419200 15976
rect 880 15432 419120 15712
rect 800 15168 419200 15432
rect 880 14888 419120 15168
rect 800 14624 419200 14888
rect 880 14344 419120 14624
rect 800 14080 419200 14344
rect 880 13800 419120 14080
rect 800 13536 419200 13800
rect 880 13256 419120 13536
rect 800 12992 419200 13256
rect 880 12712 419120 12992
rect 800 12448 419200 12712
rect 880 12168 419120 12448
rect 800 11904 419200 12168
rect 880 11624 419120 11904
rect 800 11360 419200 11624
rect 880 11080 419120 11360
rect 800 10816 419200 11080
rect 880 10536 419120 10816
rect 800 10272 419200 10536
rect 880 9992 419120 10272
rect 800 9728 419200 9992
rect 880 9448 419120 9728
rect 800 9184 419200 9448
rect 880 8904 419120 9184
rect 800 8640 419200 8904
rect 880 8360 419120 8640
rect 800 8096 419200 8360
rect 880 7816 419120 8096
rect 800 7552 419200 7816
rect 880 7272 419120 7552
rect 800 7008 419200 7272
rect 880 6728 419120 7008
rect 800 6464 419200 6728
rect 880 6184 419120 6464
rect 800 5920 419200 6184
rect 880 5640 419120 5920
rect 800 5376 419200 5640
rect 880 5096 419120 5376
rect 800 4832 419200 5096
rect 880 4552 419120 4832
rect 800 4288 419200 4552
rect 880 4008 419120 4288
rect 800 3744 419200 4008
rect 880 3464 419120 3744
rect 800 3200 419200 3464
rect 880 2920 419120 3200
rect 800 2656 419200 2920
rect 880 2376 419120 2656
rect 800 2112 419200 2376
rect 880 1832 419120 2112
rect 800 1568 419200 1832
rect 880 1288 419120 1568
rect 800 1024 419200 1288
rect 880 744 419120 1024
rect 800 480 419200 744
rect 880 307 419120 480
<< metal4 >>
rect 4208 2128 4528 125712
rect 19568 2128 19888 125712
rect 34928 2128 35248 125712
rect 50288 2128 50608 125712
rect 65648 2128 65968 125712
rect 81008 2128 81328 125712
rect 96368 2128 96688 125712
rect 111728 2128 112048 125712
rect 127088 2128 127408 125712
rect 142448 2128 142768 125712
rect 157808 2128 158128 125712
rect 173168 2128 173488 125712
rect 188528 2128 188848 125712
rect 203888 2128 204208 125712
rect 219248 2128 219568 125712
rect 234608 2128 234928 125712
rect 249968 2128 250288 125712
rect 265328 2128 265648 125712
rect 280688 2128 281008 125712
rect 296048 2128 296368 125712
rect 311408 2128 311728 125712
rect 326768 2128 327088 125712
rect 342128 2128 342448 125712
rect 357488 2128 357808 125712
rect 372848 2128 373168 125712
rect 388208 2128 388528 125712
rect 403568 2128 403888 125712
<< obsm4 >>
rect 70163 125792 416701 127669
rect 70163 2048 80928 125792
rect 81408 2048 96288 125792
rect 96768 2048 111648 125792
rect 112128 2048 127008 125792
rect 127488 2048 142368 125792
rect 142848 2048 157728 125792
rect 158208 2048 173088 125792
rect 173568 2048 188448 125792
rect 188928 2048 203808 125792
rect 204288 2048 219168 125792
rect 219648 2048 234528 125792
rect 235008 2048 249888 125792
rect 250368 2048 265248 125792
rect 265728 2048 280608 125792
rect 281088 2048 295968 125792
rect 296448 2048 311328 125792
rect 311808 2048 326688 125792
rect 327168 2048 342048 125792
rect 342528 2048 357408 125792
rect 357888 2048 372768 125792
rect 373248 2048 388128 125792
rect 388608 2048 403488 125792
rect 403968 2048 416701 125792
rect 70163 307 416701 2048
<< labels >>
rlabel metal2 s 5814 127200 5870 128000 6 curr_PC[0]
port 1 nsew signal output
rlabel metal2 s 21454 127200 21510 128000 6 curr_PC[10]
port 2 nsew signal output
rlabel metal2 s 23018 127200 23074 128000 6 curr_PC[11]
port 3 nsew signal output
rlabel metal2 s 24582 127200 24638 128000 6 curr_PC[12]
port 4 nsew signal output
rlabel metal2 s 26146 127200 26202 128000 6 curr_PC[13]
port 5 nsew signal output
rlabel metal2 s 27710 127200 27766 128000 6 curr_PC[14]
port 6 nsew signal output
rlabel metal2 s 29274 127200 29330 128000 6 curr_PC[15]
port 7 nsew signal output
rlabel metal2 s 30838 127200 30894 128000 6 curr_PC[16]
port 8 nsew signal output
rlabel metal2 s 32402 127200 32458 128000 6 curr_PC[17]
port 9 nsew signal output
rlabel metal2 s 33966 127200 34022 128000 6 curr_PC[18]
port 10 nsew signal output
rlabel metal2 s 35530 127200 35586 128000 6 curr_PC[19]
port 11 nsew signal output
rlabel metal2 s 7378 127200 7434 128000 6 curr_PC[1]
port 12 nsew signal output
rlabel metal2 s 37094 127200 37150 128000 6 curr_PC[20]
port 13 nsew signal output
rlabel metal2 s 38658 127200 38714 128000 6 curr_PC[21]
port 14 nsew signal output
rlabel metal2 s 40222 127200 40278 128000 6 curr_PC[22]
port 15 nsew signal output
rlabel metal2 s 41786 127200 41842 128000 6 curr_PC[23]
port 16 nsew signal output
rlabel metal2 s 43350 127200 43406 128000 6 curr_PC[24]
port 17 nsew signal output
rlabel metal2 s 44914 127200 44970 128000 6 curr_PC[25]
port 18 nsew signal output
rlabel metal2 s 46478 127200 46534 128000 6 curr_PC[26]
port 19 nsew signal output
rlabel metal2 s 48042 127200 48098 128000 6 curr_PC[27]
port 20 nsew signal output
rlabel metal2 s 8942 127200 8998 128000 6 curr_PC[2]
port 21 nsew signal output
rlabel metal2 s 10506 127200 10562 128000 6 curr_PC[3]
port 22 nsew signal output
rlabel metal2 s 12070 127200 12126 128000 6 curr_PC[4]
port 23 nsew signal output
rlabel metal2 s 13634 127200 13690 128000 6 curr_PC[5]
port 24 nsew signal output
rlabel metal2 s 15198 127200 15254 128000 6 curr_PC[6]
port 25 nsew signal output
rlabel metal2 s 16762 127200 16818 128000 6 curr_PC[7]
port 26 nsew signal output
rlabel metal2 s 18326 127200 18382 128000 6 curr_PC[8]
port 27 nsew signal output
rlabel metal2 s 19890 127200 19946 128000 6 curr_PC[9]
port 28 nsew signal output
rlabel metal2 s 400126 0 400182 800 6 custom_settings[0]
port 29 nsew signal input
rlabel metal2 s 403714 0 403770 800 6 custom_settings[1]
port 30 nsew signal input
rlabel metal2 s 407302 0 407358 800 6 custom_settings[2]
port 31 nsew signal input
rlabel metal2 s 410890 0 410946 800 6 custom_settings[3]
port 32 nsew signal input
rlabel metal2 s 414478 0 414534 800 6 custom_settings[4]
port 33 nsew signal input
rlabel metal2 s 118422 127200 118478 128000 6 dest_idx0[0]
port 34 nsew signal input
rlabel metal2 s 119986 127200 120042 128000 6 dest_idx0[1]
port 35 nsew signal input
rlabel metal2 s 121550 127200 121606 128000 6 dest_idx0[2]
port 36 nsew signal input
rlabel metal2 s 123114 127200 123170 128000 6 dest_idx0[3]
port 37 nsew signal input
rlabel metal2 s 124678 127200 124734 128000 6 dest_idx0[4]
port 38 nsew signal input
rlabel metal3 s 419200 24216 420000 24336 6 dest_idx1[0]
port 39 nsew signal input
rlabel metal3 s 419200 24760 420000 24880 6 dest_idx1[1]
port 40 nsew signal input
rlabel metal3 s 419200 25304 420000 25424 6 dest_idx1[2]
port 41 nsew signal input
rlabel metal3 s 419200 25848 420000 25968 6 dest_idx1[3]
port 42 nsew signal input
rlabel metal3 s 419200 26392 420000 26512 6 dest_idx1[4]
port 43 nsew signal input
rlabel metal3 s 0 24216 800 24336 6 dest_idx2[0]
port 44 nsew signal input
rlabel metal3 s 0 24760 800 24880 6 dest_idx2[1]
port 45 nsew signal input
rlabel metal3 s 0 25304 800 25424 6 dest_idx2[2]
port 46 nsew signal input
rlabel metal3 s 0 25848 800 25968 6 dest_idx2[3]
port 47 nsew signal input
rlabel metal3 s 0 26392 800 26512 6 dest_idx2[4]
port 48 nsew signal input
rlabel metal2 s 115294 127200 115350 128000 6 dest_mask0[0]
port 49 nsew signal input
rlabel metal2 s 116858 127200 116914 128000 6 dest_mask0[1]
port 50 nsew signal input
rlabel metal3 s 419200 23128 420000 23248 6 dest_mask1[0]
port 51 nsew signal input
rlabel metal3 s 419200 23672 420000 23792 6 dest_mask1[1]
port 52 nsew signal input
rlabel metal3 s 0 23128 800 23248 6 dest_mask2[0]
port 53 nsew signal input
rlabel metal3 s 0 23672 800 23792 6 dest_mask2[1]
port 54 nsew signal input
rlabel metal2 s 130934 127200 130990 128000 6 dest_pred0[0]
port 55 nsew signal input
rlabel metal2 s 132498 127200 132554 128000 6 dest_pred0[1]
port 56 nsew signal input
rlabel metal2 s 134062 127200 134118 128000 6 dest_pred0[2]
port 57 nsew signal input
rlabel metal3 s 419200 28568 420000 28688 6 dest_pred1[0]
port 58 nsew signal input
rlabel metal3 s 419200 29112 420000 29232 6 dest_pred1[1]
port 59 nsew signal input
rlabel metal3 s 419200 29656 420000 29776 6 dest_pred1[2]
port 60 nsew signal input
rlabel metal3 s 0 28568 800 28688 6 dest_pred2[0]
port 61 nsew signal input
rlabel metal3 s 0 29112 800 29232 6 dest_pred2[1]
port 62 nsew signal input
rlabel metal3 s 0 29656 800 29776 6 dest_pred2[2]
port 63 nsew signal input
rlabel metal2 s 135626 127200 135682 128000 6 dest_pred_val0
port 64 nsew signal input
rlabel metal3 s 419200 30200 420000 30320 6 dest_pred_val1
port 65 nsew signal input
rlabel metal3 s 0 30200 800 30320 6 dest_pred_val2
port 66 nsew signal input
rlabel metal2 s 65246 127200 65302 128000 6 dest_val0[0]
port 67 nsew signal input
rlabel metal2 s 80886 127200 80942 128000 6 dest_val0[10]
port 68 nsew signal input
rlabel metal2 s 82450 127200 82506 128000 6 dest_val0[11]
port 69 nsew signal input
rlabel metal2 s 84014 127200 84070 128000 6 dest_val0[12]
port 70 nsew signal input
rlabel metal2 s 85578 127200 85634 128000 6 dest_val0[13]
port 71 nsew signal input
rlabel metal2 s 87142 127200 87198 128000 6 dest_val0[14]
port 72 nsew signal input
rlabel metal2 s 88706 127200 88762 128000 6 dest_val0[15]
port 73 nsew signal input
rlabel metal2 s 90270 127200 90326 128000 6 dest_val0[16]
port 74 nsew signal input
rlabel metal2 s 91834 127200 91890 128000 6 dest_val0[17]
port 75 nsew signal input
rlabel metal2 s 93398 127200 93454 128000 6 dest_val0[18]
port 76 nsew signal input
rlabel metal2 s 94962 127200 95018 128000 6 dest_val0[19]
port 77 nsew signal input
rlabel metal2 s 66810 127200 66866 128000 6 dest_val0[1]
port 78 nsew signal input
rlabel metal2 s 96526 127200 96582 128000 6 dest_val0[20]
port 79 nsew signal input
rlabel metal2 s 98090 127200 98146 128000 6 dest_val0[21]
port 80 nsew signal input
rlabel metal2 s 99654 127200 99710 128000 6 dest_val0[22]
port 81 nsew signal input
rlabel metal2 s 101218 127200 101274 128000 6 dest_val0[23]
port 82 nsew signal input
rlabel metal2 s 102782 127200 102838 128000 6 dest_val0[24]
port 83 nsew signal input
rlabel metal2 s 104346 127200 104402 128000 6 dest_val0[25]
port 84 nsew signal input
rlabel metal2 s 105910 127200 105966 128000 6 dest_val0[26]
port 85 nsew signal input
rlabel metal2 s 107474 127200 107530 128000 6 dest_val0[27]
port 86 nsew signal input
rlabel metal2 s 109038 127200 109094 128000 6 dest_val0[28]
port 87 nsew signal input
rlabel metal2 s 110602 127200 110658 128000 6 dest_val0[29]
port 88 nsew signal input
rlabel metal2 s 68374 127200 68430 128000 6 dest_val0[2]
port 89 nsew signal input
rlabel metal2 s 112166 127200 112222 128000 6 dest_val0[30]
port 90 nsew signal input
rlabel metal2 s 113730 127200 113786 128000 6 dest_val0[31]
port 91 nsew signal input
rlabel metal2 s 69938 127200 69994 128000 6 dest_val0[3]
port 92 nsew signal input
rlabel metal2 s 71502 127200 71558 128000 6 dest_val0[4]
port 93 nsew signal input
rlabel metal2 s 73066 127200 73122 128000 6 dest_val0[5]
port 94 nsew signal input
rlabel metal2 s 74630 127200 74686 128000 6 dest_val0[6]
port 95 nsew signal input
rlabel metal2 s 76194 127200 76250 128000 6 dest_val0[7]
port 96 nsew signal input
rlabel metal2 s 77758 127200 77814 128000 6 dest_val0[8]
port 97 nsew signal input
rlabel metal2 s 79322 127200 79378 128000 6 dest_val0[9]
port 98 nsew signal input
rlabel metal3 s 419200 5720 420000 5840 6 dest_val1[0]
port 99 nsew signal input
rlabel metal3 s 419200 11160 420000 11280 6 dest_val1[10]
port 100 nsew signal input
rlabel metal3 s 419200 11704 420000 11824 6 dest_val1[11]
port 101 nsew signal input
rlabel metal3 s 419200 12248 420000 12368 6 dest_val1[12]
port 102 nsew signal input
rlabel metal3 s 419200 12792 420000 12912 6 dest_val1[13]
port 103 nsew signal input
rlabel metal3 s 419200 13336 420000 13456 6 dest_val1[14]
port 104 nsew signal input
rlabel metal3 s 419200 13880 420000 14000 6 dest_val1[15]
port 105 nsew signal input
rlabel metal3 s 419200 14424 420000 14544 6 dest_val1[16]
port 106 nsew signal input
rlabel metal3 s 419200 14968 420000 15088 6 dest_val1[17]
port 107 nsew signal input
rlabel metal3 s 419200 15512 420000 15632 6 dest_val1[18]
port 108 nsew signal input
rlabel metal3 s 419200 16056 420000 16176 6 dest_val1[19]
port 109 nsew signal input
rlabel metal3 s 419200 6264 420000 6384 6 dest_val1[1]
port 110 nsew signal input
rlabel metal3 s 419200 16600 420000 16720 6 dest_val1[20]
port 111 nsew signal input
rlabel metal3 s 419200 17144 420000 17264 6 dest_val1[21]
port 112 nsew signal input
rlabel metal3 s 419200 17688 420000 17808 6 dest_val1[22]
port 113 nsew signal input
rlabel metal3 s 419200 18232 420000 18352 6 dest_val1[23]
port 114 nsew signal input
rlabel metal3 s 419200 18776 420000 18896 6 dest_val1[24]
port 115 nsew signal input
rlabel metal3 s 419200 19320 420000 19440 6 dest_val1[25]
port 116 nsew signal input
rlabel metal3 s 419200 19864 420000 19984 6 dest_val1[26]
port 117 nsew signal input
rlabel metal3 s 419200 20408 420000 20528 6 dest_val1[27]
port 118 nsew signal input
rlabel metal3 s 419200 20952 420000 21072 6 dest_val1[28]
port 119 nsew signal input
rlabel metal3 s 419200 21496 420000 21616 6 dest_val1[29]
port 120 nsew signal input
rlabel metal3 s 419200 6808 420000 6928 6 dest_val1[2]
port 121 nsew signal input
rlabel metal3 s 419200 22040 420000 22160 6 dest_val1[30]
port 122 nsew signal input
rlabel metal3 s 419200 22584 420000 22704 6 dest_val1[31]
port 123 nsew signal input
rlabel metal3 s 419200 7352 420000 7472 6 dest_val1[3]
port 124 nsew signal input
rlabel metal3 s 419200 7896 420000 8016 6 dest_val1[4]
port 125 nsew signal input
rlabel metal3 s 419200 8440 420000 8560 6 dest_val1[5]
port 126 nsew signal input
rlabel metal3 s 419200 8984 420000 9104 6 dest_val1[6]
port 127 nsew signal input
rlabel metal3 s 419200 9528 420000 9648 6 dest_val1[7]
port 128 nsew signal input
rlabel metal3 s 419200 10072 420000 10192 6 dest_val1[8]
port 129 nsew signal input
rlabel metal3 s 419200 10616 420000 10736 6 dest_val1[9]
port 130 nsew signal input
rlabel metal3 s 0 5720 800 5840 6 dest_val2[0]
port 131 nsew signal input
rlabel metal3 s 0 11160 800 11280 6 dest_val2[10]
port 132 nsew signal input
rlabel metal3 s 0 11704 800 11824 6 dest_val2[11]
port 133 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 dest_val2[12]
port 134 nsew signal input
rlabel metal3 s 0 12792 800 12912 6 dest_val2[13]
port 135 nsew signal input
rlabel metal3 s 0 13336 800 13456 6 dest_val2[14]
port 136 nsew signal input
rlabel metal3 s 0 13880 800 14000 6 dest_val2[15]
port 137 nsew signal input
rlabel metal3 s 0 14424 800 14544 6 dest_val2[16]
port 138 nsew signal input
rlabel metal3 s 0 14968 800 15088 6 dest_val2[17]
port 139 nsew signal input
rlabel metal3 s 0 15512 800 15632 6 dest_val2[18]
port 140 nsew signal input
rlabel metal3 s 0 16056 800 16176 6 dest_val2[19]
port 141 nsew signal input
rlabel metal3 s 0 6264 800 6384 6 dest_val2[1]
port 142 nsew signal input
rlabel metal3 s 0 16600 800 16720 6 dest_val2[20]
port 143 nsew signal input
rlabel metal3 s 0 17144 800 17264 6 dest_val2[21]
port 144 nsew signal input
rlabel metal3 s 0 17688 800 17808 6 dest_val2[22]
port 145 nsew signal input
rlabel metal3 s 0 18232 800 18352 6 dest_val2[23]
port 146 nsew signal input
rlabel metal3 s 0 18776 800 18896 6 dest_val2[24]
port 147 nsew signal input
rlabel metal3 s 0 19320 800 19440 6 dest_val2[25]
port 148 nsew signal input
rlabel metal3 s 0 19864 800 19984 6 dest_val2[26]
port 149 nsew signal input
rlabel metal3 s 0 20408 800 20528 6 dest_val2[27]
port 150 nsew signal input
rlabel metal3 s 0 20952 800 21072 6 dest_val2[28]
port 151 nsew signal input
rlabel metal3 s 0 21496 800 21616 6 dest_val2[29]
port 152 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 dest_val2[2]
port 153 nsew signal input
rlabel metal3 s 0 22040 800 22160 6 dest_val2[30]
port 154 nsew signal input
rlabel metal3 s 0 22584 800 22704 6 dest_val2[31]
port 155 nsew signal input
rlabel metal3 s 0 7352 800 7472 6 dest_val2[3]
port 156 nsew signal input
rlabel metal3 s 0 7896 800 8016 6 dest_val2[4]
port 157 nsew signal input
rlabel metal3 s 0 8440 800 8560 6 dest_val2[5]
port 158 nsew signal input
rlabel metal3 s 0 8984 800 9104 6 dest_val2[6]
port 159 nsew signal input
rlabel metal3 s 0 9528 800 9648 6 dest_val2[7]
port 160 nsew signal input
rlabel metal3 s 0 10072 800 10192 6 dest_val2[8]
port 161 nsew signal input
rlabel metal3 s 0 10616 800 10736 6 dest_val2[9]
port 162 nsew signal input
rlabel metal2 s 248234 127200 248290 128000 6 eu0_busy
port 163 nsew signal input
rlabel metal2 s 249798 127200 249854 128000 6 eu0_instruction[0]
port 164 nsew signal output
rlabel metal2 s 265438 127200 265494 128000 6 eu0_instruction[10]
port 165 nsew signal output
rlabel metal2 s 267002 127200 267058 128000 6 eu0_instruction[11]
port 166 nsew signal output
rlabel metal2 s 268566 127200 268622 128000 6 eu0_instruction[12]
port 167 nsew signal output
rlabel metal2 s 270130 127200 270186 128000 6 eu0_instruction[13]
port 168 nsew signal output
rlabel metal2 s 271694 127200 271750 128000 6 eu0_instruction[14]
port 169 nsew signal output
rlabel metal2 s 273258 127200 273314 128000 6 eu0_instruction[15]
port 170 nsew signal output
rlabel metal2 s 274822 127200 274878 128000 6 eu0_instruction[16]
port 171 nsew signal output
rlabel metal2 s 276386 127200 276442 128000 6 eu0_instruction[17]
port 172 nsew signal output
rlabel metal2 s 277950 127200 278006 128000 6 eu0_instruction[18]
port 173 nsew signal output
rlabel metal2 s 279514 127200 279570 128000 6 eu0_instruction[19]
port 174 nsew signal output
rlabel metal2 s 251362 127200 251418 128000 6 eu0_instruction[1]
port 175 nsew signal output
rlabel metal2 s 281078 127200 281134 128000 6 eu0_instruction[20]
port 176 nsew signal output
rlabel metal2 s 282642 127200 282698 128000 6 eu0_instruction[21]
port 177 nsew signal output
rlabel metal2 s 284206 127200 284262 128000 6 eu0_instruction[22]
port 178 nsew signal output
rlabel metal2 s 285770 127200 285826 128000 6 eu0_instruction[23]
port 179 nsew signal output
rlabel metal2 s 287334 127200 287390 128000 6 eu0_instruction[24]
port 180 nsew signal output
rlabel metal2 s 288898 127200 288954 128000 6 eu0_instruction[25]
port 181 nsew signal output
rlabel metal2 s 290462 127200 290518 128000 6 eu0_instruction[26]
port 182 nsew signal output
rlabel metal2 s 292026 127200 292082 128000 6 eu0_instruction[27]
port 183 nsew signal output
rlabel metal2 s 293590 127200 293646 128000 6 eu0_instruction[28]
port 184 nsew signal output
rlabel metal2 s 295154 127200 295210 128000 6 eu0_instruction[29]
port 185 nsew signal output
rlabel metal2 s 252926 127200 252982 128000 6 eu0_instruction[2]
port 186 nsew signal output
rlabel metal2 s 296718 127200 296774 128000 6 eu0_instruction[30]
port 187 nsew signal output
rlabel metal2 s 298282 127200 298338 128000 6 eu0_instruction[31]
port 188 nsew signal output
rlabel metal2 s 299846 127200 299902 128000 6 eu0_instruction[32]
port 189 nsew signal output
rlabel metal2 s 301410 127200 301466 128000 6 eu0_instruction[33]
port 190 nsew signal output
rlabel metal2 s 302974 127200 303030 128000 6 eu0_instruction[34]
port 191 nsew signal output
rlabel metal2 s 304538 127200 304594 128000 6 eu0_instruction[35]
port 192 nsew signal output
rlabel metal2 s 306102 127200 306158 128000 6 eu0_instruction[36]
port 193 nsew signal output
rlabel metal2 s 307666 127200 307722 128000 6 eu0_instruction[37]
port 194 nsew signal output
rlabel metal2 s 309230 127200 309286 128000 6 eu0_instruction[38]
port 195 nsew signal output
rlabel metal2 s 310794 127200 310850 128000 6 eu0_instruction[39]
port 196 nsew signal output
rlabel metal2 s 254490 127200 254546 128000 6 eu0_instruction[3]
port 197 nsew signal output
rlabel metal2 s 312358 127200 312414 128000 6 eu0_instruction[40]
port 198 nsew signal output
rlabel metal2 s 313922 127200 313978 128000 6 eu0_instruction[41]
port 199 nsew signal output
rlabel metal2 s 256054 127200 256110 128000 6 eu0_instruction[4]
port 200 nsew signal output
rlabel metal2 s 257618 127200 257674 128000 6 eu0_instruction[5]
port 201 nsew signal output
rlabel metal2 s 259182 127200 259238 128000 6 eu0_instruction[6]
port 202 nsew signal output
rlabel metal2 s 260746 127200 260802 128000 6 eu0_instruction[7]
port 203 nsew signal output
rlabel metal2 s 262310 127200 262366 128000 6 eu0_instruction[8]
port 204 nsew signal output
rlabel metal2 s 263874 127200 263930 128000 6 eu0_instruction[9]
port 205 nsew signal output
rlabel metal3 s 419200 69368 420000 69488 6 eu1_busy
port 206 nsew signal input
rlabel metal3 s 419200 69912 420000 70032 6 eu1_instruction[0]
port 207 nsew signal output
rlabel metal3 s 419200 75352 420000 75472 6 eu1_instruction[10]
port 208 nsew signal output
rlabel metal3 s 419200 75896 420000 76016 6 eu1_instruction[11]
port 209 nsew signal output
rlabel metal3 s 419200 76440 420000 76560 6 eu1_instruction[12]
port 210 nsew signal output
rlabel metal3 s 419200 76984 420000 77104 6 eu1_instruction[13]
port 211 nsew signal output
rlabel metal3 s 419200 77528 420000 77648 6 eu1_instruction[14]
port 212 nsew signal output
rlabel metal3 s 419200 78072 420000 78192 6 eu1_instruction[15]
port 213 nsew signal output
rlabel metal3 s 419200 78616 420000 78736 6 eu1_instruction[16]
port 214 nsew signal output
rlabel metal3 s 419200 79160 420000 79280 6 eu1_instruction[17]
port 215 nsew signal output
rlabel metal3 s 419200 79704 420000 79824 6 eu1_instruction[18]
port 216 nsew signal output
rlabel metal3 s 419200 80248 420000 80368 6 eu1_instruction[19]
port 217 nsew signal output
rlabel metal3 s 419200 70456 420000 70576 6 eu1_instruction[1]
port 218 nsew signal output
rlabel metal3 s 419200 80792 420000 80912 6 eu1_instruction[20]
port 219 nsew signal output
rlabel metal3 s 419200 81336 420000 81456 6 eu1_instruction[21]
port 220 nsew signal output
rlabel metal3 s 419200 81880 420000 82000 6 eu1_instruction[22]
port 221 nsew signal output
rlabel metal3 s 419200 82424 420000 82544 6 eu1_instruction[23]
port 222 nsew signal output
rlabel metal3 s 419200 82968 420000 83088 6 eu1_instruction[24]
port 223 nsew signal output
rlabel metal3 s 419200 83512 420000 83632 6 eu1_instruction[25]
port 224 nsew signal output
rlabel metal3 s 419200 84056 420000 84176 6 eu1_instruction[26]
port 225 nsew signal output
rlabel metal3 s 419200 84600 420000 84720 6 eu1_instruction[27]
port 226 nsew signal output
rlabel metal3 s 419200 85144 420000 85264 6 eu1_instruction[28]
port 227 nsew signal output
rlabel metal3 s 419200 85688 420000 85808 6 eu1_instruction[29]
port 228 nsew signal output
rlabel metal3 s 419200 71000 420000 71120 6 eu1_instruction[2]
port 229 nsew signal output
rlabel metal3 s 419200 86232 420000 86352 6 eu1_instruction[30]
port 230 nsew signal output
rlabel metal3 s 419200 86776 420000 86896 6 eu1_instruction[31]
port 231 nsew signal output
rlabel metal3 s 419200 87320 420000 87440 6 eu1_instruction[32]
port 232 nsew signal output
rlabel metal3 s 419200 87864 420000 87984 6 eu1_instruction[33]
port 233 nsew signal output
rlabel metal3 s 419200 88408 420000 88528 6 eu1_instruction[34]
port 234 nsew signal output
rlabel metal3 s 419200 88952 420000 89072 6 eu1_instruction[35]
port 235 nsew signal output
rlabel metal3 s 419200 89496 420000 89616 6 eu1_instruction[36]
port 236 nsew signal output
rlabel metal3 s 419200 90040 420000 90160 6 eu1_instruction[37]
port 237 nsew signal output
rlabel metal3 s 419200 90584 420000 90704 6 eu1_instruction[38]
port 238 nsew signal output
rlabel metal3 s 419200 91128 420000 91248 6 eu1_instruction[39]
port 239 nsew signal output
rlabel metal3 s 419200 71544 420000 71664 6 eu1_instruction[3]
port 240 nsew signal output
rlabel metal3 s 419200 91672 420000 91792 6 eu1_instruction[40]
port 241 nsew signal output
rlabel metal3 s 419200 92216 420000 92336 6 eu1_instruction[41]
port 242 nsew signal output
rlabel metal3 s 419200 72088 420000 72208 6 eu1_instruction[4]
port 243 nsew signal output
rlabel metal3 s 419200 72632 420000 72752 6 eu1_instruction[5]
port 244 nsew signal output
rlabel metal3 s 419200 73176 420000 73296 6 eu1_instruction[6]
port 245 nsew signal output
rlabel metal3 s 419200 73720 420000 73840 6 eu1_instruction[7]
port 246 nsew signal output
rlabel metal3 s 419200 74264 420000 74384 6 eu1_instruction[8]
port 247 nsew signal output
rlabel metal3 s 419200 74808 420000 74928 6 eu1_instruction[9]
port 248 nsew signal output
rlabel metal3 s 0 69368 800 69488 6 eu2_busy
port 249 nsew signal input
rlabel metal3 s 0 69912 800 70032 6 eu2_instruction[0]
port 250 nsew signal output
rlabel metal3 s 0 75352 800 75472 6 eu2_instruction[10]
port 251 nsew signal output
rlabel metal3 s 0 75896 800 76016 6 eu2_instruction[11]
port 252 nsew signal output
rlabel metal3 s 0 76440 800 76560 6 eu2_instruction[12]
port 253 nsew signal output
rlabel metal3 s 0 76984 800 77104 6 eu2_instruction[13]
port 254 nsew signal output
rlabel metal3 s 0 77528 800 77648 6 eu2_instruction[14]
port 255 nsew signal output
rlabel metal3 s 0 78072 800 78192 6 eu2_instruction[15]
port 256 nsew signal output
rlabel metal3 s 0 78616 800 78736 6 eu2_instruction[16]
port 257 nsew signal output
rlabel metal3 s 0 79160 800 79280 6 eu2_instruction[17]
port 258 nsew signal output
rlabel metal3 s 0 79704 800 79824 6 eu2_instruction[18]
port 259 nsew signal output
rlabel metal3 s 0 80248 800 80368 6 eu2_instruction[19]
port 260 nsew signal output
rlabel metal3 s 0 70456 800 70576 6 eu2_instruction[1]
port 261 nsew signal output
rlabel metal3 s 0 80792 800 80912 6 eu2_instruction[20]
port 262 nsew signal output
rlabel metal3 s 0 81336 800 81456 6 eu2_instruction[21]
port 263 nsew signal output
rlabel metal3 s 0 81880 800 82000 6 eu2_instruction[22]
port 264 nsew signal output
rlabel metal3 s 0 82424 800 82544 6 eu2_instruction[23]
port 265 nsew signal output
rlabel metal3 s 0 82968 800 83088 6 eu2_instruction[24]
port 266 nsew signal output
rlabel metal3 s 0 83512 800 83632 6 eu2_instruction[25]
port 267 nsew signal output
rlabel metal3 s 0 84056 800 84176 6 eu2_instruction[26]
port 268 nsew signal output
rlabel metal3 s 0 84600 800 84720 6 eu2_instruction[27]
port 269 nsew signal output
rlabel metal3 s 0 85144 800 85264 6 eu2_instruction[28]
port 270 nsew signal output
rlabel metal3 s 0 85688 800 85808 6 eu2_instruction[29]
port 271 nsew signal output
rlabel metal3 s 0 71000 800 71120 6 eu2_instruction[2]
port 272 nsew signal output
rlabel metal3 s 0 86232 800 86352 6 eu2_instruction[30]
port 273 nsew signal output
rlabel metal3 s 0 86776 800 86896 6 eu2_instruction[31]
port 274 nsew signal output
rlabel metal3 s 0 87320 800 87440 6 eu2_instruction[32]
port 275 nsew signal output
rlabel metal3 s 0 87864 800 87984 6 eu2_instruction[33]
port 276 nsew signal output
rlabel metal3 s 0 88408 800 88528 6 eu2_instruction[34]
port 277 nsew signal output
rlabel metal3 s 0 88952 800 89072 6 eu2_instruction[35]
port 278 nsew signal output
rlabel metal3 s 0 89496 800 89616 6 eu2_instruction[36]
port 279 nsew signal output
rlabel metal3 s 0 90040 800 90160 6 eu2_instruction[37]
port 280 nsew signal output
rlabel metal3 s 0 90584 800 90704 6 eu2_instruction[38]
port 281 nsew signal output
rlabel metal3 s 0 91128 800 91248 6 eu2_instruction[39]
port 282 nsew signal output
rlabel metal3 s 0 71544 800 71664 6 eu2_instruction[3]
port 283 nsew signal output
rlabel metal3 s 0 91672 800 91792 6 eu2_instruction[40]
port 284 nsew signal output
rlabel metal3 s 0 92216 800 92336 6 eu2_instruction[41]
port 285 nsew signal output
rlabel metal3 s 0 72088 800 72208 6 eu2_instruction[4]
port 286 nsew signal output
rlabel metal3 s 0 72632 800 72752 6 eu2_instruction[5]
port 287 nsew signal output
rlabel metal3 s 0 73176 800 73296 6 eu2_instruction[6]
port 288 nsew signal output
rlabel metal3 s 0 73720 800 73840 6 eu2_instruction[7]
port 289 nsew signal output
rlabel metal3 s 0 74264 800 74384 6 eu2_instruction[8]
port 290 nsew signal output
rlabel metal3 s 0 74808 800 74928 6 eu2_instruction[9]
port 291 nsew signal output
rlabel metal2 s 5446 0 5502 800 6 io_in[0]
port 292 nsew signal input
rlabel metal2 s 41326 0 41382 800 6 io_in[10]
port 293 nsew signal input
rlabel metal2 s 44914 0 44970 800 6 io_in[11]
port 294 nsew signal input
rlabel metal2 s 48502 0 48558 800 6 io_in[12]
port 295 nsew signal input
rlabel metal2 s 52090 0 52146 800 6 io_in[13]
port 296 nsew signal input
rlabel metal2 s 55678 0 55734 800 6 io_in[14]
port 297 nsew signal input
rlabel metal2 s 59266 0 59322 800 6 io_in[15]
port 298 nsew signal input
rlabel metal2 s 62854 0 62910 800 6 io_in[16]
port 299 nsew signal input
rlabel metal2 s 66442 0 66498 800 6 io_in[17]
port 300 nsew signal input
rlabel metal2 s 70030 0 70086 800 6 io_in[18]
port 301 nsew signal input
rlabel metal2 s 73618 0 73674 800 6 io_in[19]
port 302 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 io_in[1]
port 303 nsew signal input
rlabel metal2 s 77206 0 77262 800 6 io_in[20]
port 304 nsew signal input
rlabel metal2 s 80794 0 80850 800 6 io_in[21]
port 305 nsew signal input
rlabel metal2 s 84382 0 84438 800 6 io_in[22]
port 306 nsew signal input
rlabel metal2 s 87970 0 88026 800 6 io_in[23]
port 307 nsew signal input
rlabel metal2 s 91558 0 91614 800 6 io_in[24]
port 308 nsew signal input
rlabel metal2 s 95146 0 95202 800 6 io_in[25]
port 309 nsew signal input
rlabel metal2 s 98734 0 98790 800 6 io_in[26]
port 310 nsew signal input
rlabel metal2 s 102322 0 102378 800 6 io_in[27]
port 311 nsew signal input
rlabel metal2 s 105910 0 105966 800 6 io_in[28]
port 312 nsew signal input
rlabel metal2 s 109498 0 109554 800 6 io_in[29]
port 313 nsew signal input
rlabel metal2 s 12622 0 12678 800 6 io_in[2]
port 314 nsew signal input
rlabel metal2 s 113086 0 113142 800 6 io_in[30]
port 315 nsew signal input
rlabel metal2 s 116674 0 116730 800 6 io_in[31]
port 316 nsew signal input
rlabel metal2 s 120262 0 120318 800 6 io_in[32]
port 317 nsew signal input
rlabel metal2 s 123850 0 123906 800 6 io_in[33]
port 318 nsew signal input
rlabel metal2 s 127438 0 127494 800 6 io_in[34]
port 319 nsew signal input
rlabel metal2 s 131026 0 131082 800 6 io_in[35]
port 320 nsew signal input
rlabel metal2 s 16210 0 16266 800 6 io_in[3]
port 321 nsew signal input
rlabel metal2 s 19798 0 19854 800 6 io_in[4]
port 322 nsew signal input
rlabel metal2 s 23386 0 23442 800 6 io_in[5]
port 323 nsew signal input
rlabel metal2 s 26974 0 27030 800 6 io_in[6]
port 324 nsew signal input
rlabel metal2 s 30562 0 30618 800 6 io_in[7]
port 325 nsew signal input
rlabel metal2 s 34150 0 34206 800 6 io_in[8]
port 326 nsew signal input
rlabel metal2 s 37738 0 37794 800 6 io_in[9]
port 327 nsew signal input
rlabel metal2 s 134614 0 134670 800 6 io_oeb[0]
port 328 nsew signal output
rlabel metal2 s 170494 0 170550 800 6 io_oeb[10]
port 329 nsew signal output
rlabel metal2 s 174082 0 174138 800 6 io_oeb[11]
port 330 nsew signal output
rlabel metal2 s 177670 0 177726 800 6 io_oeb[12]
port 331 nsew signal output
rlabel metal2 s 181258 0 181314 800 6 io_oeb[13]
port 332 nsew signal output
rlabel metal2 s 184846 0 184902 800 6 io_oeb[14]
port 333 nsew signal output
rlabel metal2 s 188434 0 188490 800 6 io_oeb[15]
port 334 nsew signal output
rlabel metal2 s 192022 0 192078 800 6 io_oeb[16]
port 335 nsew signal output
rlabel metal2 s 195610 0 195666 800 6 io_oeb[17]
port 336 nsew signal output
rlabel metal2 s 199198 0 199254 800 6 io_oeb[18]
port 337 nsew signal output
rlabel metal2 s 202786 0 202842 800 6 io_oeb[19]
port 338 nsew signal output
rlabel metal2 s 138202 0 138258 800 6 io_oeb[1]
port 339 nsew signal output
rlabel metal2 s 206374 0 206430 800 6 io_oeb[20]
port 340 nsew signal output
rlabel metal2 s 209962 0 210018 800 6 io_oeb[21]
port 341 nsew signal output
rlabel metal2 s 213550 0 213606 800 6 io_oeb[22]
port 342 nsew signal output
rlabel metal2 s 217138 0 217194 800 6 io_oeb[23]
port 343 nsew signal output
rlabel metal2 s 220726 0 220782 800 6 io_oeb[24]
port 344 nsew signal output
rlabel metal2 s 224314 0 224370 800 6 io_oeb[25]
port 345 nsew signal output
rlabel metal2 s 227902 0 227958 800 6 io_oeb[26]
port 346 nsew signal output
rlabel metal2 s 231490 0 231546 800 6 io_oeb[27]
port 347 nsew signal output
rlabel metal2 s 235078 0 235134 800 6 io_oeb[28]
port 348 nsew signal output
rlabel metal2 s 238666 0 238722 800 6 io_oeb[29]
port 349 nsew signal output
rlabel metal2 s 141790 0 141846 800 6 io_oeb[2]
port 350 nsew signal output
rlabel metal2 s 242254 0 242310 800 6 io_oeb[30]
port 351 nsew signal output
rlabel metal2 s 245842 0 245898 800 6 io_oeb[31]
port 352 nsew signal output
rlabel metal2 s 249430 0 249486 800 6 io_oeb[32]
port 353 nsew signal output
rlabel metal2 s 253018 0 253074 800 6 io_oeb[33]
port 354 nsew signal output
rlabel metal2 s 256606 0 256662 800 6 io_oeb[34]
port 355 nsew signal output
rlabel metal2 s 260194 0 260250 800 6 io_oeb[35]
port 356 nsew signal output
rlabel metal2 s 145378 0 145434 800 6 io_oeb[3]
port 357 nsew signal output
rlabel metal2 s 148966 0 149022 800 6 io_oeb[4]
port 358 nsew signal output
rlabel metal2 s 152554 0 152610 800 6 io_oeb[5]
port 359 nsew signal output
rlabel metal2 s 156142 0 156198 800 6 io_oeb[6]
port 360 nsew signal output
rlabel metal2 s 159730 0 159786 800 6 io_oeb[7]
port 361 nsew signal output
rlabel metal2 s 163318 0 163374 800 6 io_oeb[8]
port 362 nsew signal output
rlabel metal2 s 166906 0 166962 800 6 io_oeb[9]
port 363 nsew signal output
rlabel metal2 s 263782 0 263838 800 6 io_out[0]
port 364 nsew signal output
rlabel metal2 s 299662 0 299718 800 6 io_out[10]
port 365 nsew signal output
rlabel metal2 s 303250 0 303306 800 6 io_out[11]
port 366 nsew signal output
rlabel metal2 s 306838 0 306894 800 6 io_out[12]
port 367 nsew signal output
rlabel metal2 s 310426 0 310482 800 6 io_out[13]
port 368 nsew signal output
rlabel metal2 s 314014 0 314070 800 6 io_out[14]
port 369 nsew signal output
rlabel metal2 s 317602 0 317658 800 6 io_out[15]
port 370 nsew signal output
rlabel metal2 s 321190 0 321246 800 6 io_out[16]
port 371 nsew signal output
rlabel metal2 s 324778 0 324834 800 6 io_out[17]
port 372 nsew signal output
rlabel metal2 s 328366 0 328422 800 6 io_out[18]
port 373 nsew signal output
rlabel metal2 s 331954 0 332010 800 6 io_out[19]
port 374 nsew signal output
rlabel metal2 s 267370 0 267426 800 6 io_out[1]
port 375 nsew signal output
rlabel metal2 s 335542 0 335598 800 6 io_out[20]
port 376 nsew signal output
rlabel metal2 s 339130 0 339186 800 6 io_out[21]
port 377 nsew signal output
rlabel metal2 s 342718 0 342774 800 6 io_out[22]
port 378 nsew signal output
rlabel metal2 s 346306 0 346362 800 6 io_out[23]
port 379 nsew signal output
rlabel metal2 s 349894 0 349950 800 6 io_out[24]
port 380 nsew signal output
rlabel metal2 s 353482 0 353538 800 6 io_out[25]
port 381 nsew signal output
rlabel metal2 s 357070 0 357126 800 6 io_out[26]
port 382 nsew signal output
rlabel metal2 s 360658 0 360714 800 6 io_out[27]
port 383 nsew signal output
rlabel metal2 s 364246 0 364302 800 6 io_out[28]
port 384 nsew signal output
rlabel metal2 s 367834 0 367890 800 6 io_out[29]
port 385 nsew signal output
rlabel metal2 s 270958 0 271014 800 6 io_out[2]
port 386 nsew signal output
rlabel metal2 s 371422 0 371478 800 6 io_out[30]
port 387 nsew signal output
rlabel metal2 s 375010 0 375066 800 6 io_out[31]
port 388 nsew signal output
rlabel metal2 s 378598 0 378654 800 6 io_out[32]
port 389 nsew signal output
rlabel metal2 s 382186 0 382242 800 6 io_out[33]
port 390 nsew signal output
rlabel metal2 s 385774 0 385830 800 6 io_out[34]
port 391 nsew signal output
rlabel metal2 s 389362 0 389418 800 6 io_out[35]
port 392 nsew signal output
rlabel metal2 s 274546 0 274602 800 6 io_out[3]
port 393 nsew signal output
rlabel metal2 s 278134 0 278190 800 6 io_out[4]
port 394 nsew signal output
rlabel metal2 s 281722 0 281778 800 6 io_out[5]
port 395 nsew signal output
rlabel metal2 s 285310 0 285366 800 6 io_out[6]
port 396 nsew signal output
rlabel metal2 s 288898 0 288954 800 6 io_out[7]
port 397 nsew signal output
rlabel metal2 s 292486 0 292542 800 6 io_out[8]
port 398 nsew signal output
rlabel metal2 s 296074 0 296130 800 6 io_out[9]
port 399 nsew signal output
rlabel metal2 s 187238 127200 187294 128000 6 is_load0
port 400 nsew signal input
rlabel metal3 s 419200 48152 420000 48272 6 is_load1
port 401 nsew signal input
rlabel metal3 s 0 48152 800 48272 6 is_load2
port 402 nsew signal input
rlabel metal2 s 188802 127200 188858 128000 6 is_store0
port 403 nsew signal input
rlabel metal3 s 419200 48696 420000 48816 6 is_store1
port 404 nsew signal input
rlabel metal3 s 0 48696 800 48816 6 is_store2
port 405 nsew signal input
rlabel metal2 s 137190 127200 137246 128000 6 loadstore_address0[0]
port 406 nsew signal input
rlabel metal2 s 152830 127200 152886 128000 6 loadstore_address0[10]
port 407 nsew signal input
rlabel metal2 s 154394 127200 154450 128000 6 loadstore_address0[11]
port 408 nsew signal input
rlabel metal2 s 155958 127200 156014 128000 6 loadstore_address0[12]
port 409 nsew signal input
rlabel metal2 s 157522 127200 157578 128000 6 loadstore_address0[13]
port 410 nsew signal input
rlabel metal2 s 159086 127200 159142 128000 6 loadstore_address0[14]
port 411 nsew signal input
rlabel metal2 s 160650 127200 160706 128000 6 loadstore_address0[15]
port 412 nsew signal input
rlabel metal2 s 162214 127200 162270 128000 6 loadstore_address0[16]
port 413 nsew signal input
rlabel metal2 s 163778 127200 163834 128000 6 loadstore_address0[17]
port 414 nsew signal input
rlabel metal2 s 165342 127200 165398 128000 6 loadstore_address0[18]
port 415 nsew signal input
rlabel metal2 s 166906 127200 166962 128000 6 loadstore_address0[19]
port 416 nsew signal input
rlabel metal2 s 138754 127200 138810 128000 6 loadstore_address0[1]
port 417 nsew signal input
rlabel metal2 s 168470 127200 168526 128000 6 loadstore_address0[20]
port 418 nsew signal input
rlabel metal2 s 170034 127200 170090 128000 6 loadstore_address0[21]
port 419 nsew signal input
rlabel metal2 s 171598 127200 171654 128000 6 loadstore_address0[22]
port 420 nsew signal input
rlabel metal2 s 173162 127200 173218 128000 6 loadstore_address0[23]
port 421 nsew signal input
rlabel metal2 s 174726 127200 174782 128000 6 loadstore_address0[24]
port 422 nsew signal input
rlabel metal2 s 176290 127200 176346 128000 6 loadstore_address0[25]
port 423 nsew signal input
rlabel metal2 s 177854 127200 177910 128000 6 loadstore_address0[26]
port 424 nsew signal input
rlabel metal2 s 179418 127200 179474 128000 6 loadstore_address0[27]
port 425 nsew signal input
rlabel metal2 s 180982 127200 181038 128000 6 loadstore_address0[28]
port 426 nsew signal input
rlabel metal2 s 182546 127200 182602 128000 6 loadstore_address0[29]
port 427 nsew signal input
rlabel metal2 s 140318 127200 140374 128000 6 loadstore_address0[2]
port 428 nsew signal input
rlabel metal2 s 184110 127200 184166 128000 6 loadstore_address0[30]
port 429 nsew signal input
rlabel metal2 s 185674 127200 185730 128000 6 loadstore_address0[31]
port 430 nsew signal input
rlabel metal2 s 141882 127200 141938 128000 6 loadstore_address0[3]
port 431 nsew signal input
rlabel metal2 s 143446 127200 143502 128000 6 loadstore_address0[4]
port 432 nsew signal input
rlabel metal2 s 145010 127200 145066 128000 6 loadstore_address0[5]
port 433 nsew signal input
rlabel metal2 s 146574 127200 146630 128000 6 loadstore_address0[6]
port 434 nsew signal input
rlabel metal2 s 148138 127200 148194 128000 6 loadstore_address0[7]
port 435 nsew signal input
rlabel metal2 s 149702 127200 149758 128000 6 loadstore_address0[8]
port 436 nsew signal input
rlabel metal2 s 151266 127200 151322 128000 6 loadstore_address0[9]
port 437 nsew signal input
rlabel metal3 s 419200 30744 420000 30864 6 loadstore_address1[0]
port 438 nsew signal input
rlabel metal3 s 419200 36184 420000 36304 6 loadstore_address1[10]
port 439 nsew signal input
rlabel metal3 s 419200 36728 420000 36848 6 loadstore_address1[11]
port 440 nsew signal input
rlabel metal3 s 419200 37272 420000 37392 6 loadstore_address1[12]
port 441 nsew signal input
rlabel metal3 s 419200 37816 420000 37936 6 loadstore_address1[13]
port 442 nsew signal input
rlabel metal3 s 419200 38360 420000 38480 6 loadstore_address1[14]
port 443 nsew signal input
rlabel metal3 s 419200 38904 420000 39024 6 loadstore_address1[15]
port 444 nsew signal input
rlabel metal3 s 419200 39448 420000 39568 6 loadstore_address1[16]
port 445 nsew signal input
rlabel metal3 s 419200 39992 420000 40112 6 loadstore_address1[17]
port 446 nsew signal input
rlabel metal3 s 419200 40536 420000 40656 6 loadstore_address1[18]
port 447 nsew signal input
rlabel metal3 s 419200 41080 420000 41200 6 loadstore_address1[19]
port 448 nsew signal input
rlabel metal3 s 419200 31288 420000 31408 6 loadstore_address1[1]
port 449 nsew signal input
rlabel metal3 s 419200 41624 420000 41744 6 loadstore_address1[20]
port 450 nsew signal input
rlabel metal3 s 419200 42168 420000 42288 6 loadstore_address1[21]
port 451 nsew signal input
rlabel metal3 s 419200 42712 420000 42832 6 loadstore_address1[22]
port 452 nsew signal input
rlabel metal3 s 419200 43256 420000 43376 6 loadstore_address1[23]
port 453 nsew signal input
rlabel metal3 s 419200 43800 420000 43920 6 loadstore_address1[24]
port 454 nsew signal input
rlabel metal3 s 419200 44344 420000 44464 6 loadstore_address1[25]
port 455 nsew signal input
rlabel metal3 s 419200 44888 420000 45008 6 loadstore_address1[26]
port 456 nsew signal input
rlabel metal3 s 419200 45432 420000 45552 6 loadstore_address1[27]
port 457 nsew signal input
rlabel metal3 s 419200 45976 420000 46096 6 loadstore_address1[28]
port 458 nsew signal input
rlabel metal3 s 419200 46520 420000 46640 6 loadstore_address1[29]
port 459 nsew signal input
rlabel metal3 s 419200 31832 420000 31952 6 loadstore_address1[2]
port 460 nsew signal input
rlabel metal3 s 419200 47064 420000 47184 6 loadstore_address1[30]
port 461 nsew signal input
rlabel metal3 s 419200 47608 420000 47728 6 loadstore_address1[31]
port 462 nsew signal input
rlabel metal3 s 419200 32376 420000 32496 6 loadstore_address1[3]
port 463 nsew signal input
rlabel metal3 s 419200 32920 420000 33040 6 loadstore_address1[4]
port 464 nsew signal input
rlabel metal3 s 419200 33464 420000 33584 6 loadstore_address1[5]
port 465 nsew signal input
rlabel metal3 s 419200 34008 420000 34128 6 loadstore_address1[6]
port 466 nsew signal input
rlabel metal3 s 419200 34552 420000 34672 6 loadstore_address1[7]
port 467 nsew signal input
rlabel metal3 s 419200 35096 420000 35216 6 loadstore_address1[8]
port 468 nsew signal input
rlabel metal3 s 419200 35640 420000 35760 6 loadstore_address1[9]
port 469 nsew signal input
rlabel metal3 s 0 30744 800 30864 6 loadstore_address2[0]
port 470 nsew signal input
rlabel metal3 s 0 36184 800 36304 6 loadstore_address2[10]
port 471 nsew signal input
rlabel metal3 s 0 36728 800 36848 6 loadstore_address2[11]
port 472 nsew signal input
rlabel metal3 s 0 37272 800 37392 6 loadstore_address2[12]
port 473 nsew signal input
rlabel metal3 s 0 37816 800 37936 6 loadstore_address2[13]
port 474 nsew signal input
rlabel metal3 s 0 38360 800 38480 6 loadstore_address2[14]
port 475 nsew signal input
rlabel metal3 s 0 38904 800 39024 6 loadstore_address2[15]
port 476 nsew signal input
rlabel metal3 s 0 39448 800 39568 6 loadstore_address2[16]
port 477 nsew signal input
rlabel metal3 s 0 39992 800 40112 6 loadstore_address2[17]
port 478 nsew signal input
rlabel metal3 s 0 40536 800 40656 6 loadstore_address2[18]
port 479 nsew signal input
rlabel metal3 s 0 41080 800 41200 6 loadstore_address2[19]
port 480 nsew signal input
rlabel metal3 s 0 31288 800 31408 6 loadstore_address2[1]
port 481 nsew signal input
rlabel metal3 s 0 41624 800 41744 6 loadstore_address2[20]
port 482 nsew signal input
rlabel metal3 s 0 42168 800 42288 6 loadstore_address2[21]
port 483 nsew signal input
rlabel metal3 s 0 42712 800 42832 6 loadstore_address2[22]
port 484 nsew signal input
rlabel metal3 s 0 43256 800 43376 6 loadstore_address2[23]
port 485 nsew signal input
rlabel metal3 s 0 43800 800 43920 6 loadstore_address2[24]
port 486 nsew signal input
rlabel metal3 s 0 44344 800 44464 6 loadstore_address2[25]
port 487 nsew signal input
rlabel metal3 s 0 44888 800 45008 6 loadstore_address2[26]
port 488 nsew signal input
rlabel metal3 s 0 45432 800 45552 6 loadstore_address2[27]
port 489 nsew signal input
rlabel metal3 s 0 45976 800 46096 6 loadstore_address2[28]
port 490 nsew signal input
rlabel metal3 s 0 46520 800 46640 6 loadstore_address2[29]
port 491 nsew signal input
rlabel metal3 s 0 31832 800 31952 6 loadstore_address2[2]
port 492 nsew signal input
rlabel metal3 s 0 47064 800 47184 6 loadstore_address2[30]
port 493 nsew signal input
rlabel metal3 s 0 47608 800 47728 6 loadstore_address2[31]
port 494 nsew signal input
rlabel metal3 s 0 32376 800 32496 6 loadstore_address2[3]
port 495 nsew signal input
rlabel metal3 s 0 32920 800 33040 6 loadstore_address2[4]
port 496 nsew signal input
rlabel metal3 s 0 33464 800 33584 6 loadstore_address2[5]
port 497 nsew signal input
rlabel metal3 s 0 34008 800 34128 6 loadstore_address2[6]
port 498 nsew signal input
rlabel metal3 s 0 34552 800 34672 6 loadstore_address2[7]
port 499 nsew signal input
rlabel metal3 s 0 35096 800 35216 6 loadstore_address2[8]
port 500 nsew signal input
rlabel metal3 s 0 35640 800 35760 6 loadstore_address2[9]
port 501 nsew signal input
rlabel metal2 s 195058 127200 195114 128000 6 loadstore_dest0[0]
port 502 nsew signal input
rlabel metal2 s 196622 127200 196678 128000 6 loadstore_dest0[1]
port 503 nsew signal input
rlabel metal2 s 198186 127200 198242 128000 6 loadstore_dest0[2]
port 504 nsew signal input
rlabel metal2 s 199750 127200 199806 128000 6 loadstore_dest0[3]
port 505 nsew signal input
rlabel metal2 s 201314 127200 201370 128000 6 loadstore_dest0[4]
port 506 nsew signal input
rlabel metal3 s 419200 50872 420000 50992 6 loadstore_dest1[0]
port 507 nsew signal input
rlabel metal3 s 419200 51416 420000 51536 6 loadstore_dest1[1]
port 508 nsew signal input
rlabel metal3 s 419200 51960 420000 52080 6 loadstore_dest1[2]
port 509 nsew signal input
rlabel metal3 s 419200 52504 420000 52624 6 loadstore_dest1[3]
port 510 nsew signal input
rlabel metal3 s 419200 53048 420000 53168 6 loadstore_dest1[4]
port 511 nsew signal input
rlabel metal3 s 0 50872 800 50992 6 loadstore_dest2[0]
port 512 nsew signal input
rlabel metal3 s 0 51416 800 51536 6 loadstore_dest2[1]
port 513 nsew signal input
rlabel metal3 s 0 51960 800 52080 6 loadstore_dest2[2]
port 514 nsew signal input
rlabel metal3 s 0 52504 800 52624 6 loadstore_dest2[3]
port 515 nsew signal input
rlabel metal3 s 0 53048 800 53168 6 loadstore_dest2[4]
port 516 nsew signal input
rlabel metal2 s 191930 127200 191986 128000 6 loadstore_size0[0]
port 517 nsew signal input
rlabel metal2 s 193494 127200 193550 128000 6 loadstore_size0[1]
port 518 nsew signal input
rlabel metal3 s 419200 49784 420000 49904 6 loadstore_size1[0]
port 519 nsew signal input
rlabel metal3 s 419200 50328 420000 50448 6 loadstore_size1[1]
port 520 nsew signal input
rlabel metal3 s 0 49784 800 49904 6 loadstore_size2[0]
port 521 nsew signal input
rlabel metal3 s 0 50328 800 50448 6 loadstore_size2[1]
port 522 nsew signal input
rlabel metal2 s 204442 127200 204498 128000 6 new_PC0[0]
port 523 nsew signal input
rlabel metal2 s 220082 127200 220138 128000 6 new_PC0[10]
port 524 nsew signal input
rlabel metal2 s 221646 127200 221702 128000 6 new_PC0[11]
port 525 nsew signal input
rlabel metal2 s 223210 127200 223266 128000 6 new_PC0[12]
port 526 nsew signal input
rlabel metal2 s 224774 127200 224830 128000 6 new_PC0[13]
port 527 nsew signal input
rlabel metal2 s 226338 127200 226394 128000 6 new_PC0[14]
port 528 nsew signal input
rlabel metal2 s 227902 127200 227958 128000 6 new_PC0[15]
port 529 nsew signal input
rlabel metal2 s 229466 127200 229522 128000 6 new_PC0[16]
port 530 nsew signal input
rlabel metal2 s 231030 127200 231086 128000 6 new_PC0[17]
port 531 nsew signal input
rlabel metal2 s 232594 127200 232650 128000 6 new_PC0[18]
port 532 nsew signal input
rlabel metal2 s 234158 127200 234214 128000 6 new_PC0[19]
port 533 nsew signal input
rlabel metal2 s 206006 127200 206062 128000 6 new_PC0[1]
port 534 nsew signal input
rlabel metal2 s 235722 127200 235778 128000 6 new_PC0[20]
port 535 nsew signal input
rlabel metal2 s 237286 127200 237342 128000 6 new_PC0[21]
port 536 nsew signal input
rlabel metal2 s 238850 127200 238906 128000 6 new_PC0[22]
port 537 nsew signal input
rlabel metal2 s 240414 127200 240470 128000 6 new_PC0[23]
port 538 nsew signal input
rlabel metal2 s 241978 127200 242034 128000 6 new_PC0[24]
port 539 nsew signal input
rlabel metal2 s 243542 127200 243598 128000 6 new_PC0[25]
port 540 nsew signal input
rlabel metal2 s 245106 127200 245162 128000 6 new_PC0[26]
port 541 nsew signal input
rlabel metal2 s 246670 127200 246726 128000 6 new_PC0[27]
port 542 nsew signal input
rlabel metal2 s 207570 127200 207626 128000 6 new_PC0[2]
port 543 nsew signal input
rlabel metal2 s 209134 127200 209190 128000 6 new_PC0[3]
port 544 nsew signal input
rlabel metal2 s 210698 127200 210754 128000 6 new_PC0[4]
port 545 nsew signal input
rlabel metal2 s 212262 127200 212318 128000 6 new_PC0[5]
port 546 nsew signal input
rlabel metal2 s 213826 127200 213882 128000 6 new_PC0[6]
port 547 nsew signal input
rlabel metal2 s 215390 127200 215446 128000 6 new_PC0[7]
port 548 nsew signal input
rlabel metal2 s 216954 127200 217010 128000 6 new_PC0[8]
port 549 nsew signal input
rlabel metal2 s 218518 127200 218574 128000 6 new_PC0[9]
port 550 nsew signal input
rlabel metal3 s 419200 54136 420000 54256 6 new_PC1[0]
port 551 nsew signal input
rlabel metal3 s 419200 59576 420000 59696 6 new_PC1[10]
port 552 nsew signal input
rlabel metal3 s 419200 60120 420000 60240 6 new_PC1[11]
port 553 nsew signal input
rlabel metal3 s 419200 60664 420000 60784 6 new_PC1[12]
port 554 nsew signal input
rlabel metal3 s 419200 61208 420000 61328 6 new_PC1[13]
port 555 nsew signal input
rlabel metal3 s 419200 61752 420000 61872 6 new_PC1[14]
port 556 nsew signal input
rlabel metal3 s 419200 62296 420000 62416 6 new_PC1[15]
port 557 nsew signal input
rlabel metal3 s 419200 62840 420000 62960 6 new_PC1[16]
port 558 nsew signal input
rlabel metal3 s 419200 63384 420000 63504 6 new_PC1[17]
port 559 nsew signal input
rlabel metal3 s 419200 63928 420000 64048 6 new_PC1[18]
port 560 nsew signal input
rlabel metal3 s 419200 64472 420000 64592 6 new_PC1[19]
port 561 nsew signal input
rlabel metal3 s 419200 54680 420000 54800 6 new_PC1[1]
port 562 nsew signal input
rlabel metal3 s 419200 65016 420000 65136 6 new_PC1[20]
port 563 nsew signal input
rlabel metal3 s 419200 65560 420000 65680 6 new_PC1[21]
port 564 nsew signal input
rlabel metal3 s 419200 66104 420000 66224 6 new_PC1[22]
port 565 nsew signal input
rlabel metal3 s 419200 66648 420000 66768 6 new_PC1[23]
port 566 nsew signal input
rlabel metal3 s 419200 67192 420000 67312 6 new_PC1[24]
port 567 nsew signal input
rlabel metal3 s 419200 67736 420000 67856 6 new_PC1[25]
port 568 nsew signal input
rlabel metal3 s 419200 68280 420000 68400 6 new_PC1[26]
port 569 nsew signal input
rlabel metal3 s 419200 68824 420000 68944 6 new_PC1[27]
port 570 nsew signal input
rlabel metal3 s 419200 55224 420000 55344 6 new_PC1[2]
port 571 nsew signal input
rlabel metal3 s 419200 55768 420000 55888 6 new_PC1[3]
port 572 nsew signal input
rlabel metal3 s 419200 56312 420000 56432 6 new_PC1[4]
port 573 nsew signal input
rlabel metal3 s 419200 56856 420000 56976 6 new_PC1[5]
port 574 nsew signal input
rlabel metal3 s 419200 57400 420000 57520 6 new_PC1[6]
port 575 nsew signal input
rlabel metal3 s 419200 57944 420000 58064 6 new_PC1[7]
port 576 nsew signal input
rlabel metal3 s 419200 58488 420000 58608 6 new_PC1[8]
port 577 nsew signal input
rlabel metal3 s 419200 59032 420000 59152 6 new_PC1[9]
port 578 nsew signal input
rlabel metal3 s 0 54136 800 54256 6 new_PC2[0]
port 579 nsew signal input
rlabel metal3 s 0 59576 800 59696 6 new_PC2[10]
port 580 nsew signal input
rlabel metal3 s 0 60120 800 60240 6 new_PC2[11]
port 581 nsew signal input
rlabel metal3 s 0 60664 800 60784 6 new_PC2[12]
port 582 nsew signal input
rlabel metal3 s 0 61208 800 61328 6 new_PC2[13]
port 583 nsew signal input
rlabel metal3 s 0 61752 800 61872 6 new_PC2[14]
port 584 nsew signal input
rlabel metal3 s 0 62296 800 62416 6 new_PC2[15]
port 585 nsew signal input
rlabel metal3 s 0 62840 800 62960 6 new_PC2[16]
port 586 nsew signal input
rlabel metal3 s 0 63384 800 63504 6 new_PC2[17]
port 587 nsew signal input
rlabel metal3 s 0 63928 800 64048 6 new_PC2[18]
port 588 nsew signal input
rlabel metal3 s 0 64472 800 64592 6 new_PC2[19]
port 589 nsew signal input
rlabel metal3 s 0 54680 800 54800 6 new_PC2[1]
port 590 nsew signal input
rlabel metal3 s 0 65016 800 65136 6 new_PC2[20]
port 591 nsew signal input
rlabel metal3 s 0 65560 800 65680 6 new_PC2[21]
port 592 nsew signal input
rlabel metal3 s 0 66104 800 66224 6 new_PC2[22]
port 593 nsew signal input
rlabel metal3 s 0 66648 800 66768 6 new_PC2[23]
port 594 nsew signal input
rlabel metal3 s 0 67192 800 67312 6 new_PC2[24]
port 595 nsew signal input
rlabel metal3 s 0 67736 800 67856 6 new_PC2[25]
port 596 nsew signal input
rlabel metal3 s 0 68280 800 68400 6 new_PC2[26]
port 597 nsew signal input
rlabel metal3 s 0 68824 800 68944 6 new_PC2[27]
port 598 nsew signal input
rlabel metal3 s 0 55224 800 55344 6 new_PC2[2]
port 599 nsew signal input
rlabel metal3 s 0 55768 800 55888 6 new_PC2[3]
port 600 nsew signal input
rlabel metal3 s 0 56312 800 56432 6 new_PC2[4]
port 601 nsew signal input
rlabel metal3 s 0 56856 800 56976 6 new_PC2[5]
port 602 nsew signal input
rlabel metal3 s 0 57400 800 57520 6 new_PC2[6]
port 603 nsew signal input
rlabel metal3 s 0 57944 800 58064 6 new_PC2[7]
port 604 nsew signal input
rlabel metal3 s 0 58488 800 58608 6 new_PC2[8]
port 605 nsew signal input
rlabel metal3 s 0 59032 800 59152 6 new_PC2[9]
port 606 nsew signal input
rlabel metal2 s 126242 127200 126298 128000 6 pred_idx0[0]
port 607 nsew signal input
rlabel metal2 s 127806 127200 127862 128000 6 pred_idx0[1]
port 608 nsew signal input
rlabel metal2 s 129370 127200 129426 128000 6 pred_idx0[2]
port 609 nsew signal input
rlabel metal3 s 419200 26936 420000 27056 6 pred_idx1[0]
port 610 nsew signal input
rlabel metal3 s 419200 27480 420000 27600 6 pred_idx1[1]
port 611 nsew signal input
rlabel metal3 s 419200 28024 420000 28144 6 pred_idx1[2]
port 612 nsew signal input
rlabel metal3 s 0 26936 800 27056 6 pred_idx2[0]
port 613 nsew signal input
rlabel metal3 s 0 27480 800 27600 6 pred_idx2[1]
port 614 nsew signal input
rlabel metal3 s 0 28024 800 28144 6 pred_idx2[2]
port 615 nsew signal input
rlabel metal2 s 415582 127200 415638 128000 6 pred_val0
port 616 nsew signal output
rlabel metal3 s 419200 127576 420000 127696 6 pred_val1
port 617 nsew signal output
rlabel metal3 s 0 127576 800 127696 6 pred_val2
port 618 nsew signal output
rlabel metal2 s 49606 127200 49662 128000 6 reg1_idx0[0]
port 619 nsew signal input
rlabel metal2 s 51170 127200 51226 128000 6 reg1_idx0[1]
port 620 nsew signal input
rlabel metal2 s 52734 127200 52790 128000 6 reg1_idx0[2]
port 621 nsew signal input
rlabel metal2 s 54298 127200 54354 128000 6 reg1_idx0[3]
port 622 nsew signal input
rlabel metal2 s 55862 127200 55918 128000 6 reg1_idx0[4]
port 623 nsew signal input
rlabel metal3 s 419200 280 420000 400 6 reg1_idx1[0]
port 624 nsew signal input
rlabel metal3 s 419200 824 420000 944 6 reg1_idx1[1]
port 625 nsew signal input
rlabel metal3 s 419200 1368 420000 1488 6 reg1_idx1[2]
port 626 nsew signal input
rlabel metal3 s 419200 1912 420000 2032 6 reg1_idx1[3]
port 627 nsew signal input
rlabel metal3 s 419200 2456 420000 2576 6 reg1_idx1[4]
port 628 nsew signal input
rlabel metal3 s 0 280 800 400 6 reg1_idx2[0]
port 629 nsew signal input
rlabel metal3 s 0 824 800 944 6 reg1_idx2[1]
port 630 nsew signal input
rlabel metal3 s 0 1368 800 1488 6 reg1_idx2[2]
port 631 nsew signal input
rlabel metal3 s 0 1912 800 2032 6 reg1_idx2[3]
port 632 nsew signal input
rlabel metal3 s 0 2456 800 2576 6 reg1_idx2[4]
port 633 nsew signal input
rlabel metal2 s 315486 127200 315542 128000 6 reg1_val0[0]
port 634 nsew signal output
rlabel metal2 s 331126 127200 331182 128000 6 reg1_val0[10]
port 635 nsew signal output
rlabel metal2 s 332690 127200 332746 128000 6 reg1_val0[11]
port 636 nsew signal output
rlabel metal2 s 334254 127200 334310 128000 6 reg1_val0[12]
port 637 nsew signal output
rlabel metal2 s 335818 127200 335874 128000 6 reg1_val0[13]
port 638 nsew signal output
rlabel metal2 s 337382 127200 337438 128000 6 reg1_val0[14]
port 639 nsew signal output
rlabel metal2 s 338946 127200 339002 128000 6 reg1_val0[15]
port 640 nsew signal output
rlabel metal2 s 340510 127200 340566 128000 6 reg1_val0[16]
port 641 nsew signal output
rlabel metal2 s 342074 127200 342130 128000 6 reg1_val0[17]
port 642 nsew signal output
rlabel metal2 s 343638 127200 343694 128000 6 reg1_val0[18]
port 643 nsew signal output
rlabel metal2 s 345202 127200 345258 128000 6 reg1_val0[19]
port 644 nsew signal output
rlabel metal2 s 317050 127200 317106 128000 6 reg1_val0[1]
port 645 nsew signal output
rlabel metal2 s 346766 127200 346822 128000 6 reg1_val0[20]
port 646 nsew signal output
rlabel metal2 s 348330 127200 348386 128000 6 reg1_val0[21]
port 647 nsew signal output
rlabel metal2 s 349894 127200 349950 128000 6 reg1_val0[22]
port 648 nsew signal output
rlabel metal2 s 351458 127200 351514 128000 6 reg1_val0[23]
port 649 nsew signal output
rlabel metal2 s 353022 127200 353078 128000 6 reg1_val0[24]
port 650 nsew signal output
rlabel metal2 s 354586 127200 354642 128000 6 reg1_val0[25]
port 651 nsew signal output
rlabel metal2 s 356150 127200 356206 128000 6 reg1_val0[26]
port 652 nsew signal output
rlabel metal2 s 357714 127200 357770 128000 6 reg1_val0[27]
port 653 nsew signal output
rlabel metal2 s 359278 127200 359334 128000 6 reg1_val0[28]
port 654 nsew signal output
rlabel metal2 s 360842 127200 360898 128000 6 reg1_val0[29]
port 655 nsew signal output
rlabel metal2 s 318614 127200 318670 128000 6 reg1_val0[2]
port 656 nsew signal output
rlabel metal2 s 362406 127200 362462 128000 6 reg1_val0[30]
port 657 nsew signal output
rlabel metal2 s 363970 127200 364026 128000 6 reg1_val0[31]
port 658 nsew signal output
rlabel metal2 s 320178 127200 320234 128000 6 reg1_val0[3]
port 659 nsew signal output
rlabel metal2 s 321742 127200 321798 128000 6 reg1_val0[4]
port 660 nsew signal output
rlabel metal2 s 323306 127200 323362 128000 6 reg1_val0[5]
port 661 nsew signal output
rlabel metal2 s 324870 127200 324926 128000 6 reg1_val0[6]
port 662 nsew signal output
rlabel metal2 s 326434 127200 326490 128000 6 reg1_val0[7]
port 663 nsew signal output
rlabel metal2 s 327998 127200 328054 128000 6 reg1_val0[8]
port 664 nsew signal output
rlabel metal2 s 329562 127200 329618 128000 6 reg1_val0[9]
port 665 nsew signal output
rlabel metal3 s 419200 92760 420000 92880 6 reg1_val1[0]
port 666 nsew signal output
rlabel metal3 s 419200 98200 420000 98320 6 reg1_val1[10]
port 667 nsew signal output
rlabel metal3 s 419200 98744 420000 98864 6 reg1_val1[11]
port 668 nsew signal output
rlabel metal3 s 419200 99288 420000 99408 6 reg1_val1[12]
port 669 nsew signal output
rlabel metal3 s 419200 99832 420000 99952 6 reg1_val1[13]
port 670 nsew signal output
rlabel metal3 s 419200 100376 420000 100496 6 reg1_val1[14]
port 671 nsew signal output
rlabel metal3 s 419200 100920 420000 101040 6 reg1_val1[15]
port 672 nsew signal output
rlabel metal3 s 419200 101464 420000 101584 6 reg1_val1[16]
port 673 nsew signal output
rlabel metal3 s 419200 102008 420000 102128 6 reg1_val1[17]
port 674 nsew signal output
rlabel metal3 s 419200 102552 420000 102672 6 reg1_val1[18]
port 675 nsew signal output
rlabel metal3 s 419200 103096 420000 103216 6 reg1_val1[19]
port 676 nsew signal output
rlabel metal3 s 419200 93304 420000 93424 6 reg1_val1[1]
port 677 nsew signal output
rlabel metal3 s 419200 103640 420000 103760 6 reg1_val1[20]
port 678 nsew signal output
rlabel metal3 s 419200 104184 420000 104304 6 reg1_val1[21]
port 679 nsew signal output
rlabel metal3 s 419200 104728 420000 104848 6 reg1_val1[22]
port 680 nsew signal output
rlabel metal3 s 419200 105272 420000 105392 6 reg1_val1[23]
port 681 nsew signal output
rlabel metal3 s 419200 105816 420000 105936 6 reg1_val1[24]
port 682 nsew signal output
rlabel metal3 s 419200 106360 420000 106480 6 reg1_val1[25]
port 683 nsew signal output
rlabel metal3 s 419200 106904 420000 107024 6 reg1_val1[26]
port 684 nsew signal output
rlabel metal3 s 419200 107448 420000 107568 6 reg1_val1[27]
port 685 nsew signal output
rlabel metal3 s 419200 107992 420000 108112 6 reg1_val1[28]
port 686 nsew signal output
rlabel metal3 s 419200 108536 420000 108656 6 reg1_val1[29]
port 687 nsew signal output
rlabel metal3 s 419200 93848 420000 93968 6 reg1_val1[2]
port 688 nsew signal output
rlabel metal3 s 419200 109080 420000 109200 6 reg1_val1[30]
port 689 nsew signal output
rlabel metal3 s 419200 109624 420000 109744 6 reg1_val1[31]
port 690 nsew signal output
rlabel metal3 s 419200 94392 420000 94512 6 reg1_val1[3]
port 691 nsew signal output
rlabel metal3 s 419200 94936 420000 95056 6 reg1_val1[4]
port 692 nsew signal output
rlabel metal3 s 419200 95480 420000 95600 6 reg1_val1[5]
port 693 nsew signal output
rlabel metal3 s 419200 96024 420000 96144 6 reg1_val1[6]
port 694 nsew signal output
rlabel metal3 s 419200 96568 420000 96688 6 reg1_val1[7]
port 695 nsew signal output
rlabel metal3 s 419200 97112 420000 97232 6 reg1_val1[8]
port 696 nsew signal output
rlabel metal3 s 419200 97656 420000 97776 6 reg1_val1[9]
port 697 nsew signal output
rlabel metal3 s 0 92760 800 92880 6 reg1_val2[0]
port 698 nsew signal output
rlabel metal3 s 0 98200 800 98320 6 reg1_val2[10]
port 699 nsew signal output
rlabel metal3 s 0 98744 800 98864 6 reg1_val2[11]
port 700 nsew signal output
rlabel metal3 s 0 99288 800 99408 6 reg1_val2[12]
port 701 nsew signal output
rlabel metal3 s 0 99832 800 99952 6 reg1_val2[13]
port 702 nsew signal output
rlabel metal3 s 0 100376 800 100496 6 reg1_val2[14]
port 703 nsew signal output
rlabel metal3 s 0 100920 800 101040 6 reg1_val2[15]
port 704 nsew signal output
rlabel metal3 s 0 101464 800 101584 6 reg1_val2[16]
port 705 nsew signal output
rlabel metal3 s 0 102008 800 102128 6 reg1_val2[17]
port 706 nsew signal output
rlabel metal3 s 0 102552 800 102672 6 reg1_val2[18]
port 707 nsew signal output
rlabel metal3 s 0 103096 800 103216 6 reg1_val2[19]
port 708 nsew signal output
rlabel metal3 s 0 93304 800 93424 6 reg1_val2[1]
port 709 nsew signal output
rlabel metal3 s 0 103640 800 103760 6 reg1_val2[20]
port 710 nsew signal output
rlabel metal3 s 0 104184 800 104304 6 reg1_val2[21]
port 711 nsew signal output
rlabel metal3 s 0 104728 800 104848 6 reg1_val2[22]
port 712 nsew signal output
rlabel metal3 s 0 105272 800 105392 6 reg1_val2[23]
port 713 nsew signal output
rlabel metal3 s 0 105816 800 105936 6 reg1_val2[24]
port 714 nsew signal output
rlabel metal3 s 0 106360 800 106480 6 reg1_val2[25]
port 715 nsew signal output
rlabel metal3 s 0 106904 800 107024 6 reg1_val2[26]
port 716 nsew signal output
rlabel metal3 s 0 107448 800 107568 6 reg1_val2[27]
port 717 nsew signal output
rlabel metal3 s 0 107992 800 108112 6 reg1_val2[28]
port 718 nsew signal output
rlabel metal3 s 0 108536 800 108656 6 reg1_val2[29]
port 719 nsew signal output
rlabel metal3 s 0 93848 800 93968 6 reg1_val2[2]
port 720 nsew signal output
rlabel metal3 s 0 109080 800 109200 6 reg1_val2[30]
port 721 nsew signal output
rlabel metal3 s 0 109624 800 109744 6 reg1_val2[31]
port 722 nsew signal output
rlabel metal3 s 0 94392 800 94512 6 reg1_val2[3]
port 723 nsew signal output
rlabel metal3 s 0 94936 800 95056 6 reg1_val2[4]
port 724 nsew signal output
rlabel metal3 s 0 95480 800 95600 6 reg1_val2[5]
port 725 nsew signal output
rlabel metal3 s 0 96024 800 96144 6 reg1_val2[6]
port 726 nsew signal output
rlabel metal3 s 0 96568 800 96688 6 reg1_val2[7]
port 727 nsew signal output
rlabel metal3 s 0 97112 800 97232 6 reg1_val2[8]
port 728 nsew signal output
rlabel metal3 s 0 97656 800 97776 6 reg1_val2[9]
port 729 nsew signal output
rlabel metal2 s 57426 127200 57482 128000 6 reg2_idx0[0]
port 730 nsew signal input
rlabel metal2 s 58990 127200 59046 128000 6 reg2_idx0[1]
port 731 nsew signal input
rlabel metal2 s 60554 127200 60610 128000 6 reg2_idx0[2]
port 732 nsew signal input
rlabel metal2 s 62118 127200 62174 128000 6 reg2_idx0[3]
port 733 nsew signal input
rlabel metal2 s 63682 127200 63738 128000 6 reg2_idx0[4]
port 734 nsew signal input
rlabel metal3 s 419200 3000 420000 3120 6 reg2_idx1[0]
port 735 nsew signal input
rlabel metal3 s 419200 3544 420000 3664 6 reg2_idx1[1]
port 736 nsew signal input
rlabel metal3 s 419200 4088 420000 4208 6 reg2_idx1[2]
port 737 nsew signal input
rlabel metal3 s 419200 4632 420000 4752 6 reg2_idx1[3]
port 738 nsew signal input
rlabel metal3 s 419200 5176 420000 5296 6 reg2_idx1[4]
port 739 nsew signal input
rlabel metal3 s 0 3000 800 3120 6 reg2_idx2[0]
port 740 nsew signal input
rlabel metal3 s 0 3544 800 3664 6 reg2_idx2[1]
port 741 nsew signal input
rlabel metal3 s 0 4088 800 4208 6 reg2_idx2[2]
port 742 nsew signal input
rlabel metal3 s 0 4632 800 4752 6 reg2_idx2[3]
port 743 nsew signal input
rlabel metal3 s 0 5176 800 5296 6 reg2_idx2[4]
port 744 nsew signal input
rlabel metal2 s 365534 127200 365590 128000 6 reg2_val0[0]
port 745 nsew signal output
rlabel metal2 s 381174 127200 381230 128000 6 reg2_val0[10]
port 746 nsew signal output
rlabel metal2 s 382738 127200 382794 128000 6 reg2_val0[11]
port 747 nsew signal output
rlabel metal2 s 384302 127200 384358 128000 6 reg2_val0[12]
port 748 nsew signal output
rlabel metal2 s 385866 127200 385922 128000 6 reg2_val0[13]
port 749 nsew signal output
rlabel metal2 s 387430 127200 387486 128000 6 reg2_val0[14]
port 750 nsew signal output
rlabel metal2 s 388994 127200 389050 128000 6 reg2_val0[15]
port 751 nsew signal output
rlabel metal2 s 390558 127200 390614 128000 6 reg2_val0[16]
port 752 nsew signal output
rlabel metal2 s 392122 127200 392178 128000 6 reg2_val0[17]
port 753 nsew signal output
rlabel metal2 s 393686 127200 393742 128000 6 reg2_val0[18]
port 754 nsew signal output
rlabel metal2 s 395250 127200 395306 128000 6 reg2_val0[19]
port 755 nsew signal output
rlabel metal2 s 367098 127200 367154 128000 6 reg2_val0[1]
port 756 nsew signal output
rlabel metal2 s 396814 127200 396870 128000 6 reg2_val0[20]
port 757 nsew signal output
rlabel metal2 s 398378 127200 398434 128000 6 reg2_val0[21]
port 758 nsew signal output
rlabel metal2 s 399942 127200 399998 128000 6 reg2_val0[22]
port 759 nsew signal output
rlabel metal2 s 401506 127200 401562 128000 6 reg2_val0[23]
port 760 nsew signal output
rlabel metal2 s 403070 127200 403126 128000 6 reg2_val0[24]
port 761 nsew signal output
rlabel metal2 s 404634 127200 404690 128000 6 reg2_val0[25]
port 762 nsew signal output
rlabel metal2 s 406198 127200 406254 128000 6 reg2_val0[26]
port 763 nsew signal output
rlabel metal2 s 407762 127200 407818 128000 6 reg2_val0[27]
port 764 nsew signal output
rlabel metal2 s 409326 127200 409382 128000 6 reg2_val0[28]
port 765 nsew signal output
rlabel metal2 s 410890 127200 410946 128000 6 reg2_val0[29]
port 766 nsew signal output
rlabel metal2 s 368662 127200 368718 128000 6 reg2_val0[2]
port 767 nsew signal output
rlabel metal2 s 412454 127200 412510 128000 6 reg2_val0[30]
port 768 nsew signal output
rlabel metal2 s 414018 127200 414074 128000 6 reg2_val0[31]
port 769 nsew signal output
rlabel metal2 s 370226 127200 370282 128000 6 reg2_val0[3]
port 770 nsew signal output
rlabel metal2 s 371790 127200 371846 128000 6 reg2_val0[4]
port 771 nsew signal output
rlabel metal2 s 373354 127200 373410 128000 6 reg2_val0[5]
port 772 nsew signal output
rlabel metal2 s 374918 127200 374974 128000 6 reg2_val0[6]
port 773 nsew signal output
rlabel metal2 s 376482 127200 376538 128000 6 reg2_val0[7]
port 774 nsew signal output
rlabel metal2 s 378046 127200 378102 128000 6 reg2_val0[8]
port 775 nsew signal output
rlabel metal2 s 379610 127200 379666 128000 6 reg2_val0[9]
port 776 nsew signal output
rlabel metal3 s 419200 110168 420000 110288 6 reg2_val1[0]
port 777 nsew signal output
rlabel metal3 s 419200 115608 420000 115728 6 reg2_val1[10]
port 778 nsew signal output
rlabel metal3 s 419200 116152 420000 116272 6 reg2_val1[11]
port 779 nsew signal output
rlabel metal3 s 419200 116696 420000 116816 6 reg2_val1[12]
port 780 nsew signal output
rlabel metal3 s 419200 117240 420000 117360 6 reg2_val1[13]
port 781 nsew signal output
rlabel metal3 s 419200 117784 420000 117904 6 reg2_val1[14]
port 782 nsew signal output
rlabel metal3 s 419200 118328 420000 118448 6 reg2_val1[15]
port 783 nsew signal output
rlabel metal3 s 419200 118872 420000 118992 6 reg2_val1[16]
port 784 nsew signal output
rlabel metal3 s 419200 119416 420000 119536 6 reg2_val1[17]
port 785 nsew signal output
rlabel metal3 s 419200 119960 420000 120080 6 reg2_val1[18]
port 786 nsew signal output
rlabel metal3 s 419200 120504 420000 120624 6 reg2_val1[19]
port 787 nsew signal output
rlabel metal3 s 419200 110712 420000 110832 6 reg2_val1[1]
port 788 nsew signal output
rlabel metal3 s 419200 121048 420000 121168 6 reg2_val1[20]
port 789 nsew signal output
rlabel metal3 s 419200 121592 420000 121712 6 reg2_val1[21]
port 790 nsew signal output
rlabel metal3 s 419200 122136 420000 122256 6 reg2_val1[22]
port 791 nsew signal output
rlabel metal3 s 419200 122680 420000 122800 6 reg2_val1[23]
port 792 nsew signal output
rlabel metal3 s 419200 123224 420000 123344 6 reg2_val1[24]
port 793 nsew signal output
rlabel metal3 s 419200 123768 420000 123888 6 reg2_val1[25]
port 794 nsew signal output
rlabel metal3 s 419200 124312 420000 124432 6 reg2_val1[26]
port 795 nsew signal output
rlabel metal3 s 419200 124856 420000 124976 6 reg2_val1[27]
port 796 nsew signal output
rlabel metal3 s 419200 125400 420000 125520 6 reg2_val1[28]
port 797 nsew signal output
rlabel metal3 s 419200 125944 420000 126064 6 reg2_val1[29]
port 798 nsew signal output
rlabel metal3 s 419200 111256 420000 111376 6 reg2_val1[2]
port 799 nsew signal output
rlabel metal3 s 419200 126488 420000 126608 6 reg2_val1[30]
port 800 nsew signal output
rlabel metal3 s 419200 127032 420000 127152 6 reg2_val1[31]
port 801 nsew signal output
rlabel metal3 s 419200 111800 420000 111920 6 reg2_val1[3]
port 802 nsew signal output
rlabel metal3 s 419200 112344 420000 112464 6 reg2_val1[4]
port 803 nsew signal output
rlabel metal3 s 419200 112888 420000 113008 6 reg2_val1[5]
port 804 nsew signal output
rlabel metal3 s 419200 113432 420000 113552 6 reg2_val1[6]
port 805 nsew signal output
rlabel metal3 s 419200 113976 420000 114096 6 reg2_val1[7]
port 806 nsew signal output
rlabel metal3 s 419200 114520 420000 114640 6 reg2_val1[8]
port 807 nsew signal output
rlabel metal3 s 419200 115064 420000 115184 6 reg2_val1[9]
port 808 nsew signal output
rlabel metal3 s 0 110168 800 110288 6 reg2_val2[0]
port 809 nsew signal output
rlabel metal3 s 0 115608 800 115728 6 reg2_val2[10]
port 810 nsew signal output
rlabel metal3 s 0 116152 800 116272 6 reg2_val2[11]
port 811 nsew signal output
rlabel metal3 s 0 116696 800 116816 6 reg2_val2[12]
port 812 nsew signal output
rlabel metal3 s 0 117240 800 117360 6 reg2_val2[13]
port 813 nsew signal output
rlabel metal3 s 0 117784 800 117904 6 reg2_val2[14]
port 814 nsew signal output
rlabel metal3 s 0 118328 800 118448 6 reg2_val2[15]
port 815 nsew signal output
rlabel metal3 s 0 118872 800 118992 6 reg2_val2[16]
port 816 nsew signal output
rlabel metal3 s 0 119416 800 119536 6 reg2_val2[17]
port 817 nsew signal output
rlabel metal3 s 0 119960 800 120080 6 reg2_val2[18]
port 818 nsew signal output
rlabel metal3 s 0 120504 800 120624 6 reg2_val2[19]
port 819 nsew signal output
rlabel metal3 s 0 110712 800 110832 6 reg2_val2[1]
port 820 nsew signal output
rlabel metal3 s 0 121048 800 121168 6 reg2_val2[20]
port 821 nsew signal output
rlabel metal3 s 0 121592 800 121712 6 reg2_val2[21]
port 822 nsew signal output
rlabel metal3 s 0 122136 800 122256 6 reg2_val2[22]
port 823 nsew signal output
rlabel metal3 s 0 122680 800 122800 6 reg2_val2[23]
port 824 nsew signal output
rlabel metal3 s 0 123224 800 123344 6 reg2_val2[24]
port 825 nsew signal output
rlabel metal3 s 0 123768 800 123888 6 reg2_val2[25]
port 826 nsew signal output
rlabel metal3 s 0 124312 800 124432 6 reg2_val2[26]
port 827 nsew signal output
rlabel metal3 s 0 124856 800 124976 6 reg2_val2[27]
port 828 nsew signal output
rlabel metal3 s 0 125400 800 125520 6 reg2_val2[28]
port 829 nsew signal output
rlabel metal3 s 0 125944 800 126064 6 reg2_val2[29]
port 830 nsew signal output
rlabel metal3 s 0 111256 800 111376 6 reg2_val2[2]
port 831 nsew signal output
rlabel metal3 s 0 126488 800 126608 6 reg2_val2[30]
port 832 nsew signal output
rlabel metal3 s 0 127032 800 127152 6 reg2_val2[31]
port 833 nsew signal output
rlabel metal3 s 0 111800 800 111920 6 reg2_val2[3]
port 834 nsew signal output
rlabel metal3 s 0 112344 800 112464 6 reg2_val2[4]
port 835 nsew signal output
rlabel metal3 s 0 112888 800 113008 6 reg2_val2[5]
port 836 nsew signal output
rlabel metal3 s 0 113432 800 113552 6 reg2_val2[6]
port 837 nsew signal output
rlabel metal3 s 0 113976 800 114096 6 reg2_val2[7]
port 838 nsew signal output
rlabel metal3 s 0 114520 800 114640 6 reg2_val2[8]
port 839 nsew signal output
rlabel metal3 s 0 115064 800 115184 6 reg2_val2[9]
port 840 nsew signal output
rlabel metal2 s 4250 127200 4306 128000 6 rst_eu
port 841 nsew signal output
rlabel metal2 s 396538 0 396594 800 6 rst_n
port 842 nsew signal input
rlabel metal2 s 190366 127200 190422 128000 6 sign_extend0
port 843 nsew signal input
rlabel metal3 s 419200 49240 420000 49360 6 sign_extend1
port 844 nsew signal input
rlabel metal3 s 0 49240 800 49360 6 sign_extend2
port 845 nsew signal input
rlabel metal2 s 202878 127200 202934 128000 6 take_branch0
port 846 nsew signal input
rlabel metal3 s 419200 53592 420000 53712 6 take_branch1
port 847 nsew signal input
rlabel metal3 s 0 53592 800 53712 6 take_branch2
port 848 nsew signal input
rlabel metal4 s 4208 2128 4528 125712 6 vccd1
port 849 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 125712 6 vccd1
port 849 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 125712 6 vccd1
port 849 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 125712 6 vccd1
port 849 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 125712 6 vccd1
port 849 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 125712 6 vccd1
port 849 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 125712 6 vccd1
port 849 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 125712 6 vccd1
port 849 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 125712 6 vccd1
port 849 nsew power bidirectional
rlabel metal4 s 280688 2128 281008 125712 6 vccd1
port 849 nsew power bidirectional
rlabel metal4 s 311408 2128 311728 125712 6 vccd1
port 849 nsew power bidirectional
rlabel metal4 s 342128 2128 342448 125712 6 vccd1
port 849 nsew power bidirectional
rlabel metal4 s 372848 2128 373168 125712 6 vccd1
port 849 nsew power bidirectional
rlabel metal4 s 403568 2128 403888 125712 6 vccd1
port 849 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 125712 6 vssd1
port 850 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 125712 6 vssd1
port 850 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 125712 6 vssd1
port 850 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 125712 6 vssd1
port 850 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 125712 6 vssd1
port 850 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 125712 6 vssd1
port 850 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 125712 6 vssd1
port 850 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 125712 6 vssd1
port 850 nsew ground bidirectional
rlabel metal4 s 265328 2128 265648 125712 6 vssd1
port 850 nsew ground bidirectional
rlabel metal4 s 296048 2128 296368 125712 6 vssd1
port 850 nsew ground bidirectional
rlabel metal4 s 326768 2128 327088 125712 6 vssd1
port 850 nsew ground bidirectional
rlabel metal4 s 357488 2128 357808 125712 6 vssd1
port 850 nsew ground bidirectional
rlabel metal4 s 388208 2128 388528 125712 6 vssd1
port 850 nsew ground bidirectional
rlabel metal2 s 392950 0 393006 800 6 wb_clk_i
port 851 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 420000 128000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 94922248
string GDS_FILE /home/tholin/Desktop/ci2406-rej-pommedeterrible-tholin/openlane/VLIW/runs/24_06_01_14_51/results/signoff/vliw.magic.gds
string GDS_START 1290044
<< end >>

