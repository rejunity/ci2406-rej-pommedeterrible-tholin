* NGSPICE file created from ci2406_z80.ext - technology: sky130B

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_2 abstract view
.subckt sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_4 abstract view
.subckt sky130_fd_sc_hd__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_4 abstract view
.subckt sky130_fd_sc_hd__and2b_4 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_2 abstract view
.subckt sky130_fd_sc_hd__o41ai_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_4 abstract view
.subckt sky130_fd_sc_hd__o2111a_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_4 abstract view
.subckt sky130_fd_sc_hd__a41o_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_4 abstract view
.subckt sky130_fd_sc_hd__o41a_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

.subckt ci2406_z80 custom_settings[0] custom_settings[1] io_in[0] io_in[10] io_in[11]
+ io_in[12] io_in[13] io_in[14] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19]
+ io_in[1] io_in[20] io_in[21] io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[27]
+ io_in[28] io_in[29] io_in[2] io_in[30] io_in[31] io_in[32] io_in[33] io_in[34] io_in[35]
+ io_in[3] io_in[4] io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10]
+ io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18]
+ io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25]
+ io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32]
+ io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[3]
+ io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] rst_n vccd1 vssd1 wb_clk_i
XFILLER_0_94_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3155_ _3193_/B _3379_/B vssd1 vssd1 vccd1 vccd1 _5560_/C sky130_fd_sc_hd__or2_1
XANTENNA__5530__S _5553_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3086_ _6258_/Q _6257_/Q vssd1 vssd1 vccd1 vccd1 _4214_/B sky130_fd_sc_hd__and2_4
XFILLER_0_89_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4640__A1 _6340_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3988_ _6339_/Q _3988_/B vssd1 vssd1 vccd1 vccd1 _3988_/X sky130_fd_sc_hd__or2_1
XFILLER_0_57_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5727_ hold21/X _4243_/B _5727_/S vssd1 vssd1 vccd1 vccd1 hold22/A sky130_fd_sc_hd__mux2_1
XFILLER_0_17_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5658_ _5695_/A1 _3062_/A _5571_/Y _5657_/X vssd1 vssd1 vccd1 vccd1 _5658_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_32_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4609_ _6403_/D _4609_/B vssd1 vssd1 vccd1 vccd1 _4609_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_60_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5589_ _5599_/A _5603_/B _5602_/B _5691_/S vssd1 vssd1 vccd1 vccd1 _5589_/X sky130_fd_sc_hd__and4_2
XFILLER_0_32_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5705__S _6060_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold351 _5977_/X vssd1 vssd1 vccd1 vccd1 _5978_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold340 _6284_/Q vssd1 vssd1 vccd1 vccd1 hold340/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold362 _4293_/X vssd1 vssd1 vccd1 vccd1 _6079_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3733__B _4070_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold384 _5496_/X vssd1 vssd1 vccd1 vccd1 _6328_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold373 _6276_/Q vssd1 vssd1 vccd1 vccd1 hold373/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold395 _6374_/Q vssd1 vssd1 vccd1 vccd1 _5778_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_fanout75_A _3718_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4845__A _6323_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5592__C1 _5673_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3370__A1 _4228_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3643__B _5978_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5647__B1 _5676_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3122__A1 _3254_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4870__B2 _4863_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4960_ _6443_/Q _5056_/A2 _4959_/X vssd1 vssd1 vccd1 vccd1 _4960_/X sky130_fd_sc_hd__a21o_1
XANTENNA__3976__A3 _6339_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3911_ _6216_/Q _3784_/X _3786_/X _6153_/Q vssd1 vssd1 vccd1 vccd1 _3911_/X sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_48_wb_clk_i_A clkbuf_leaf_6_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_4891_ _5849_/S _4890_/X _4883_/X vssd1 vssd1 vccd1 vccd1 _4891_/X sky130_fd_sc_hd__a21o_1
XANTENNA__5586__A _5691_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3842_ _4394_/A _3866_/B vssd1 vssd1 vccd1 vccd1 _3870_/B sky130_fd_sc_hd__or2_1
XFILLER_0_73_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3773_ _5325_/A _3773_/B vssd1 vssd1 vccd1 vccd1 _3773_/X sky130_fd_sc_hd__or2_1
XFILLER_0_42_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5512_ _5512_/A _5512_/B vssd1 vssd1 vccd1 vccd1 _5512_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5443_ _5441_/A _5442_/X _5371_/A vssd1 vssd1 vccd1 vccd1 _5443_/X sky130_fd_sc_hd__o21a_1
XANTENNA__4689__A1 _6032_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5374_ _5368_/Y _5371_/Y _5373_/X _5560_/D vssd1 vssd1 vccd1 vccd1 _5374_/X sky130_fd_sc_hd__a2bb2o_1
XANTENNA__3834__A _3862_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4784__S1 _5358_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4325_ _5053_/S _4324_/X _5727_/S vssd1 vssd1 vccd1 vccd1 _6085_/D sky130_fd_sc_hd__mux2_1
Xfanout138 hold655/X vssd1 vssd1 vccd1 vccd1 _4070_/A sky130_fd_sc_hd__buf_4
Xfanout127 _3611_/A vssd1 vssd1 vccd1 vccd1 _5265_/A sky130_fd_sc_hd__buf_4
Xfanout116 _6427_/Q vssd1 vssd1 vccd1 vccd1 _5553_/S sky130_fd_sc_hd__buf_8
XFILLER_0_10_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout105 _4732_/S vssd1 vssd1 vccd1 vccd1 _6064_/S sky130_fd_sc_hd__clkbuf_8
Xfanout149 _4284_/A vssd1 vssd1 vccd1 vccd1 _4135_/S sky130_fd_sc_hd__buf_2
X_4256_ _3254_/A _3502_/A _4255_/Y _3725_/B vssd1 vssd1 vccd1 vccd1 _4256_/X sky130_fd_sc_hd__a31o_1
X_3207_ _3549_/A _5270_/B _3599_/A _5270_/C vssd1 vssd1 vccd1 vccd1 _5293_/A sky130_fd_sc_hd__a211o_1
X_4187_ _6343_/Q _5328_/C _3747_/B _4186_/Y vssd1 vssd1 vccd1 vccd1 _4187_/X sky130_fd_sc_hd__o211a_1
X_3138_ _3254_/A _3289_/A _3549_/A _3183_/B vssd1 vssd1 vccd1 vccd1 _3379_/B sky130_fd_sc_hd__or4bb_4
XFILLER_0_96_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6063__A0 _4193_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3069_ _5989_/A vssd1 vssd1 vccd1 vccd1 _5069_/A sky130_fd_sc_hd__inv_2
XFILLER_0_92_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5169__A2 _5447_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4604__S _4604_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3447__C _5978_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5435__S _5518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold170 _4336_/X vssd1 vssd1 vccd1 vccd1 _6098_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold192 _3461_/X vssd1 vssd1 vccd1 vccd1 _6206_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold181 _6171_/Q vssd1 vssd1 vccd1 vccd1 hold181/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4301__B1 _5695_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5170__S _5192_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4514__S _4518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3654__A _3654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4540__B1 _5317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5090_ _6301_/Q _5088_/B _6291_/Q _6304_/Q vssd1 vssd1 vccd1 vccd1 _5090_/X sky130_fd_sc_hd__o211a_1
X_4110_ _4394_/A _4110_/B vssd1 vssd1 vccd1 vccd1 _4112_/A sky130_fd_sc_hd__nor2_1
X_4041_ _4042_/A _3746_/X _3985_/A _5211_/C _4040_/A vssd1 vssd1 vccd1 vccd1 _4041_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_75_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6335__RESET_B fanout174/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_4_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_5992_ _6054_/B vssd1 vssd1 vccd1 vccd1 _5992_/Y sky130_fd_sc_hd__inv_2
X_4943_ _6327_/Q _6328_/Q _4943_/C vssd1 vssd1 vccd1 vccd1 _4981_/C sky130_fd_sc_hd__and3_1
XFILLER_0_59_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4874_ _4873_/X _6324_/Q _5825_/S vssd1 vssd1 vccd1 vccd1 _4874_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_6_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3825_ _4111_/A _3826_/B vssd1 vssd1 vccd1 vccd1 _3825_/X sky130_fd_sc_hd__and2_1
XANTENNA_fanout125_A _4214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3756_ _6336_/Q _4188_/C _3746_/X vssd1 vssd1 vccd1 vccd1 _3756_/X sky130_fd_sc_hd__a21o_1
XANTENNA__3564__A _6487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3687_ _6428_/Q _3687_/B vssd1 vssd1 vccd1 vccd1 _3687_/Y sky130_fd_sc_hd__nand2_1
X_5426_ _5426_/A _5426_/B vssd1 vssd1 vccd1 vccd1 _5427_/B sky130_fd_sc_hd__xor2_1
X_5357_ _3359_/B _4758_/C _4323_/B _4322_/Y vssd1 vssd1 vccd1 vccd1 _5357_/Y sky130_fd_sc_hd__o31ai_1
XFILLER_0_10_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5288_ _6256_/Q _3144_/X _3116_/X vssd1 vssd1 vccd1 vccd1 _5288_/Y sky130_fd_sc_hd__o21ai_1
X_4308_ _4309_/A _4313_/D _4313_/B vssd1 vssd1 vccd1 vccd1 _4310_/B sky130_fd_sc_hd__a21oi_1
X_4239_ _3656_/A _4541_/A _3952_/B _5096_/D _4221_/X vssd1 vssd1 vccd1 vccd1 _4239_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_0_97_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4062__A2 _6341_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4334__S _4336_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3474__A _5560_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5078__A1 _4284_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4509__S _4509_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3800__A2 _3779_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3368__B _3369_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3610_ _3645_/B _3606_/Y _4309_/A vssd1 vssd1 vccd1 vccd1 _3610_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_9_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4590_ _6420_/Q _4569_/X _4570_/X _6271_/Q vssd1 vssd1 vccd1 vccd1 _4590_/X sky130_fd_sc_hd__a22o_1
X_3541_ _3541_/A _5354_/B vssd1 vssd1 vccd1 vccd1 _6119_/D sky130_fd_sc_hd__and2_1
XFILLER_0_3_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3384__A _3611_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6260_ _6291_/CLK _6260_/D fanout177/X vssd1 vssd1 vccd1 vccd1 _6260_/Q sky130_fd_sc_hd__dfrtp_1
X_3472_ _3473_/A _3473_/B vssd1 vssd1 vccd1 vccd1 _5739_/A sky130_fd_sc_hd__and2_2
XANTENNA__4739__S1 _5358_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5211_ _5211_/A _5211_/B _5211_/C _5211_/D vssd1 vssd1 vccd1 vccd1 _5212_/C sky130_fd_sc_hd__or4_1
X_6191_ _6407_/CLK hold72/X vssd1 vssd1 vccd1 vccd1 hold71/A sky130_fd_sc_hd__dfxtp_1
X_5142_ _5142_/A _5142_/B vssd1 vssd1 vccd1 vccd1 _5143_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_43_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5073_ hold623/X _5247_/B _4188_/C vssd1 vssd1 vccd1 vccd1 _5241_/S sky130_fd_sc_hd__a21oi_4
X_4024_ _6292_/Q _4066_/B _4073_/C _4023_/Y vssd1 vssd1 vccd1 vccd1 _4025_/B sky130_fd_sc_hd__o22a_1
XFILLER_0_94_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5975_ input7/X hold644/X _5975_/S vssd1 vssd1 vccd1 vccd1 _6423_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_47_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4926_ _6416_/Q _4925_/X _5060_/S vssd1 vssd1 vccd1 vccd1 _4926_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_74_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4857_ _6323_/Q _5852_/S _4856_/X _5557_/S vssd1 vssd1 vccd1 vccd1 _4857_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_74_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3808_ _6134_/Q _3789_/X _3791_/X _6413_/Q vssd1 vssd1 vccd1 vccd1 _3808_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3555__A1 _4224_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4788_ _5058_/S _4788_/B vssd1 vssd1 vccd1 vccd1 _4788_/X sky130_fd_sc_hd__or2_1
XFILLER_0_7_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4201__C1 _5676_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3739_ _6303_/Q _3740_/B vssd1 vssd1 vccd1 vccd1 _3760_/B sky130_fd_sc_hd__and2_1
XFILLER_0_70_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6389_ _6430_/CLK _6389_/D fanout172/X vssd1 vssd1 vccd1 vccd1 _6389_/Q sky130_fd_sc_hd__dfrtp_4
X_5409_ _5450_/A _5408_/B _5408_/C vssd1 vssd1 vccd1 vccd1 _5410_/B sky130_fd_sc_hd__a21o_1
XANTENNA__5713__S _6064_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6257__RESET_B fanout179/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4329__S _4336_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5232__A1 _5242_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4999__S _6315_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5299__A1 _4228_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5578__B _5578_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5760_ _5773_/A _5760_/B vssd1 vssd1 vccd1 vccd1 _5760_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_8_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4711_ hold502/X _4304_/A _4727_/S vssd1 vssd1 vccd1 vccd1 _4711_/X sky130_fd_sc_hd__mux2_1
X_5691_ _4204_/X _5690_/X _5691_/S vssd1 vssd1 vccd1 vccd1 _5691_/X sky130_fd_sc_hd__mux2_1
X_4642_ _5715_/B _4636_/Y _4641_/X hold310/X _4635_/Y vssd1 vssd1 vccd1 vccd1 _4642_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_0_71_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4702__S _4732_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4573_ _5695_/A1 hold429/X _4546_/Y _4572_/X vssd1 vssd1 vccd1 vccd1 _4573_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_4_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3524_ _6118_/Q _5258_/B _5256_/A vssd1 vssd1 vccd1 vccd1 _3524_/X sky130_fd_sc_hd__and3_1
X_6312_ _6401_/CLK _6312_/D fanout179/X vssd1 vssd1 vccd1 vccd1 _6312_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3455_ hold31/X _3449_/X _3464_/A vssd1 vssd1 vccd1 vccd1 hold32/A sky130_fd_sc_hd__a21o_1
X_6243_ _6421_/CLK _6243_/D vssd1 vssd1 vccd1 vccd1 _6243_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_12_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4938__A _5054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3386_ _3386_/A _3386_/B vssd1 vssd1 vccd1 vccd1 _3599_/C sky130_fd_sc_hd__or2_1
X_6174_ _6408_/CLK hold82/X vssd1 vssd1 vccd1 vccd1 hold81/A sky130_fd_sc_hd__dfxtp_1
X_5125_ _5125_/A _5125_/B vssd1 vssd1 vccd1 vccd1 _5128_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_98_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5056_ _6448_/Q _5056_/A2 _5055_/X vssd1 vssd1 vccd1 vccd1 _5056_/X sky130_fd_sc_hd__a21o_1
XANTENNA__4265__A2 _4222_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4673__A _6026_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4007_ _4004_/X _4005_/X _4006_/X _4427_/S vssd1 vssd1 vccd1 vccd1 _4007_/X sky130_fd_sc_hd__a22o_2
XANTENNA__5462__A1 _5715_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_356 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5214__A1 _5560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5958_ _6405_/Q _3639_/C _3627_/Y _3639_/A vssd1 vssd1 vccd1 vccd1 _5958_/X sky130_fd_sc_hd__a22o_1
X_4909_ _6423_/Q _4758_/X _4902_/X _3361_/X _4907_/X vssd1 vssd1 vccd1 vccd1 _4909_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_35_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5889_ _5889_/A _5889_/B vssd1 vssd1 vccd1 vccd1 _5889_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__5708__S _6064_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold669_A _6292_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold41 hold41/A vssd1 vssd1 vccd1 vccd1 hold41/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold30 hold30/A vssd1 vssd1 vccd1 vccd1 hold30/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 hold74/A vssd1 vssd1 vccd1 vccd1 hold74/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold63 hold63/A vssd1 vssd1 vccd1 vccd1 hold63/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 hold52/A vssd1 vssd1 vccd1 vccd1 hold52/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4256__A2 _3502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold96 hold96/A vssd1 vssd1 vccd1 vccd1 hold96/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 hold85/A vssd1 vssd1 vccd1 vccd1 hold85/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_85_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4964__A0 _6418_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3231__A3 _3573_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_14_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6204_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_81_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_5 _4820_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3240_ _4320_/B _3479_/B vssd1 vssd1 vccd1 vccd1 _5292_/B sky130_fd_sc_hd__or2_1
XFILLER_0_67_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3171_ _3525_/A _3220_/A _3379_/B vssd1 vssd1 vccd1 vccd1 _3171_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__3381__B _6389_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5692__A1 _6378_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5444__A1 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6447__SET_B fanout168/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5812_ _5813_/A _5813_/B _5811_/X vssd1 vssd1 vccd1 vccd1 _5821_/B sky130_fd_sc_hd__o21ba_1
XFILLER_0_8_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5743_ _5236_/S _3067_/Y _3580_/A _5735_/X vssd1 vssd1 vccd1 vccd1 _5745_/B sky130_fd_sc_hd__o31a_1
XFILLER_0_84_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4432__S _4437_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5674_ _5674_/A _5674_/B vssd1 vssd1 vccd1 vccd1 _5674_/X sky130_fd_sc_hd__or2_1
X_4625_ input2/X _4631_/B vssd1 vssd1 vccd1 vccd1 _4625_/X sky130_fd_sc_hd__and2_1
XFILLER_0_72_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4556_ _4224_/A _5096_/D _3307_/Y _3572_/A vssd1 vssd1 vccd1 vccd1 _4556_/X sky130_fd_sc_hd__a211o_1
Xhold500 _6247_/Q vssd1 vssd1 vccd1 vccd1 hold500/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold511 _5912_/X vssd1 vssd1 vccd1 vccd1 _6384_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3507_ hold69/X _3507_/B _3507_/C hold37/X vssd1 vssd1 vccd1 vccd1 _3507_/X sky130_fd_sc_hd__or4_1
Xhold544 _6390_/Q vssd1 vssd1 vccd1 vccd1 _3043_/A sky130_fd_sc_hd__buf_1
Xhold533 _4603_/X vssd1 vssd1 vccd1 vccd1 _6248_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold522 _6327_/Q vssd1 vssd1 vccd1 vccd1 hold522/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4668__A _6022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold566 _5945_/X vssd1 vssd1 vccd1 vccd1 hold566/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold588 _6432_/Q vssd1 vssd1 vccd1 vccd1 hold588/X sky130_fd_sc_hd__buf_1
Xhold577 _6332_/Q vssd1 vssd1 vccd1 vccd1 hold577/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold555 _6041_/X vssd1 vssd1 vccd1 vccd1 _6443_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4487_ hold41/X _4399_/X _4491_/S vssd1 vssd1 vccd1 vccd1 hold42/A sky130_fd_sc_hd__mux2_1
X_3438_ hold269/X hold264/X _3438_/S vssd1 vssd1 vccd1 vccd1 _3438_/X sky130_fd_sc_hd__mux2_1
Xhold599 _6294_/Q vssd1 vssd1 vccd1 vccd1 hold599/X sky130_fd_sc_hd__dlygate4sd3_1
X_6226_ _6271_/CLK _6226_/D fanout170/X vssd1 vssd1 vccd1 vccd1 _6226_/Q sky130_fd_sc_hd__dfstp_1
X_3369_ _4679_/C _3369_/B vssd1 vssd1 vccd1 vccd1 _3595_/D sky130_fd_sc_hd__or2_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6157_ _6444_/CLK hold86/X vssd1 vssd1 vccd1 vccd1 hold85/A sky130_fd_sc_hd__dfxtp_1
X_5108_ _4160_/B _4163_/Y _5107_/X vssd1 vssd1 vccd1 vccd1 _5108_/Y sky130_fd_sc_hd__o21ai_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6088_ _6204_/CLK _6088_/D fanout174/X vssd1 vssd1 vccd1 vccd1 _6088_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__5435__A1 _4863_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3446__B1 _5956_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5039_ _6332_/Q _6333_/Q _5039_/C vssd1 vssd1 vccd1 vccd1 _5059_/B sky130_fd_sc_hd__and3_1
XANTENNA__3749__A1 _3952_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4946__A0 _6417_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4342__S _4345_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput42 _6266_/Q vssd1 vssd1 vccd1 vccd1 io_out[27] sky130_fd_sc_hd__buf_12
XANTENNA__3482__A _3482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput31 _6286_/Q vssd1 vssd1 vccd1 vccd1 io_out[17] sky130_fd_sc_hd__buf_12
Xoutput20 _6486_/X vssd1 vssd1 vccd1 vccd1 io_oeb[27] sky130_fd_sc_hd__buf_12
Xoutput53 _6277_/Q vssd1 vssd1 vccd1 vccd1 io_out[8] sky130_fd_sc_hd__buf_12
XFILLER_0_53_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4517__S _4518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_38_wb_clk_i_A clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_85_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4410_ hold5/X _4425_/A2 _4088_/Y _4409_/Y _5597_/B vssd1 vssd1 vccd1 vccd1 _4410_/X
+ sky130_fd_sc_hd__o221a_1
X_5390_ _5388_/X _5389_/X _5560_/D vssd1 vssd1 vccd1 vccd1 _5390_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4341_ hold107/X _4007_/X _4345_/S vssd1 vssd1 vccd1 vccd1 _4341_/X sky130_fd_sc_hd__mux2_1
X_4272_ _3510_/B _3654_/A _5728_/B _4271_/X vssd1 vssd1 vccd1 vccd1 _4273_/D sky130_fd_sc_hd__a31o_1
X_3223_ _3278_/A _3566_/B vssd1 vssd1 vccd1 vccd1 _3431_/A sky130_fd_sc_hd__nor2_1
X_6011_ _3046_/A _6009_/X _6010_/Y hold455/X _5995_/Y vssd1 vssd1 vccd1 vccd1 _6011_/X
+ sky130_fd_sc_hd__o32a_1
XANTENNA__3676__B1 _3566_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3154_ _3683_/C _3206_/B vssd1 vssd1 vccd1 vccd1 _5325_/A sky130_fd_sc_hd__nand2_2
XANTENNA__5417__B2 _5560_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3085_ _3686_/A _3491_/B _3541_/A _5935_/A vssd1 vssd1 vccd1 vccd1 _3359_/B sky130_fd_sc_hd__o31a_2
XANTENNA__4427__S _4427_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3987_ _3748_/Y _4188_/C _3988_/B vssd1 vssd1 vccd1 vccd1 _3987_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_9_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5726_ hold35/X _5725_/Y _5727_/S vssd1 vssd1 vccd1 vccd1 hold36/A sky130_fd_sc_hd__mux2_1
XFILLER_0_45_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5657_ _5657_/A _5657_/B vssd1 vssd1 vccd1 vccd1 _5657_/X sky130_fd_sc_hd__or2_1
X_4608_ _6402_/Q hold316/X _4546_/Y _4607_/X vssd1 vssd1 vccd1 vccd1 _4608_/X sky130_fd_sc_hd__a22o_1
X_5588_ _5603_/A _5610_/A _5603_/D vssd1 vssd1 vccd1 vccd1 _5588_/X sky130_fd_sc_hd__and3_2
XFILLER_0_13_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold352 _5985_/X vssd1 vssd1 vccd1 vccd1 _6428_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4539_ hold468/X _6298_/Q _4539_/S vssd1 vssd1 vccd1 vccd1 _4539_/X sky130_fd_sc_hd__mux2_1
Xhold341 _4954_/X vssd1 vssd1 vccd1 vccd1 _6284_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold330 _6275_/Q vssd1 vssd1 vccd1 vccd1 hold330/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold363 _6285_/Q vssd1 vssd1 vccd1 vccd1 hold363/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold385 _6278_/Q vssd1 vssd1 vccd1 vccd1 hold385/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold374 _4803_/X vssd1 vssd1 vccd1 vccd1 _6276_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold396 _5789_/X vssd1 vssd1 vccd1 vccd1 _6374_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6209_ _6209_/CLK hold74/X vssd1 vssd1 vccd1 vccd1 hold73/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__5656__A1 _6271_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3667__B1 _5096_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5721__S _5723_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4092__B1 _3794_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5592__B1 _3718_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output49_A _3647_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4622__A2 _4615_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3830__B1 _3794_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4890_ _4887_/X _4888_/X _4889_/X _4796_/B _6377_/Q vssd1 vssd1 vccd1 vccd1 _4890_/X
+ sky130_fd_sc_hd__o32a_1
X_3910_ _3724_/A _6036_/A _4391_/A2 vssd1 vssd1 vccd1 vccd1 _3910_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_58_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3841_ _3866_/B vssd1 vssd1 vccd1 vccd1 _3841_/Y sky130_fd_sc_hd__inv_2
X_3772_ _4309_/A _3772_/B vssd1 vssd1 vccd1 vccd1 _3773_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_13_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5511_ _5503_/A _5503_/B _5502_/A vssd1 vssd1 vccd1 vccd1 _5512_/B sky130_fd_sc_hd__a21o_1
XANTENNA__4138__A1 _4255_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4138__B2 _6342_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5442_ _3952_/A _6324_/Q _5442_/S vssd1 vssd1 vccd1 vccd1 _5442_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5335__B1 _5977_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5373_ hold573/X input9/X _5469_/S vssd1 vssd1 vccd1 vccd1 _5373_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4689__A2 _4731_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5107__A _6249_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4324_ _5561_/A _4322_/Y _4323_/X _3363_/A vssd1 vssd1 vccd1 vccd1 _4324_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_10_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout128 _3337_/A vssd1 vssd1 vccd1 vccd1 _3611_/A sky130_fd_sc_hd__buf_4
Xfanout117 hold422/X vssd1 vssd1 vccd1 vccd1 _3473_/A sky130_fd_sc_hd__buf_8
Xfanout106 _5472_/S vssd1 vssd1 vccd1 vccd1 _5727_/S sky130_fd_sc_hd__clkbuf_8
Xfanout139 _6256_/Q vssd1 vssd1 vccd1 vccd1 _3656_/A sky130_fd_sc_hd__clkbuf_8
X_4255_ _4541_/B _4255_/B vssd1 vssd1 vccd1 vccd1 _4255_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__5541__S _5553_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4186_ _6301_/Q _5328_/C vssd1 vssd1 vccd1 vccd1 _4186_/Y sky130_fd_sc_hd__nand2_1
X_3206_ _3206_/A _3206_/B vssd1 vssd1 vccd1 vccd1 _5270_/C sky130_fd_sc_hd__and2_1
X_3137_ _3549_/A _5303_/B _3135_/X vssd1 vssd1 vccd1 vccd1 _3137_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3068_ _6418_/Q vssd1 vssd1 vccd1 vccd1 _5393_/B sky130_fd_sc_hd__inv_2
XFILLER_0_65_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3821__B1 _3781_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3297__A _3573_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5100__B1_N _5193_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5716__S _5723_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5709_ hold19/X _3930_/B _6060_/S vssd1 vssd1 vccd1 vccd1 hold20/A sky130_fd_sc_hd__mux2_1
XANTENNA__5877__A1 _6381_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold171 _6204_/Q vssd1 vssd1 vccd1 vccd1 _3507_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold160 _4490_/X vssd1 vssd1 vccd1 vccd1 _6190_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold182 _4469_/X vssd1 vssd1 vccd1 vccd1 _6171_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold193 _6182_/Q vssd1 vssd1 vccd1 vccd1 hold193/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5629__A1 _6269_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4301__A1 _4305_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4683__A1_N _5740_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5801__A1 _5815_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4698__A1_N _6269_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5801__B2 _5747_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4040_ _4040_/A _5110_/A vssd1 vssd1 vccd1 vccd1 _4046_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_91_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5991_ _5991_/A _5991_/B vssd1 vssd1 vccd1 vccd1 _6054_/B sky130_fd_sc_hd__and2_4
XANTENNA__5597__A _6314_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4705__S _4727_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4942_ _4938_/B _4941_/X _5058_/S vssd1 vssd1 vccd1 vccd1 _4942_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3803__B1 _3794_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6375__RESET_B fanout169/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4873_ _5849_/S _4872_/X _4864_/X vssd1 vssd1 vccd1 vccd1 _4873_/X sky130_fd_sc_hd__a21o_1
XANTENNA__6304__RESET_B fanout180/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3824_ _3824_/A _3824_/B vssd1 vssd1 vccd1 vccd1 _3826_/B sky130_fd_sc_hd__or2_2
X_3755_ _3759_/A _6303_/Q _3755_/C _3938_/A vssd1 vssd1 vccd1 vccd1 _3755_/X sky130_fd_sc_hd__or4_1
XFILLER_0_15_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3582__A2 _5315_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3686_ _3686_/A _6428_/Q _3686_/C vssd1 vssd1 vccd1 vccd1 _3700_/B sky130_fd_sc_hd__and3_2
XANTENNA__4440__S _4446_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5859__A1 _6380_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout118_A _6402_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5425_ _5410_/B _5412_/B _5410_/A vssd1 vssd1 vccd1 vccd1 _5426_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_64_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4531__A1 _6274_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5356_ _5578_/B _3505_/Y _5354_/X _3363_/A vssd1 vssd1 vccd1 vccd1 _5356_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_49_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5287_ _5715_/B hold635/X _5275_/X _5321_/S vssd1 vssd1 vccd1 vccd1 _5287_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3580__A _3580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4307_ _6082_/Q _4307_/B vssd1 vssd1 vccd1 vccd1 _4313_/D sky130_fd_sc_hd__and2_1
X_4238_ _3530_/D _4236_/X _4237_/X vssd1 vssd1 vccd1 vccd1 _4238_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__4295__A0 _6269_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4169_ _5087_/A _5217_/A _6343_/Q _3740_/Y _4168_/X vssd1 vssd1 vccd1 vccd1 _5109_/B
+ sky130_fd_sc_hd__o41a_2
XFILLER_0_77_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4598__A1 _5695_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4598__B2 _4597_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4770__A1 _4637_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3474__B _5975_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5181__S _5447_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5078__A2 _4070_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3490__A _5472_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_39_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6383_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_88_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5210__A _6242_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3540_ _3529_/Y _3536_/X _3538_/X hold359/X vssd1 vssd1 vccd1 vccd1 _3540_/X sky130_fd_sc_hd__a2bb2o_1
XANTENNA__3665__A _5158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3384__B _4734_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5210_ _6242_/Q _5210_/B _5210_/C vssd1 vssd1 vccd1 vccd1 _5219_/D sky130_fd_sc_hd__or3_1
X_3471_ _3471_/A _3471_/B _3471_/C _3471_/D vssd1 vssd1 vccd1 vccd1 _6396_/D sky130_fd_sc_hd__or4_1
XANTENNA__3316__A2 _3309_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6190_ _6408_/CLK _6190_/D vssd1 vssd1 vccd1 vccd1 _6190_/Q sky130_fd_sc_hd__dfxtp_1
X_5141_ _6246_/Q _6247_/Q vssd1 vssd1 vccd1 vccd1 _5142_/B sky130_fd_sc_hd__xor2_1
X_5072_ _6032_/A _5243_/S vssd1 vssd1 vccd1 vccd1 _5072_/Y sky130_fd_sc_hd__nor2_1
X_4023_ _6292_/Q _6295_/Q vssd1 vssd1 vccd1 vccd1 _4023_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4435__S _4437_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5777__B1 _5735_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5974_ input5/X hold643/X _5975_/S vssd1 vssd1 vccd1 vccd1 _6422_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_47_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4925_ _6327_/Q _4943_/C vssd1 vssd1 vccd1 vccd1 _4925_/X sky130_fd_sc_hd__xor2_1
X_4856_ _5773_/A _4855_/X _4844_/X vssd1 vssd1 vccd1 vccd1 _4856_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_7_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3807_ _6190_/Q _3779_/X _3781_/X hold136/X _3806_/X vssd1 vssd1 vccd1 vccd1 _3810_/A
+ sky130_fd_sc_hd__a221o_1
X_4787_ _6372_/Q _6320_/Q _4901_/S vssd1 vssd1 vccd1 vccd1 _4787_/X sky130_fd_sc_hd__mux2_1
X_3738_ _3738_/A _3738_/B vssd1 vssd1 vccd1 vccd1 _3738_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_30_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3669_ _5096_/B _3663_/X _3668_/X vssd1 vssd1 vccd1 vccd1 _3669_/X sky130_fd_sc_hd__o21a_1
X_6388_ _6430_/CLK _6388_/D fanout172/X vssd1 vssd1 vccd1 vccd1 _6388_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__4504__A1 _4392_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5408_ _5450_/A _5408_/B _5408_/C vssd1 vssd1 vccd1 vccd1 _5410_/A sky130_fd_sc_hd__nand3_1
XANTENNA__3712__C1 _3365_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5339_ _5339_/A _5977_/S _5339_/C _5339_/D vssd1 vssd1 vccd1 vccd1 _5339_/X sky130_fd_sc_hd__or4_1
XANTENNA__3514__S _5472_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6009__A1 _5560_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold447_A _6290_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4345__S _4345_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3469__B _5978_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5940__B1 _5935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5299__A2 _3770_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5208__C1 _6304_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6036__A _6036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3234__A1 _3573_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4710_ _6271_/Q _4681_/X _4709_/X _5029_/S vssd1 vssd1 vccd1 vccd1 _4710_/X sky130_fd_sc_hd__a22o_1
X_5690_ _5689_/X _4426_/X _5690_/S vssd1 vssd1 vccd1 vccd1 _5690_/X sky130_fd_sc_hd__mux2_1
X_4641_ _3691_/B _4640_/X _4673_/B vssd1 vssd1 vccd1 vccd1 _4641_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_4_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4572_ _6433_/Q _4567_/Y _4568_/X _6441_/Q _4571_/X vssd1 vssd1 vccd1 vccd1 _4572_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_4_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3523_ _3572_/A _3164_/Y _5584_/A1 vssd1 vssd1 vccd1 vccd1 _3523_/X sky130_fd_sc_hd__o21a_1
X_6311_ _6428_/CLK _6311_/D fanout173/X vssd1 vssd1 vccd1 vccd1 _6311_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3454_ _4558_/A _3581_/A _3457_/C vssd1 vssd1 vccd1 vccd1 _3464_/A sky130_fd_sc_hd__and3_1
X_6242_ _6297_/CLK _6242_/D vssd1 vssd1 vccd1 vccd1 _6242_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__4938__B _4938_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3385_ _4541_/B _5480_/D vssd1 vssd1 vccd1 vccd1 _3385_/Y sky130_fd_sc_hd__nand2_1
X_6173_ _6181_/CLK hold88/X vssd1 vssd1 vccd1 vccd1 hold87/A sky130_fd_sc_hd__dfxtp_1
X_5124_ _5124_/A _5124_/B vssd1 vssd1 vccd1 vccd1 _5125_/B sky130_fd_sc_hd__xnor2_1
X_5055_ _6274_/Q _4758_/X _5054_/B _4757_/Y vssd1 vssd1 vccd1 vccd1 _5055_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_46_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4006_ hold271/X hold107/X hold231/X hold163/X _5676_/C1 _4200_/S vssd1 vssd1 vccd1
+ vccd1 _4006_/X sky130_fd_sc_hd__mux4_2
XFILLER_0_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5462__A2 _6423_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5214__A2 _6297_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5957_ _5715_/B _5956_/Y _3443_/A vssd1 vssd1 vccd1 vccd1 _6402_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_75_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4908_ _6440_/Q _4756_/Y _4757_/Y _4900_/B _4754_/X vssd1 vssd1 vccd1 vccd1 _4908_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_90_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5888_ _5888_/A _5888_/B vssd1 vssd1 vccd1 vccd1 _5892_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_7_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4839_ _4299_/A _4313_/C _5068_/S vssd1 vssd1 vccd1 vccd1 _4839_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3697__D1 _3611_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4567__C _4604_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold31 hold31/A vssd1 vssd1 vccd1 vccd1 hold31/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold20 hold20/A vssd1 vssd1 vccd1 vccd1 hold20/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 hold53/A vssd1 vssd1 vccd1 vccd1 hold53/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 hold64/A vssd1 vssd1 vccd1 vccd1 hold64/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 hold42/A vssd1 vssd1 vccd1 vccd1 hold42/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 hold75/A vssd1 vssd1 vccd1 vccd1 hold75/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold86 hold86/A vssd1 vssd1 vccd1 vccd1 hold86/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 hold97/A vssd1 vssd1 vccd1 vccd1 hold97/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_28_wb_clk_i_A _6404_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4716__A1 _6272_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4716__B2 _5371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_6 _5280_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3170_ _3502_/A _4222_/B _5328_/B _3600_/B vssd1 vssd1 vccd1 vccd1 _3170_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_83_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5589__B _5603_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xci2406_z80_210 vssd1 vssd1 vccd1 vccd1 io_oeb[4] ci2406_z80_210/LO sky130_fd_sc_hd__conb_1
XFILLER_0_16_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5811_ _5821_/A _5811_/B vssd1 vssd1 vccd1 vccd1 _5811_/X sky130_fd_sc_hd__or2_1
XFILLER_0_29_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4713__S _4731_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5742_ _5742_/A vssd1 vssd1 vccd1 vccd1 _5742_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_84_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5673_ _6134_/Q _6313_/Q _4384_/S _6213_/Q _5673_/C1 vssd1 vssd1 vccd1 vccd1 _5674_/B
+ sky130_fd_sc_hd__o221a_1
X_4624_ _3525_/A _4615_/X _4617_/Y _4623_/X vssd1 vssd1 vccd1 vccd1 _6254_/D sky130_fd_sc_hd__o22a_1
XFILLER_0_13_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4555_ _4217_/X _4548_/X _4553_/X _4554_/X vssd1 vssd1 vccd1 vccd1 _4555_/X sky130_fd_sc_hd__o31a_1
Xhold501 _4598_/X vssd1 vssd1 vccd1 vccd1 _6247_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout100_A _4639_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold545 _5947_/X vssd1 vssd1 vccd1 vccd1 hold545/X sky130_fd_sc_hd__dlygate4sd3_1
X_3506_ _3486_/B _3505_/Y _5354_/B _3491_/B vssd1 vssd1 vccd1 vccd1 _6117_/D sky130_fd_sc_hd__a2bb2o_1
Xhold512 _6331_/Q vssd1 vssd1 vccd1 vccd1 _5526_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold534 _6365_/Q vssd1 vssd1 vccd1 vccd1 hold534/X sky130_fd_sc_hd__buf_1
Xhold523 _5487_/X vssd1 vssd1 vccd1 vccd1 _6327_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold556 _6394_/Q vssd1 vssd1 vccd1 vccd1 _5728_/A sky130_fd_sc_hd__buf_1
XANTENNA__3572__B _3770_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold567 _5946_/X vssd1 vssd1 vccd1 vccd1 _6390_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4486_ hold39/X _4392_/X _4491_/S vssd1 vssd1 vccd1 vccd1 hold40/A sky130_fd_sc_hd__mux2_1
Xhold578 _5540_/X vssd1 vssd1 vccd1 vccd1 _6332_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold589 _3641_/X vssd1 vssd1 vccd1 vccd1 _6432_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3437_ hold306/X _3435_/Y _3436_/X vssd1 vssd1 vccd1 vccd1 _3437_/X sky130_fd_sc_hd__a21o_1
X_6225_ _6271_/CLK _6225_/D fanout170/X vssd1 vssd1 vccd1 vccd1 _6225_/Q sky130_fd_sc_hd__dfstp_1
X_3368_ _4679_/C _3369_/B vssd1 vssd1 vccd1 vccd1 _3511_/A sky130_fd_sc_hd__nor2_2
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6156_ _6331_/CLK _6156_/D vssd1 vssd1 vccd1 vccd1 _6156_/Q sky130_fd_sc_hd__dfxtp_1
X_5107_ _6249_/Q _5107_/B _4160_/B vssd1 vssd1 vccd1 vccd1 _5107_/X sky130_fd_sc_hd__or3b_1
XANTENNA__4684__A _5226_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6087_ _6204_/CLK _6087_/D fanout174/X vssd1 vssd1 vccd1 vccd1 _6087_/Q sky130_fd_sc_hd__dfrtp_1
X_3299_ _5325_/A _5256_/A _3299_/C vssd1 vssd1 vccd1 vccd1 _3299_/X sky130_fd_sc_hd__and3_1
XANTENNA__4643__A0 _6243_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3446__A1 _5560_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5038_ _6057_/C _5037_/X _5058_/S vssd1 vssd1 vccd1 vccd1 _5038_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_79_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3997__A2 _3784_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5719__S _5723_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3382__B1 _4541_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput43 _6260_/Q vssd1 vssd1 vccd1 vccd1 io_out[28] sky130_fd_sc_hd__buf_12
XANTENNA__3482__B _5560_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput32 _6287_/Q vssd1 vssd1 vccd1 vccd1 io_out[18] sky130_fd_sc_hd__buf_12
Xoutput21 _6487_/X vssd1 vssd1 vccd1 vccd1 io_oeb[28] sky130_fd_sc_hd__buf_12
XANTENNA__5659__C1 _5675_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput54 _6275_/Q vssd1 vssd1 vccd1 vccd1 io_out[9] sky130_fd_sc_hd__buf_12
XANTENNA__4594__A _4594_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5362__B2 _4214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3912__A2 _3779_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4340_ hold63/X _3965_/X _4345_/S vssd1 vssd1 vccd1 vccd1 hold64/A sky130_fd_sc_hd__mux2_1
X_4271_ _3656_/A _5323_/C _4269_/X _5563_/C _4216_/A vssd1 vssd1 vccd1 vccd1 _4271_/X
+ sky130_fd_sc_hd__a311o_1
X_3222_ _3254_/A _3566_/A _3566_/B vssd1 vssd1 vccd1 vccd1 _5158_/A sky130_fd_sc_hd__or3_4
XANTENNA__6329__RESET_B fanout168/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6010_ _6044_/A _6026_/B vssd1 vssd1 vccd1 vccd1 _6010_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__3676__A1 _3254_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3153_ _3683_/C _3206_/B vssd1 vssd1 vccd1 vccd1 _3661_/A sky130_fd_sc_hd__and2_2
XANTENNA__4708__S _5447_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4443__S _4446_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout148_A _4284_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3986_ _5209_/A _5123_/B _5216_/D _3761_/A vssd1 vssd1 vccd1 vccd1 _3986_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_76_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4928__A1 _6379_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5725_ _5725_/A _5725_/B vssd1 vssd1 vccd1 vccd1 _5725_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_94_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5656_ _6271_/Q _5589_/X _5610_/X hold399/X _5655_/X vssd1 vssd1 vccd1 vccd1 _5657_/B
+ sky130_fd_sc_hd__a221o_1
X_4607_ _4564_/A _4604_/X _4606_/X vssd1 vssd1 vccd1 vccd1 _4607_/X sky130_fd_sc_hd__a21o_1
XANTENNA__4679__A _4679_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5587_ _5599_/A _5610_/A _5691_/S vssd1 vssd1 vccd1 vccd1 _5587_/X sky130_fd_sc_hd__and3_2
XFILLER_0_13_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold320 _4859_/X vssd1 vssd1 vccd1 vccd1 _6279_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4538_ hold459/X _6297_/Q _4539_/S vssd1 vssd1 vccd1 vccd1 _4538_/X sky130_fd_sc_hd__mux2_1
Xhold353 _6345_/Q vssd1 vssd1 vccd1 vccd1 _3080_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold331 _4782_/X vssd1 vssd1 vccd1 vccd1 _6275_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold342 _6352_/Q vssd1 vssd1 vccd1 vccd1 _3078_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold375 _6337_/Q vssd1 vssd1 vccd1 vccd1 _3907_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold364 _4972_/X vssd1 vssd1 vccd1 vccd1 _6285_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold386 _4840_/X vssd1 vssd1 vccd1 vccd1 _6278_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4469_ _4399_/X hold181/X _4473_/S vssd1 vssd1 vccd1 vccd1 _4469_/X sky130_fd_sc_hd__mux2_1
X_6208_ _6344_/CLK hold58/X vssd1 vssd1 vccd1 vccd1 hold57/A sky130_fd_sc_hd__dfxtp_1
Xhold397 _6360_/Q vssd1 vssd1 vccd1 vccd1 hold397/X sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6139_ _6218_/CLK _6139_/D vssd1 vssd1 vccd1 vccd1 _6139_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5449__S _5553_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4353__S _4360_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4552__C1 _4222_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5647__A2 _4198_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3840_ _3863_/A _3839_/X _3836_/Y _3834_/Y vssd1 vssd1 vccd1 vccd1 _3866_/B sky130_fd_sc_hd__o2bb2a_2
XANTENNA__6044__A _6044_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5583__A1 _5096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3771_ _3772_/B vssd1 vssd1 vccd1 vccd1 _3771_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_6_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4386__A2 _4382_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5510_ _5554_/A _5510_/B vssd1 vssd1 vccd1 vccd1 _5512_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_89_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5441_ _5441_/A _5441_/B vssd1 vssd1 vccd1 vccd1 _5441_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__5335__A1 _5725_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5372_ _5739_/A _5372_/B _5372_/C vssd1 vssd1 vccd1 vccd1 _5469_/S sky130_fd_sc_hd__and3_4
XFILLER_0_10_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4323_ _4323_/A _4323_/B vssd1 vssd1 vccd1 vccd1 _4323_/X sky130_fd_sc_hd__or2_1
XFILLER_0_10_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout129 _3337_/A vssd1 vssd1 vccd1 vccd1 _5578_/A sky130_fd_sc_hd__clkbuf_8
Xfanout107 _4732_/S vssd1 vssd1 vccd1 vccd1 _5472_/S sky130_fd_sc_hd__buf_4
XFILLER_0_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout118 _6402_/Q vssd1 vssd1 vccd1 vccd1 _3046_/A sky130_fd_sc_hd__clkbuf_8
X_4254_ _3152_/A _5315_/A _4273_/A _4252_/X _5563_/B vssd1 vssd1 vccd1 vccd1 _4254_/X
+ sky130_fd_sc_hd__a2111o_1
XANTENNA__3850__B _3850_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4185_ _5217_/A _4081_/S _4184_/X _3323_/X vssd1 vssd1 vccd1 vccd1 _5212_/B sky130_fd_sc_hd__a211o_1
X_3205_ _3290_/B _4679_/D vssd1 vssd1 vccd1 vccd1 _4747_/C sky130_fd_sc_hd__or2_1
X_3136_ _3254_/A _3136_/B _3293_/B vssd1 vssd1 vccd1 vccd1 _5303_/B sky130_fd_sc_hd__or3_4
X_3067_ _6416_/Q vssd1 vssd1 vccd1 vccd1 _3067_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_89_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3969_ _5088_/B _3969_/B vssd1 vssd1 vccd1 vccd1 _3969_/X sky130_fd_sc_hd__or2_1
X_5708_ hold13/X _3916_/Y _6064_/S vssd1 vssd1 vccd1 vccd1 hold14/A sky130_fd_sc_hd__mux2_1
XANTENNA__4901__S _4901_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5639_ _5638_/X _5635_/X _4006_/X _4398_/X _5691_/S _5690_/S vssd1 vssd1 vccd1 vccd1
+ _5639_/X sky130_fd_sc_hd__mux4_2
Xhold150 _4455_/X vssd1 vssd1 vccd1 vccd1 _6159_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold161 _6210_/Q vssd1 vssd1 vccd1 vccd1 hold161/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 _3456_/X vssd1 vssd1 vccd1 vccd1 _6204_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold183 _6154_/Q vssd1 vssd1 vccd1 vccd1 hold183/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold194 _4481_/X vssd1 vssd1 vccd1 vccd1 _6182_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout80_A _4319_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3101__A_N _3183_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold644_A _6423_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3488__A _4541_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5565__A1 _3656_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5565__B2 _5578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3576__B1 _5313_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4811__S _5058_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5990_ _3611_/A _6428_/Q _5739_/A vssd1 vssd1 vccd1 vccd1 _5991_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_91_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3264__C1 _3632_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4941_ _6380_/Q _6328_/Q _6315_/Q vssd1 vssd1 vccd1 vccd1 _4941_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5597__B _5597_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3398__A _5258_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4872_ _4867_/X _4870_/X _4871_/X _4796_/B _6376_/Q vssd1 vssd1 vccd1 vccd1 _4872_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_0_86_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3823_ _6180_/Q _3715_/X _3794_/X _6211_/Q _3822_/X vssd1 vssd1 vccd1 vccd1 _3824_/B
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5556__B2 _5441_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3754_ _6303_/Q _6301_/Q _5087_/A _6304_/Q vssd1 vssd1 vccd1 vccd1 _4188_/C sky130_fd_sc_hd__and4b_4
XFILLER_0_61_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_9_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6428_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__4721__S _4727_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3685_ _5518_/S _3687_/B vssd1 vssd1 vccd1 vccd1 _4197_/B sky130_fd_sc_hd__nand2_8
XFILLER_0_30_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5424_ _5422_/X _5424_/B vssd1 vssd1 vccd1 vccd1 _5426_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_100_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5355_ _3656_/A _3505_/Y _5354_/X _3363_/B vssd1 vssd1 vccd1 vccd1 _5355_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_57_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5286_ _5715_/B _5746_/A vssd1 vssd1 vccd1 vccd1 _5321_/S sky130_fd_sc_hd__nor2_2
X_4306_ _4304_/A _4301_/X _4305_/X _6064_/S vssd1 vssd1 vccd1 vccd1 _4306_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4819__B1 _5728_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4237_ _3289_/A _6118_/Q _5584_/A1 vssd1 vssd1 vccd1 vccd1 _4237_/X sky130_fd_sc_hd__a21o_1
X_4168_ _3740_/Y _4162_/X _4163_/Y _4167_/X vssd1 vssd1 vccd1 vccd1 _4168_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_97_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6066__3 _6270_/CLK vssd1 vssd1 vccd1 vccd1 _6124_/CLK sky130_fd_sc_hd__inv_2
X_3119_ _4679_/A _3220_/A vssd1 vssd1 vccd1 vccd1 _4522_/D sky130_fd_sc_hd__or2_2
X_4099_ _3724_/A _5253_/B _4088_/Y vssd1 vssd1 vccd1 vccd1 _4099_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_77_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5547__B2 _5377_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3490__B _4287_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5235__A0 _6298_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3470_ hold69/X hold47/X _3507_/C hold33/X _3449_/X vssd1 vssd1 vccd1 vccd1 _3471_/D
+ sky130_fd_sc_hd__o41a_1
XFILLER_0_10_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5140_ _5140_/A _5140_/B vssd1 vssd1 vccd1 vccd1 _5143_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__4286__C_N _4727_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5071_ _5243_/S vssd1 vssd1 vccd1 vccd1 _5098_/A sky130_fd_sc_hd__inv_2
XFILLER_0_19_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4022_ _4022_/A _4022_/B vssd1 vssd1 vccd1 vccd1 _4022_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5973_ input4/X hold642/X _5975_/S vssd1 vssd1 vccd1 vccd1 _6421_/D sky130_fd_sc_hd__mux2_1
XANTENNA__5777__A1 _5236_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4924_ _4920_/B _4923_/X _5058_/S vssd1 vssd1 vccd1 vccd1 _4924_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_59_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4855_ _6323_/Q _5928_/A2 _5850_/B1 _4854_/X vssd1 vssd1 vccd1 vccd1 _4855_/X sky130_fd_sc_hd__a22o_1
XANTENNA_fanout130_A _4309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4786_ _4785_/X _4784_/X _5053_/S vssd1 vssd1 vccd1 vccd1 _4788_/B sky130_fd_sc_hd__mux2_2
XANTENNA__4451__S _4455_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3806_ hold89/A _3784_/X _3786_/X hold81/A vssd1 vssd1 vccd1 vccd1 _3806_/X sky130_fd_sc_hd__a22o_1
X_3737_ _3738_/A _3738_/B vssd1 vssd1 vccd1 vccd1 _3737_/X sky130_fd_sc_hd__or2_1
XFILLER_0_7_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3668_ _3668_/A _4220_/B _3668_/C vssd1 vssd1 vccd1 vccd1 _3668_/X sky130_fd_sc_hd__or3_2
XFILLER_0_15_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3599_ _3599_/A _3657_/A _3599_/C vssd1 vssd1 vccd1 vccd1 _5272_/B sky130_fd_sc_hd__or3_1
X_6387_ _6430_/CLK _6387_/D fanout172/X vssd1 vssd1 vccd1 vccd1 _6387_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_0_11_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5407_ _6436_/Q _4830_/B _5553_/S vssd1 vssd1 vccd1 vccd1 _5408_/C sky130_fd_sc_hd__mux2_1
XFILLER_0_100_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5338_ _5988_/B _5337_/Y _5727_/S vssd1 vssd1 vccd1 vccd1 _5338_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_100_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5269_ _5322_/A _5715_/C _4734_/C _3511_/A vssd1 vssd1 vccd1 vccd1 _5273_/B sky130_fd_sc_hd__a211o_1
XFILLER_0_76_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_18_wb_clk_i_A _6404_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6016__A2_N _6054_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6266__RESET_B fanout177/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5192__S _5192_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4259__A1 _3594_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6036__B _6063_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3234__A2 _4228_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4640_ _4638_/X _6340_/Q _4675_/S vssd1 vssd1 vccd1 vccd1 _4640_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6052__A _6052_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6310_ _6433_/CLK _6310_/D fanout173/X vssd1 vssd1 vccd1 vccd1 _6310_/Q sky130_fd_sc_hd__dfrtp_1
X_4571_ _6416_/Q _4569_/X _4570_/X _6267_/Q _4566_/Y vssd1 vssd1 vccd1 vccd1 _4571_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_24_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3522_ _5293_/A _3515_/X _3521_/X _3530_/D vssd1 vssd1 vccd1 vccd1 _3522_/X sky130_fd_sc_hd__o31a_1
XFILLER_0_4_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3453_ _3466_/B _3453_/B vssd1 vssd1 vccd1 vccd1 _3457_/C sky130_fd_sc_hd__and2b_1
XFILLER_0_12_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6241_ _6290_/CLK _6241_/D fanout166/X vssd1 vssd1 vccd1 vccd1 _6241_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA__4300__A _4313_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6172_ _6412_/CLK _6172_/D vssd1 vssd1 vccd1 vccd1 _6172_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3170__A1 _3502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5123_ _5209_/B _5123_/B vssd1 vssd1 vccd1 vccd1 _5124_/B sky130_fd_sc_hd__xnor2_1
X_3384_ _3611_/A _4734_/B vssd1 vssd1 vccd1 vccd1 _3384_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__5830__S _5933_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5054_ _5054_/A _5054_/B vssd1 vssd1 vccd1 vccd1 _5054_/Y sky130_fd_sc_hd__nand2_1
X_4005_ hold9/X _4425_/A2 _5597_/B vssd1 vssd1 vccd1 vccd1 _4005_/X sky130_fd_sc_hd__o21a_1
XANTENNA__4446__S _4446_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4670__A1 _6244_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout178_A fanout181/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5956_ _5977_/S _5956_/B vssd1 vssd1 vccd1 vccd1 _5956_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_47_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5887_ _5887_/A _5926_/A vssd1 vssd1 vccd1 vccd1 _5888_/B sky130_fd_sc_hd__or2_1
X_4907_ _4809_/B _4906_/Y _4903_/X _4867_/B vssd1 vssd1 vccd1 vccd1 _4907_/X sky130_fd_sc_hd__o211a_1
X_4838_ _6322_/Q _5852_/S _4837_/X _5557_/S vssd1 vssd1 vccd1 vccd1 _4838_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_28_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4769_ _4772_/A _4772_/B _5272_/C _4769_/D vssd1 vssd1 vccd1 vccd1 _4769_/X sky130_fd_sc_hd__or4_2
XANTENNA__5922__B2 _5747_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5922__A1 _5932_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6439_ _6448_/CLK _6439_/D fanout181/X vssd1 vssd1 vccd1 vccd1 _6439_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_0_101_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3697__C1 _5518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold32 hold32/A vssd1 vssd1 vccd1 vccd1 hold32/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 hold21/A vssd1 vssd1 vccd1 vccd1 hold21/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold10 hold10/A vssd1 vssd1 vccd1 vccd1 hold10/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 hold43/A vssd1 vssd1 vccd1 vccd1 hold43/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 hold54/A vssd1 vssd1 vccd1 vccd1 hold54/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 hold65/A vssd1 vssd1 vccd1 vccd1 hold65/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold76 hold76/A vssd1 vssd1 vccd1 vccd1 hold76/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4356__S _4360_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold87 hold87/A vssd1 vssd1 vccd1 vccd1 hold87/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold98 hold98/A vssd1 vssd1 vccd1 vccd1 hold98/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_7 _6274_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5429__B1 _5371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_23_wb_clk_i _6404_/CLK vssd1 vssd1 vccd1 vccd1 _6291_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_16_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4652__A1 _5715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xci2406_z80_200 vssd1 vssd1 vccd1 vccd1 ci2406_z80_200/HI io_oeb[19] sky130_fd_sc_hd__conb_1
Xci2406_z80_211 vssd1 vssd1 vccd1 vccd1 io_oeb[30] ci2406_z80_211/LO sky130_fd_sc_hd__conb_1
XFILLER_0_76_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5810_ _6376_/Q _5810_/B vssd1 vssd1 vccd1 vccd1 _5811_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_91_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6117__RESET_B fanout173/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5741_ _5931_/S _5932_/S _5731_/X vssd1 vssd1 vccd1 vccd1 _5742_/A sky130_fd_sc_hd__a21oi_4
XFILLER_0_29_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5672_ _6413_/Q _6313_/Q _4384_/S _6182_/Q _3721_/Y vssd1 vssd1 vccd1 vccd1 _5674_/A
+ sky130_fd_sc_hd__o221a_1
X_4623_ input3/X _4631_/B vssd1 vssd1 vccd1 vccd1 _4623_/X sky130_fd_sc_hd__and2_1
X_4554_ _3549_/A _4211_/C _3725_/B vssd1 vssd1 vccd1 vccd1 _4554_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_12_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold502 _6364_/Q vssd1 vssd1 vccd1 vccd1 hold502/X sky130_fd_sc_hd__dlygate4sd3_1
X_3505_ _3505_/A _3505_/B vssd1 vssd1 vccd1 vccd1 _3505_/Y sky130_fd_sc_hd__nand2_1
Xhold524 _6330_/Q vssd1 vssd1 vccd1 vccd1 _5514_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold513 _5529_/X vssd1 vssd1 vccd1 vccd1 _6331_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold535 _5721_/X vssd1 vssd1 vccd1 vccd1 _6365_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5126__A _6292_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6224_ _6305_/CLK _6224_/D fanout179/X vssd1 vssd1 vccd1 vccd1 _6224_/Q sky130_fd_sc_hd__dfrtp_1
Xhold557 _3644_/Y vssd1 vssd1 vccd1 vccd1 _6394_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold546 _5948_/X vssd1 vssd1 vccd1 vccd1 _6391_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold568 _6317_/Q vssd1 vssd1 vccd1 vccd1 _3363_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4485_ hold274/X _4380_/X _4491_/S vssd1 vssd1 vccd1 vccd1 _4485_/X sky130_fd_sc_hd__mux2_1
Xhold579 _6320_/Q vssd1 vssd1 vccd1 vccd1 hold579/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3436_ _5518_/S _3436_/B _3438_/S vssd1 vssd1 vccd1 vccd1 _3436_/X sky130_fd_sc_hd__and3_1
XFILLER_0_0_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3367_ _3658_/B _3367_/B vssd1 vssd1 vccd1 vccd1 _3426_/B sky130_fd_sc_hd__nand2_1
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6155_ _6218_/CLK _6155_/D vssd1 vssd1 vccd1 vccd1 _6155_/Q sky130_fd_sc_hd__dfxtp_1
X_6086_ _6204_/CLK _6086_/D fanout174/X vssd1 vssd1 vccd1 vccd1 _6086_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__4684__B _5553_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5106_ hold669/X _5105_/X _5447_/S vssd1 vssd1 vccd1 vccd1 _6292_/D sky130_fd_sc_hd__mux2_1
X_3298_ _3344_/A _3297_/X _3296_/X vssd1 vssd1 vccd1 vccd1 _3299_/C sky130_fd_sc_hd__o21a_1
X_5037_ _6385_/Q _6333_/Q _6315_/Q vssd1 vssd1 vccd1 vccd1 _5037_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4643__A1 _6337_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3446__A2 _3443_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3749__A3 _5715_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5939_ _5265_/A _3623_/A _3625_/B _5938_/X vssd1 vssd1 vccd1 vccd1 _6387_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_63_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3906__A0 _6417_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput33 _6288_/Q vssd1 vssd1 vccd1 vccd1 io_out[19] sky130_fd_sc_hd__buf_12
XANTENNA__4006__S0 _5676_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput22 _6487_/A vssd1 vssd1 vccd1 vccd1 io_oeb[29] sky130_fd_sc_hd__buf_12
XANTENNA__5659__B1 _5676_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput44 _6259_/Q vssd1 vssd1 vccd1 vccd1 io_out[29] sky130_fd_sc_hd__buf_12
XFILLER_0_9_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5470__S _5560_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4594__B _4604_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5831__B1 _5735_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6281__RESET_B fanout169/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4270_ _4747_/C _4270_/B vssd1 vssd1 vccd1 vccd1 _5563_/C sky130_fd_sc_hd__nor2_1
X_3221_ _4257_/B _3566_/B vssd1 vssd1 vccd1 vccd1 _4346_/A sky130_fd_sc_hd__or2_2
XANTENNA__4322__B1 _4323_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3676__A2 _5578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3152_ _3152_/A _3373_/A vssd1 vssd1 vccd1 vccd1 _3152_/Y sky130_fd_sc_hd__nand2_1
X_3083_ _3083_/A vssd1 vssd1 vccd1 vccd1 _6406_/D sky130_fd_sc_hd__inv_2
XANTENNA__3428__A2 _4734_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4724__S _5240_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3848__B _3862_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3985_ _3985_/A _5211_/B vssd1 vssd1 vccd1 vccd1 _3985_/X sky130_fd_sc_hd__and2_1
XFILLER_0_45_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5724_ _6274_/Q hold157/X _5724_/S vssd1 vssd1 vccd1 vccd1 _5724_/X sky130_fd_sc_hd__mux2_1
X_5655_ _6383_/Q _5600_/X _5652_/X _5594_/Y vssd1 vssd1 vccd1 vccd1 _5655_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_32_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4606_ _6440_/Q _4567_/Y _4568_/X _6448_/Q _4605_/X vssd1 vssd1 vccd1 vccd1 _4606_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4679__B _5560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold310 _6259_/Q vssd1 vssd1 vccd1 vccd1 hold310/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5586_ _5691_/S vssd1 vssd1 vccd1 vccd1 _5603_/D sky130_fd_sc_hd__inv_2
Xhold332 _6266_/Q vssd1 vssd1 vccd1 vccd1 hold332/X sky130_fd_sc_hd__dlygate4sd3_1
X_4537_ hold478/X _6296_/Q _4539_/S vssd1 vssd1 vccd1 vccd1 _4537_/X sky130_fd_sc_hd__mux2_1
Xhold321 _6077_/Q vssd1 vssd1 vccd1 vccd1 hold321/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold343 _6344_/Q vssd1 vssd1 vccd1 vccd1 _3079_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold354 _5698_/X vssd1 vssd1 vccd1 vccd1 _5699_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold376 _5621_/X vssd1 vssd1 vccd1 vccd1 _6337_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4468_ _4392_/X hold43/X _4473_/S vssd1 vssd1 vccd1 vccd1 hold44/A sky130_fd_sc_hd__mux2_1
Xhold365 _6338_/Q vssd1 vssd1 vccd1 vccd1 _3061_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_7_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold387 _6442_/Q vssd1 vssd1 vccd1 vccd1 hold387/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_3419_ _5324_/A _3297_/X _3661_/A _4318_/B _5322_/D vssd1 vssd1 vccd1 vccd1 _3419_/X
+ sky130_fd_sc_hd__a2111o_1
X_6207_ _6344_/CLK _6207_/D vssd1 vssd1 vccd1 vccd1 _6207_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold398 _5716_/X vssd1 vssd1 vccd1 vccd1 _6360_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6138_ _6194_/CLK _6138_/D vssd1 vssd1 vccd1 vccd1 _6138_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4864__A1 _6324_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4399_ _4427_/S _4398_/X _4397_/X vssd1 vssd1 vccd1 vccd1 _4399_/X sky130_fd_sc_hd__a21o_2
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6069_ _6181_/CLK _6069_/D vssd1 vssd1 vccd1 vccd1 _6069_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4092__A2 _3715_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5592__A2 _4382_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4855__A1 _6323_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5280__A1 _3656_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3830__A2 _3715_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6044__B _6063_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3770_ _3770_/A _6390_/Q _6391_/Q vssd1 vssd1 vccd1 vccd1 _3772_/B sky130_fd_sc_hd__or3b_2
XFILLER_0_13_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5440_ _5440_/A _5440_/B vssd1 vssd1 vccd1 vccd1 _5441_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5371_ _5371_/A _5441_/A vssd1 vssd1 vccd1 vccd1 _5371_/Y sky130_fd_sc_hd__nand2_1
X_4322_ _5058_/S _4323_/B _4323_/A vssd1 vssd1 vccd1 vccd1 _4322_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_10_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4253_ _5578_/A _3426_/A _4209_/Y vssd1 vssd1 vccd1 vccd1 _5563_/B sky130_fd_sc_hd__a21o_1
Xfanout119 hold612/X vssd1 vssd1 vccd1 vccd1 _5339_/A sky130_fd_sc_hd__buf_4
Xfanout108 _5347_/A vssd1 vssd1 vccd1 vccd1 _5447_/S sky130_fd_sc_hd__buf_6
XANTENNA__4719__S _4731_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3204_ _3290_/B _4679_/D vssd1 vssd1 vccd1 vccd1 _3599_/A sky130_fd_sc_hd__nor2_1
X_4184_ _4679_/A _6248_/Q _3216_/A _4183_/Y vssd1 vssd1 vccd1 vccd1 _4184_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_38_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3135_ _3289_/A _3573_/A _3534_/A vssd1 vssd1 vccd1 vccd1 _3135_/X sky130_fd_sc_hd__or3_1
X_3066_ _3066_/A vssd1 vssd1 vccd1 vccd1 _5347_/B sky130_fd_sc_hd__inv_2
XANTENNA__4454__S _4455_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3821__A2 _3779_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5023__A1 _5061_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3968_ _3970_/A _3970_/B vssd1 vssd1 vccd1 vccd1 _3969_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_92_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5023__B2 _4867_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5707_ _5707_/A vssd1 vssd1 vccd1 vccd1 _6352_/D sky130_fd_sc_hd__inv_2
X_3899_ _6243_/Q _6244_/Q _6245_/Q vssd1 vssd1 vccd1 vccd1 _4071_/C sky130_fd_sc_hd__o21a_1
XANTENNA__3594__A _3594_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5638_ _5638_/A _5638_/B vssd1 vssd1 vccd1 vccd1 _5638_/X sky130_fd_sc_hd__or2_1
X_5569_ _5603_/C vssd1 vssd1 vccd1 vccd1 _5602_/B sky130_fd_sc_hd__inv_2
XFILLER_0_13_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold140 _6158_/Q vssd1 vssd1 vccd1 vccd1 hold140/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold162 _4505_/X vssd1 vssd1 vccd1 vccd1 _6210_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold151 _6214_/Q vssd1 vssd1 vccd1 vccd1 hold151/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 _6224_/Q vssd1 vssd1 vccd1 vccd1 _4616_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold184 _4450_/X vssd1 vssd1 vccd1 vccd1 _6154_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 _6106_/Q vssd1 vssd1 vccd1 vccd1 hold173/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3760__C _6304_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6039__B1 _6063_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4065__A2 _6247_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3769__A _4224_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold637_A _6416_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3488__B _5975_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4773__B1 _4639_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3500__A1 _4214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3264__B1 _3654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4940_ _6442_/Q _5056_/A2 _4939_/X vssd1 vssd1 vccd1 vccd1 _4940_/X sky130_fd_sc_hd__a21o_1
XANTENNA__3803__A2 _3715_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5005__A1 _5061_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4871_ _6421_/Q _4758_/X _4869_/X _5061_/A1 vssd1 vssd1 vccd1 vccd1 _4871_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_46_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5005__B2 _4867_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3822_ _6132_/Q _3789_/X _3791_/X _6411_/Q vssd1 vssd1 vccd1 vccd1 _3822_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3567__A1 _6293_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5556__A2 _5377_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3753_ _4679_/A _6243_/Q _3752_/X vssd1 vssd1 vccd1 vccd1 _5130_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_27_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3684_ _3686_/A _5518_/S _3686_/C vssd1 vssd1 vccd1 vccd1 _3684_/X sky130_fd_sc_hd__and3_1
XANTENNA__3319__A1 _4637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5423_ _5450_/A _5422_/B _5422_/C vssd1 vssd1 vccd1 vccd1 _5424_/B sky130_fd_sc_hd__a21o_1
X_5354_ _5354_/A _5354_/B vssd1 vssd1 vccd1 vccd1 _5354_/X sky130_fd_sc_hd__or2_1
X_4305_ _6271_/Q _4304_/Y _4305_/S vssd1 vssd1 vccd1 vccd1 _4305_/X sky130_fd_sc_hd__mux2_1
X_5285_ _5275_/X _5283_/A _5284_/X hold113/X _5560_/B vssd1 vssd1 vccd1 vccd1 _5285_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_10_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4449__S _4455_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4819__A1 _5054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4236_ _4222_/B _4217_/X _4234_/X _4235_/X vssd1 vssd1 vccd1 vccd1 _4236_/X sky130_fd_sc_hd__o31a_1
XFILLER_0_4_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4167_ _3741_/X _4164_/X _4166_/B _4166_/Y _5087_/B vssd1 vssd1 vccd1 vccd1 _4167_/X
+ sky130_fd_sc_hd__a32o_1
X_3118_ _4744_/A _3183_/B _4744_/B vssd1 vssd1 vccd1 vccd1 _3220_/A sky130_fd_sc_hd__or3_4
XFILLER_0_65_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4047__A2 _6420_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4098_ _4098_/A _4098_/B vssd1 vssd1 vccd1 vccd1 _5253_/B sky130_fd_sc_hd__xnor2_1
X_3049_ _6401_/Q vssd1 vssd1 vccd1 vccd1 _3049_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_81_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3101__B _3254_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_47_wb_clk_i_A clkbuf_leaf_6_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__4867__B _4867_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4359__S _4360_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3099__A_N _4284_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_48_wb_clk_i clkbuf_leaf_6_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6354_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_64_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout90 _5784_/S vssd1 vssd1 vccd1 vccd1 _5849_/S sky130_fd_sc_hd__buf_4
XFILLER_0_36_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4841__S0 _5051_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5171__A0 _6270_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5455__A2_N _5377_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5070_ _5988_/B _5988_/C _6028_/A _5988_/A vssd1 vssd1 vccd1 vccd1 _5243_/S sky130_fd_sc_hd__or4b_4
XANTENNA__5474__A1 _4920_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4021_ _4021_/A _4021_/B vssd1 vssd1 vccd1 vccd1 _4022_/B sky130_fd_sc_hd__nor2_1
X_5972_ input2/X hold645/X _5975_/S vssd1 vssd1 vccd1 vccd1 _6420_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_59_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5777__A2 _6419_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4923_ _6379_/Q _6327_/Q _6315_/Q vssd1 vssd1 vccd1 vccd1 _4923_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5828__S _5931_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4732__S _4732_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4854_ _6323_/Q _4752_/X _4852_/X _4853_/X vssd1 vssd1 vccd1 vccd1 _4854_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_74_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4785_ _6161_/Q _6408_/Q hold67/A _6177_/Q _4326_/B _5358_/A0 vssd1 vssd1 vccd1 vccd1
+ _4785_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_7_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4201__A2 _4198_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3805_ _4111_/A _3805_/B vssd1 vssd1 vccd1 vccd1 _4423_/A sky130_fd_sc_hd__xnor2_1
X_3736_ _3938_/A _3735_/X _3736_/S vssd1 vssd1 vccd1 vccd1 _3738_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_55_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3667_ _3224_/X _4745_/B _5096_/B vssd1 vssd1 vccd1 vccd1 _3668_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_42_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3598_ _4522_/B _3600_/B _3600_/C vssd1 vssd1 vccd1 vccd1 _4743_/C sky130_fd_sc_hd__a21o_1
X_6386_ _6386_/CLK _6386_/D fanout166/X vssd1 vssd1 vccd1 vccd1 _6386_/Q sky130_fd_sc_hd__dfrtp_4
X_5406_ _5715_/A _6419_/Q vssd1 vssd1 vccd1 vccd1 _5408_/B sky130_fd_sc_hd__or2_1
XFILLER_0_100_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3712__A1 _3473_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5337_ _4568_/B _5332_/Y _5977_/S vssd1 vssd1 vccd1 vccd1 _5337_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_11_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5268_ _4224_/A _3572_/A _5266_/X _5267_/X _3574_/B vssd1 vssd1 vccd1 vccd1 _5268_/X
+ sky130_fd_sc_hd__a221o_1
X_4219_ _3254_/A _6118_/Q _3530_/D _4218_/X vssd1 vssd1 vccd1 vccd1 _4219_/X sky130_fd_sc_hd__a22o_1
X_5199_ _3759_/A _5196_/X _5198_/X vssd1 vssd1 vccd1 vccd1 _5199_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__3476__B1 _4309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3112__A _3254_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4728__B1 _5075_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4823__S0 _5358_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_3_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3703__A1 _3473_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5456__A1 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6436__SET_B fanout171/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6052__B _6063_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4570_ _4604_/S _4570_/B vssd1 vssd1 vccd1 vccd1 _4570_/X sky130_fd_sc_hd__and2_2
XFILLER_0_4_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3521_ _3600_/A _5291_/A _3521_/C _3521_/D vssd1 vssd1 vccd1 vccd1 _3521_/X sky130_fd_sc_hd__or4_1
XFILLER_0_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4788__A _5058_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3452_ _3469_/A _3452_/B vssd1 vssd1 vccd1 vccd1 _3453_/B sky130_fd_sc_hd__nor2_1
X_6240_ _6297_/CLK _6240_/D fanout176/X vssd1 vssd1 vccd1 vccd1 _6240_/Q sky130_fd_sc_hd__dfstp_1
X_3383_ _3657_/A _3418_/B vssd1 vssd1 vccd1 vccd1 _3394_/C sky130_fd_sc_hd__and2_1
X_6171_ _6410_/CLK _6171_/D vssd1 vssd1 vccd1 vccd1 _6171_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5695__A1 _5695_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3170__A2 _4222_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5122_ _5122_/A _5219_/B vssd1 vssd1 vccd1 vccd1 _5124_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_41_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5053_ _5052_/X _5051_/X _5053_/S vssd1 vssd1 vccd1 vccd1 _5054_/B sky130_fd_sc_hd__mux2_2
XANTENNA__4727__S _4727_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4004_ _3724_/A _5253_/A _3995_/Y vssd1 vssd1 vccd1 vccd1 _4004_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_79_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5955_ _4616_/A _3639_/C _3641_/B vssd1 vssd1 vccd1 vccd1 _5955_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_1_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5886_ _5887_/A _5926_/A vssd1 vssd1 vccd1 vccd1 _5888_/A sky130_fd_sc_hd__nand2_1
XANTENNA__4462__S _4464_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4906_ _4943_/C vssd1 vssd1 vccd1 vccd1 _4906_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_47_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4837_ _5773_/A _4836_/X _4826_/X vssd1 vssd1 vccd1 vccd1 _4837_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_90_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4805__S0 _5358_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4768_ _4768_/A _4768_/B vssd1 vssd1 vccd1 vccd1 _4769_/D sky130_fd_sc_hd__nand2_1
X_3719_ _6335_/Q _5597_/B vssd1 vssd1 vccd1 vccd1 _3719_/X sky130_fd_sc_hd__or2_1
X_4699_ _6269_/Q _4681_/X _4698_/X _5371_/A vssd1 vssd1 vccd1 vccd1 _4699_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_101_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6438_ _6445_/CLK _6438_/D fanout171/X vssd1 vssd1 vccd1 vccd1 _6438_/Q sky130_fd_sc_hd__dfstp_2
XANTENNA__4210__B _5258_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5686__A1 _6274_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3107__A _5258_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6369_ _6430_/CLK hold36/X vssd1 vssd1 vccd1 vccd1 hold35/A sky130_fd_sc_hd__dfxtp_1
Xhold22 hold22/A vssd1 vssd1 vccd1 vccd1 hold22/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold11 hold11/A vssd1 vssd1 vccd1 vccd1 hold11/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 hold33/A vssd1 vssd1 vccd1 vccd1 hold33/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 hold55/A vssd1 vssd1 vccd1 vccd1 hold55/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 hold44/A vssd1 vssd1 vccd1 vccd1 hold44/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 hold77/A vssd1 vssd1 vccd1 vccd1 hold77/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 hold99/A vssd1 vssd1 vccd1 vccd1 hold99/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 hold88/A vssd1 vssd1 vccd1 vccd1 hold88/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 hold66/A vssd1 vssd1 vccd1 vccd1 hold66/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5992__A _6054_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_8 _6117_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5931__S _5931_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5429__A1 _5441_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5589__D _5691_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xci2406_z80_201 vssd1 vssd1 vccd1 vccd1 ci2406_z80_201/HI io_oeb[20] sky130_fd_sc_hd__conb_1
Xci2406_z80_212 vssd1 vssd1 vccd1 vccd1 io_oeb[31] ci2406_z80_212/LO sky130_fd_sc_hd__conb_1
XFILLER_0_76_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5740_ _5740_/A _5746_/B vssd1 vssd1 vccd1 vccd1 _5815_/S sky130_fd_sc_hd__nor2_2
XFILLER_0_8_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5671_ _5695_/A1 _4056_/A _5571_/Y _5670_/X vssd1 vssd1 vccd1 vccd1 _5671_/X sky130_fd_sc_hd__a22o_1
X_4622_ _4744_/B _4615_/X _4617_/Y _4621_/X vssd1 vssd1 vccd1 vccd1 _6253_/D sky130_fd_sc_hd__o22a_1
XFILLER_0_72_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4553_ _3549_/A _3511_/A _4767_/B _4550_/Y _4552_/X vssd1 vssd1 vccd1 vccd1 _4553_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_0_13_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold514 _6255_/Q vssd1 vssd1 vccd1 vccd1 hold514/X sky130_fd_sc_hd__dlygate4sd3_1
X_3504_ hold249/X _3503_/X _5472_/S vssd1 vssd1 vccd1 vccd1 _3504_/X sky130_fd_sc_hd__mux2_1
X_4484_ hold105/X _4367_/X _4491_/S vssd1 vssd1 vccd1 vccd1 _4484_/X sky130_fd_sc_hd__mux2_1
Xhold525 _5517_/X vssd1 vssd1 vccd1 vccd1 _6330_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold503 _5720_/X vssd1 vssd1 vccd1 vccd1 _6364_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold536 _6440_/Q vssd1 vssd1 vccd1 vccd1 hold536/X sky130_fd_sc_hd__dlygate4sd3_1
X_6223_ _6403_/CLK _6223_/D fanout179/X vssd1 vssd1 vccd1 vccd1 _6223_/Q sky130_fd_sc_hd__dfrtp_1
X_3435_ _3438_/S vssd1 vssd1 vccd1 vccd1 _3435_/Y sky130_fd_sc_hd__inv_2
Xhold569 _5356_/X vssd1 vssd1 vccd1 vccd1 _6317_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold547 _6383_/Q vssd1 vssd1 vccd1 vccd1 _5887_/A sky130_fd_sc_hd__buf_1
Xhold558 _6329_/Q vssd1 vssd1 vccd1 vccd1 hold558/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5668__A1 _6384_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3366_ _5061_/A1 _3362_/X _4279_/A vssd1 vssd1 vccd1 vccd1 _4901_/S sky130_fd_sc_hd__o21ai_4
X_6154_ _6194_/CLK _6154_/D vssd1 vssd1 vccd1 vccd1 _6154_/Q sky130_fd_sc_hd__dfxtp_1
X_3297_ _3573_/A _4541_/A _4541_/C vssd1 vssd1 vccd1 vccd1 _3297_/X sky130_fd_sc_hd__and3_2
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5105_ _3909_/Y _5098_/A _5098_/Y _5104_/X vssd1 vssd1 vccd1 vccd1 _5105_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4457__S _4464_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6085_ _6433_/CLK _6085_/D vssd1 vssd1 vccd1 vccd1 _6085_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5036_ _6447_/Q _5056_/A2 _5035_/X vssd1 vssd1 vccd1 vccd1 _5036_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5938_ hold565/X _5949_/B _5936_/Y _5937_/Y _3625_/A vssd1 vssd1 vccd1 vccd1 _5938_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__6123__D _6127_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5869_ _5889_/A _5869_/B vssd1 vssd1 vccd1 vccd1 _5869_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4221__A _4637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5317__A _5317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput23 _4732_/S vssd1 vssd1 vccd1 vccd1 io_out[0] sky130_fd_sc_hd__buf_12
Xoutput34 _6415_/Q vssd1 vssd1 vccd1 vccd1 io_out[1] sky130_fd_sc_hd__buf_12
XFILLER_0_31_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput45 _3648_/X vssd1 vssd1 vccd1 vccd1 io_out[2] sky130_fd_sc_hd__buf_12
XANTENNA_hold667_A _6313_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5831__A1 _5236_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3300__A _3656_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6250__RESET_B fanout179/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3220_ _3220_/A _3566_/B vssd1 vssd1 vccd1 vccd1 _5097_/B sky130_fd_sc_hd__or2_4
XANTENNA__4322__A1 _5058_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3151_ _3152_/A _3373_/A vssd1 vssd1 vccd1 vccd1 _3232_/C sky130_fd_sc_hd__and2_1
X_3082_ _3082_/A vssd1 vssd1 vccd1 vccd1 _6404_/D sky130_fd_sc_hd__inv_2
XFILLER_0_89_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3984_ _6244_/Q _6246_/Q _4135_/S vssd1 vssd1 vccd1 vccd1 _5211_/B sky130_fd_sc_hd__mux2_1
XANTENNA__3210__A _4284_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5723_ _6274_/Q hold560/X _5723_/S vssd1 vssd1 vccd1 vccd1 _5723_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_72_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5654_ _6437_/Q _5588_/X _5603_/X _6375_/Q _5653_/X vssd1 vssd1 vccd1 vccd1 _5657_/A
+ sky130_fd_sc_hd__a221o_1
X_4605_ _6423_/Q _4569_/X _4570_/X _6274_/Q vssd1 vssd1 vccd1 vccd1 _4605_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4561__A1 _3183_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5585_ _3183_/B _5573_/X _5584_/X _5952_/A vssd1 vssd1 vccd1 vccd1 _5691_/S sky130_fd_sc_hd__a22o_4
Xhold311 _4642_/X vssd1 vssd1 vccd1 vccd1 _6259_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold300 _6411_/Q vssd1 vssd1 vccd1 vccd1 hold300/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold333 _4677_/X vssd1 vssd1 vccd1 vccd1 _6266_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold344 _6263_/Q vssd1 vssd1 vccd1 vccd1 hold344/X sky130_fd_sc_hd__dlygate4sd3_1
X_4536_ hold482/X _6295_/Q _4539_/S vssd1 vssd1 vccd1 vccd1 _4536_/X sky130_fd_sc_hd__mux2_1
Xhold322 _4282_/X vssd1 vssd1 vccd1 vccd1 _6077_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold355 _6264_/Q vssd1 vssd1 vccd1 vccd1 hold355/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold366 _5632_/X vssd1 vssd1 vccd1 vccd1 _6338_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4467_ _4380_/X hold67/X _4473_/S vssd1 vssd1 vccd1 vccd1 hold68/A sky130_fd_sc_hd__mux2_1
XANTENNA__4976__A _5054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold377 _6361_/Q vssd1 vssd1 vccd1 vccd1 hold377/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6206_ _6397_/CLK _6206_/D fanout174/X vssd1 vssd1 vccd1 vccd1 _6206_/Q sky130_fd_sc_hd__dfrtp_1
X_3418_ _3418_/A _3418_/B vssd1 vssd1 vccd1 vccd1 _3418_/Y sky130_fd_sc_hd__nor2_1
Xhold388 _6037_/X vssd1 vssd1 vccd1 vccd1 _6442_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold399 _6445_/Q vssd1 vssd1 vccd1 vccd1 hold399/X sky130_fd_sc_hd__buf_1
X_4398_ hold181/X hold59/X hold285/X hold41/X _5673_/C1 _4384_/S vssd1 vssd1 vccd1
+ vccd1 _4398_/X sky130_fd_sc_hd__mux4_2
X_3349_ _3349_/A _3349_/B _3348_/X vssd1 vssd1 vccd1 vccd1 _3349_/X sky130_fd_sc_hd__or3b_1
X_6137_ _6217_/CLK _6137_/D vssd1 vssd1 vccd1 vccd1 _6137_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4864__A2 _4752_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6068_ _6221_/CLK _6068_/D vssd1 vssd1 vccd1 vccd1 _6068_/Q sky130_fd_sc_hd__dfxtp_1
X_5019_ _6384_/Q _6332_/Q _6315_/Q vssd1 vssd1 vccd1 vccd1 _5019_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4915__S _5029_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5600__A _5603_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6079__RESET_B fanout169/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4552__B2 _5733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4068__B1 _5217_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5804__A1 _6324_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3815__B1 _3791_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4825__S _5053_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6431__RESET_B fanout178/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4126__A _6248_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3684__B _5518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4543__A1 _5096_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5370_ _6392_/Q _5518_/S vssd1 vssd1 vccd1 vccd1 _5377_/A sky130_fd_sc_hd__nand2_4
XFILLER_0_22_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4321_ _4321_/A _4321_/B vssd1 vssd1 vccd1 vccd1 _4323_/B sky130_fd_sc_hd__nand2_1
X_4252_ _4228_/A _3654_/A _5323_/C _4251_/X vssd1 vssd1 vccd1 vccd1 _4252_/X sky130_fd_sc_hd__a31o_1
XANTENNA__5099__A2 _6292_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout109 _4732_/S vssd1 vssd1 vccd1 vccd1 _5347_/A sky130_fd_sc_hd__buf_4
XFILLER_0_10_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3203_ _5322_/A _5292_/A vssd1 vssd1 vccd1 vccd1 _3281_/A sky130_fd_sc_hd__or2_1
X_4183_ _4679_/A _4183_/B vssd1 vssd1 vccd1 vccd1 _4183_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3134_ _3091_/X _3116_/X _3125_/X _3133_/X vssd1 vssd1 vccd1 vccd1 _3197_/A sky130_fd_sc_hd__o211ai_1
X_3065_ _6295_/Q vssd1 vssd1 vccd1 vccd1 _3065_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3806__B1 _3786_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5420__A _5715_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3967_ _5088_/B _6339_/Q vssd1 vssd1 vccd1 vccd1 _3970_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_70_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4470__S _4473_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5706_ _3078_/Y _3798_/B _6060_/S vssd1 vssd1 vccd1 vccd1 _5707_/A sky130_fd_sc_hd__mux2_1
X_3898_ _3896_/S _3746_/X _3895_/X _3897_/X vssd1 vssd1 vccd1 vccd1 _3898_/X sky130_fd_sc_hd__a211o_1
XANTENNA__3594__B _5733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5637_ _6094_/Q _4382_/B _4200_/S _6139_/Q _5673_/C1 vssd1 vssd1 vccd1 vccd1 _5638_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_79_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4534__A1 _6293_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5568_ _5935_/A _5568_/B vssd1 vssd1 vccd1 vccd1 _5603_/C sky130_fd_sc_hd__nor2_2
XANTENNA__5731__B1 _3477_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4519_ _4767_/A _4520_/B vssd1 vssd1 vccd1 vccd1 _5075_/B sky130_fd_sc_hd__and2_4
XANTENNA_clkbuf_leaf_37_wb_clk_i_A clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold141 _6189_/Q vssd1 vssd1 vccd1 vccd1 hold141/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold152 _4509_/X vssd1 vssd1 vccd1 vccd1 _6214_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold130 _6409_/Q vssd1 vssd1 vccd1 vccd1 hold130/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold185 _6137_/Q vssd1 vssd1 vccd1 vccd1 hold185/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold163 _6111_/Q vssd1 vssd1 vccd1 vccd1 hold163/X sky130_fd_sc_hd__dlygate4sd3_1
X_5499_ _6443_/Q _4958_/B _5518_/S vssd1 vssd1 vccd1 vccd1 _5501_/B sky130_fd_sc_hd__mux2_1
Xhold174 _4345_/X vssd1 vssd1 vccd1 vccd1 _6106_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold196 _3539_/X vssd1 vssd1 vccd1 vccd1 _6224_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6039__A1 _6057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold365_A _6338_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5262__A2 _5578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4065__A3 _6341_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3769__B _5322_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold532_A _6248_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5970__A0 input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4525__A1 _6268_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5722__A0 _6273_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3264__A1 _3611_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4870_ _6438_/Q _4756_/Y _4757_/Y _4863_/B _4754_/X vssd1 vssd1 vccd1 vccd1 _4870_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_74_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3821_ hold93/A _3779_/X _3781_/X hold61/A _3820_/X vssd1 vssd1 vccd1 vccd1 _3824_/A
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3567__A2 _5158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3752_ _5217_/A _3216_/A _3751_/X _3525_/B _4135_/S vssd1 vssd1 vccd1 vccd1 _3752_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_6_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3683_ _4767_/A _3683_/B _3683_/C vssd1 vssd1 vccd1 vccd1 _3687_/B sky130_fd_sc_hd__and3_2
XFILLER_0_2_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5422_ _5450_/A _5422_/B _5422_/C vssd1 vssd1 vccd1 vccd1 _5422_/X sky130_fd_sc_hd__and3_1
X_5353_ _5353_/A _5353_/B vssd1 vssd1 vccd1 vccd1 _6315_/D sky130_fd_sc_hd__or2_1
XFILLER_0_49_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4304_ _4304_/A _4304_/B vssd1 vssd1 vccd1 vccd1 _4304_/Y sky130_fd_sc_hd__nor2_1
X_5284_ _6389_/Q _6117_/Q _5347_/A vssd1 vssd1 vccd1 vccd1 _5284_/X sky130_fd_sc_hd__and3_1
XANTENNA__4819__A2 _4807_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4235_ _6256_/Q _3952_/B _4211_/C _3725_/B vssd1 vssd1 vccd1 vccd1 _4235_/X sky130_fd_sc_hd__a31o_1
X_4166_ _5087_/A _4166_/B vssd1 vssd1 vccd1 vccd1 _4166_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_4_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3117_ _3254_/A _3183_/B vssd1 vssd1 vccd1 vccd1 _3289_/C sky130_fd_sc_hd__nor2_1
XANTENNA__5150__A _6304_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4097_ _4022_/A _4022_/B _4021_/A vssd1 vssd1 vccd1 vccd1 _4098_/B sky130_fd_sc_hd__a21oi_1
X_3048_ _5728_/A vssd1 vssd1 vccd1 vccd1 _3048_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_77_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4999_ _6383_/Q _6331_/Q _6315_/Q vssd1 vssd1 vccd1 vccd1 _4999_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_33_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4691__B1 _5075_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5943__B1 _5096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout91 _5029_/S vssd1 vssd1 vccd1 vccd1 _5557_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_0_24_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout80 _4319_/X vssd1 vssd1 vccd1 vccd1 _5054_/A sky130_fd_sc_hd__buf_4
XFILLER_0_64_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4841__S1 _5052_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_17_wb_clk_i _6404_/CLK vssd1 vssd1 vccd1 vccd1 _6401_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_101_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3721__A2 _4382_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4020_ _4111_/A _4020_/B vssd1 vssd1 vccd1 vccd1 _4021_/B sky130_fd_sc_hd__nor2_1
XANTENNA__4793__B _4867_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5971_ input3/X hold641/X _5975_/S vssd1 vssd1 vccd1 vccd1 _6419_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_47_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4985__A1 _5061_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5777__A3 _3580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4922_ _6441_/Q _5056_/A2 _4921_/X vssd1 vssd1 vccd1 vccd1 _4922_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_47_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4985__B2 _4867_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4853_ _6375_/Q _4796_/B _5927_/S vssd1 vssd1 vccd1 vccd1 _4853_/X sky130_fd_sc_hd__o21a_1
X_4784_ _6185_/Q hold75/A _6145_/Q hold57/A _4326_/B _5358_/A0 vssd1 vssd1 vccd1 vccd1
+ _4784_/X sky130_fd_sc_hd__mux4_1
X_3804_ _3804_/A _3804_/B _3804_/C vssd1 vssd1 vccd1 vccd1 _3805_/B sky130_fd_sc_hd__or3_2
X_3735_ _6301_/Q _3938_/A vssd1 vssd1 vccd1 vccd1 _3735_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_15_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5844__S _5933_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3666_ _3666_/A vssd1 vssd1 vccd1 vccd1 _4220_/B sky130_fd_sc_hd__inv_2
XANTENNA_fanout116_A _6427_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5405_ hold585/X _5404_/X _5447_/S vssd1 vssd1 vccd1 vccd1 _5405_/X sky130_fd_sc_hd__mux2_1
X_3597_ _3597_/A vssd1 vssd1 vccd1 vccd1 _3597_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_62_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6385_ _6386_/CLK _6385_/D fanout167/X vssd1 vssd1 vccd1 vccd1 _6385_/Q sky130_fd_sc_hd__dfrtp_4
X_5336_ _5988_/A _5335_/Y _5727_/S vssd1 vssd1 vccd1 vccd1 _5336_/X sky130_fd_sc_hd__mux2_1
X_5267_ _3572_/A _3770_/A _5317_/B _4224_/A vssd1 vssd1 vccd1 vccd1 _5267_/X sky130_fd_sc_hd__a211o_1
X_4218_ _3152_/A _5733_/A _3770_/A _4212_/X _4217_/X vssd1 vssd1 vccd1 vccd1 _4218_/X
+ sky130_fd_sc_hd__a311o_1
X_5198_ _3985_/A _5211_/D _5149_/X _6296_/Q _5197_/X vssd1 vssd1 vccd1 vccd1 _5198_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3476__A1 _5553_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4149_ _4148_/X hold197/X _4206_/S vssd1 vssd1 vccd1 vccd1 _6074_/D sky130_fd_sc_hd__mux2_1
XANTENNA__6126__D _6126_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4923__S _6315_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4224__A _4224_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4823__S1 _4326_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3782__B _3862_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6204__RESET_B fanout174/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4664__A0 _6337_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5613__C1 _5675_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3234__A4 _3566_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4134__A _4255_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3520_ _3520_/A _4734_/C _4541_/D _4347_/C vssd1 vssd1 vccd1 vccd1 _3521_/D sky130_fd_sc_hd__or4_1
XFILLER_0_97_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4788__B _4788_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5144__A1 _6337_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5144__B2 _6338_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3451_ _5935_/A _6392_/Q _3451_/C _5978_/A vssd1 vssd1 vccd1 vccd1 _3452_/B sky130_fd_sc_hd__or4_1
XFILLER_0_12_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3382_ _3337_/B _5480_/D _4541_/B vssd1 vssd1 vccd1 vccd1 _3418_/B sky130_fd_sc_hd__o21a_1
X_6170_ _6414_/CLK hold44/X vssd1 vssd1 vccd1 vccd1 hold43/A sky130_fd_sc_hd__dfxtp_1
X_5121_ _5121_/A _5121_/B vssd1 vssd1 vccd1 vccd1 _5125_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5052_ _6222_/Q _6159_/Q _6199_/Q _6075_/Q _5358_/A0 _5052_/S1 vssd1 vssd1 vccd1
+ vccd1 _5052_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4003_ _4009_/B _4003_/B vssd1 vssd1 vccd1 vccd1 _5253_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__4309__A _4309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3213__A _4228_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4028__B _6340_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5954_ _3467_/X _3621_/A _3625_/B hold621/X _5952_/Y vssd1 vssd1 vccd1 vccd1 _5954_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_0_87_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5885_ _5876_/A _5884_/X _5933_/S vssd1 vssd1 vccd1 vccd1 _5885_/X sky130_fd_sc_hd__mux2_1
X_4905_ _6321_/Q _6322_/Q _4905_/C _4905_/D vssd1 vssd1 vccd1 vccd1 _4943_/C sky130_fd_sc_hd__and4_2
XFILLER_0_47_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4836_ _6322_/Q _5825_/S _5850_/B1 _4835_/X vssd1 vssd1 vccd1 vccd1 _4836_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4805__S1 _4326_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4767_ _4767_/A _4767_/B _4767_/C vssd1 vssd1 vccd1 vccd1 _4768_/B sky130_fd_sc_hd__and3_1
XFILLER_0_7_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3718_ _6313_/Q _4382_/C vssd1 vssd1 vccd1 vccd1 _3718_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__6442__SET_B fanout171/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4698_ _6269_/Q _4680_/X _5075_/B hold451/X vssd1 vssd1 vccd1 vccd1 _4698_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_101_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3649_ _6127_/Q _6123_/Q input1/X vssd1 vssd1 vccd1 vccd1 _3649_/X sky130_fd_sc_hd__mux2_1
X_6437_ _6445_/CLK _6437_/D fanout171/X vssd1 vssd1 vccd1 vccd1 _6437_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_0_101_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6368_ _6368_/CLK _6368_/D fanout169/X vssd1 vssd1 vccd1 vccd1 _6368_/Q sky130_fd_sc_hd__dfrtp_1
X_5319_ _5715_/B hold623/X _5321_/S _5318_/X vssd1 vssd1 vccd1 vccd1 _6305_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_87_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3697__A1 _5096_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4894__A0 _6325_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6299_ _6399_/CLK _6299_/D vssd1 vssd1 vccd1 vccd1 _6299_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5603__A _5603_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold23 hold23/A vssd1 vssd1 vccd1 vccd1 hold23/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold12 hold12/A vssd1 vssd1 vccd1 vccd1 hold12/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 hold34/A vssd1 vssd1 vccd1 vccd1 hold34/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 hold56/A vssd1 vssd1 vccd1 vccd1 hold56/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 hold45/A vssd1 vssd1 vccd1 vccd1 hold45/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 hold67/A vssd1 vssd1 vccd1 vccd1 hold67/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 hold78/A vssd1 vssd1 vccd1 vccd1 hold78/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold89 hold89/A vssd1 vssd1 vccd1 vccd1 hold89/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold612_A _6402_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5374__B2 _5560_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_9 _4349_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4885__A0 _4882_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3033__A _3183_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xci2406_z80_202 vssd1 vssd1 vccd1 vccd1 ci2406_z80_202/HI io_oeb[21] sky130_fd_sc_hd__conb_1
XFILLER_0_16_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xci2406_z80_213 vssd1 vssd1 vccd1 vccd1 io_oeb[35] ci2406_z80_213/LO sky130_fd_sc_hd__conb_1
XFILLER_0_29_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3612__A1 _4309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_32_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6343_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_17_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5670_ _5670_/A _5670_/B vssd1 vssd1 vccd1 vccd1 _5670_/X sky130_fd_sc_hd__or2_1
X_4621_ input6/X _4631_/B vssd1 vssd1 vccd1 vccd1 _4621_/X sky130_fd_sc_hd__and2_1
XFILLER_0_72_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5394__S _5553_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4552_ _3549_/A _5324_/A _4551_/Y _5733_/A _4222_/B vssd1 vssd1 vccd1 vccd1 _4552_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_25_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3503_ _3530_/D _3500_/X _3537_/B _6118_/Q _3501_/Y vssd1 vssd1 vccd1 vccd1 _3503_/X
+ sky130_fd_sc_hd__a221o_1
Xhold515 _3569_/Y vssd1 vssd1 vccd1 vccd1 _6399_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold526 _6334_/Q vssd1 vssd1 vccd1 vccd1 hold526/X sky130_fd_sc_hd__dlygate4sd3_1
X_4483_ _4483_/A _5959_/B vssd1 vssd1 vccd1 vccd1 _4491_/S sky130_fd_sc_hd__nor2_4
Xhold504 _6377_/Q vssd1 vssd1 vccd1 vccd1 hold504/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3434_ _5935_/A _3434_/B _3434_/C _3433_/X vssd1 vssd1 vccd1 vccd1 _3438_/S sky130_fd_sc_hd__or4b_2
Xhold559 _5508_/X vssd1 vssd1 vccd1 vccd1 _6329_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold548 _5899_/X vssd1 vssd1 vccd1 vccd1 _6383_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6222_ _6444_/CLK _6222_/D vssd1 vssd1 vccd1 vccd1 _6222_/Q sky130_fd_sc_hd__dfxtp_1
Xhold537 _6027_/X vssd1 vssd1 vccd1 vccd1 _6440_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3679__A1 _3164_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4876__A0 _6324_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3365_ _3365_/A _3365_/B vssd1 vssd1 vccd1 vccd1 _4279_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_0_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6153_ _6217_/CLK _6153_/D vssd1 vssd1 vccd1 vccd1 _6153_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4628__B1 _4617_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3296_ _5578_/A _5258_/B _3233_/D vssd1 vssd1 vccd1 vccd1 _3296_/X sky130_fd_sc_hd__a21o_1
X_5104_ _5102_/Y _5103_/X _5099_/X vssd1 vssd1 vccd1 vccd1 _5104_/X sky130_fd_sc_hd__a21o_1
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6084_ _6368_/CLK _6084_/D fanout169/X vssd1 vssd1 vccd1 vccd1 _6084_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5035_ _6273_/Q _4758_/X _6057_/C _4757_/Y vssd1 vssd1 vccd1 vccd1 _5035_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_79_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4473__S _4473_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5937_ _5952_/A _5937_/B vssd1 vssd1 vccd1 vccd1 _5937_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_48_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4800__B1 _5728_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5868_ _5889_/A _5869_/B vssd1 vssd1 vccd1 vccd1 _5868_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_63_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5799_ _5773_/A _5798_/X _4844_/X vssd1 vssd1 vccd1 vccd1 _5799_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_35_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4819_ _5054_/A _4807_/X _5728_/D vssd1 vssd1 vccd1 vccd1 _4819_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_16_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5317__B _5317_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5659__A2 _4198_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput24 _6276_/Q vssd1 vssd1 vccd1 vccd1 io_out[10] sky130_fd_sc_hd__buf_12
XFILLER_0_101_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput46 _3048_/Y vssd1 vssd1 vccd1 vccd1 io_out[32] sky130_fd_sc_hd__buf_12
Xoutput35 _6289_/Q vssd1 vssd1 vccd1 vccd1 io_out[20] sky130_fd_sc_hd__buf_12
XANTENNA_fanout96_A _5740_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4648__S _4674_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5831__A2 _6423_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4709__A1_N _6271_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3150_ _6257_/Q _6258_/Q vssd1 vssd1 vccd1 vccd1 _3233_/D sky130_fd_sc_hd__nand2b_2
X_3081_ _5949_/C vssd1 vssd1 vccd1 vccd1 _3081_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_27_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4293__S _6064_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5035__B1 _6057_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3983_ _6339_/Q _6343_/Q _6301_/Q vssd1 vssd1 vccd1 vccd1 _5216_/D sky130_fd_sc_hd__mux2_1
XANTENNA__3210__B _5226_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5722_ _6273_/Q hold405/X _5723_/S vssd1 vssd1 vccd1 vccd1 _5722_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_84_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5653_ _6295_/Q _5587_/X _5602_/X _6420_/Q vssd1 vssd1 vccd1 vccd1 _5653_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_45_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6378__RESET_B fanout168/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5584_ _5584_/A1 _5576_/X _5583_/X _3530_/D vssd1 vssd1 vccd1 vccd1 _5584_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_60_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6307__RESET_B fanout173/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4604_ _4156_/B _3805_/B _4604_/S vssd1 vssd1 vccd1 vccd1 _4604_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4679__D _4679_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4535_ hold480/X _6294_/Q _4539_/S vssd1 vssd1 vccd1 vccd1 _4535_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_13_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold301 _6410_/Q vssd1 vssd1 vccd1 vccd1 hold301/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4561__A2 _5313_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold334 _6265_/Q vssd1 vssd1 vccd1 vccd1 hold334/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_27_wb_clk_i_A _6404_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold312 _6260_/Q vssd1 vssd1 vccd1 vccd1 hold312/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold323 _6081_/Q vssd1 vssd1 vccd1 vccd1 _4299_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold367 _6403_/Q vssd1 vssd1 vccd1 vccd1 _4609_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold356 _4667_/X vssd1 vssd1 vccd1 vccd1 _6264_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold345 _4662_/X vssd1 vssd1 vccd1 vccd1 _6263_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4466_ _4367_/X hold53/X _4473_/S vssd1 vssd1 vccd1 vccd1 hold54/A sky130_fd_sc_hd__mux2_1
Xhold378 _5717_/X vssd1 vssd1 vccd1 vccd1 _6361_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4849__A0 _4843_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6205_ _6397_/CLK hold48/X fanout174/X vssd1 vssd1 vccd1 vccd1 hold47/A sky130_fd_sc_hd__dfrtp_1
X_3417_ _4747_/D _3377_/Y _4541_/B vssd1 vssd1 vccd1 vccd1 _3417_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_68_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4468__S _4473_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold389 _6286_/Q vssd1 vssd1 vccd1 vccd1 hold389/X sky130_fd_sc_hd__dlygate4sd3_1
X_4397_ hold15/X _4425_/A2 _3995_/Y _4396_/Y _5597_/B vssd1 vssd1 vccd1 vccd1 _4397_/X
+ sky130_fd_sc_hd__o221a_1
X_3348_ _3418_/A _3657_/B _3346_/Y _3342_/X vssd1 vssd1 vccd1 vccd1 _3348_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6136_ _6221_/CLK _6136_/D vssd1 vssd1 vccd1 vccd1 _6136_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3279_ _3683_/C _3238_/C _4320_/B _3242_/B _5322_/D vssd1 vssd1 vccd1 vccd1 _3592_/A
+ sky130_fd_sc_hd__a2111o_1
X_5018_ _6446_/Q _5056_/A2 _5017_/X vssd1 vssd1 vccd1 vccd1 _5018_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_67_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5329__A1 _4224_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5328__A _6390_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4935__S0 _5051_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3790__B _3850_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5998__A _6032_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4068__A1 _6247_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6400__RESET_B fanout178/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4320_ _4767_/A _4320_/B vssd1 vssd1 vccd1 vccd1 _4321_/B sky130_fd_sc_hd__nand2_1
X_4251_ _3254_/A _5315_/B _4216_/A _4222_/B vssd1 vssd1 vccd1 vccd1 _4251_/X sky130_fd_sc_hd__a211o_1
XANTENNA__4288__S _4305_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3202_ _5480_/C _5322_/B vssd1 vssd1 vccd1 vccd1 _5292_/A sky130_fd_sc_hd__or2_1
XFILLER_0_38_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3205__B _4679_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4182_ _5217_/A _3761_/A _5219_/C _3758_/Y vssd1 vssd1 vccd1 vccd1 _4182_/X sky130_fd_sc_hd__a22o_1
X_3133_ _3193_/B _3237_/A _3126_/X vssd1 vssd1 vccd1 vccd1 _3133_/X sky130_fd_sc_hd__a21o_1
X_3064_ _6292_/Q vssd1 vssd1 vccd1 vccd1 _3064_/Y sky130_fd_sc_hd__inv_2
XANTENNA__5420__B _6420_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout146_A _4224_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4231__A1 _4224_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3966_ _3965_/X hold175/X _4206_/S vssd1 vssd1 vccd1 vccd1 _3966_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_18_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5705_ hold7/X _3805_/B _6060_/S vssd1 vssd1 vccd1 vccd1 hold8/A sky130_fd_sc_hd__mux2_1
XFILLER_0_92_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3897_ _3746_/X _3896_/X _3907_/A vssd1 vssd1 vccd1 vccd1 _3897_/X sky130_fd_sc_hd__o21a_1
X_5636_ _6195_/Q _4198_/B _4200_/S _6071_/Q _5675_/C1 vssd1 vssd1 vccd1 vccd1 _5638_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_33_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5567_ _3530_/D _5564_/X _5566_/Y _4637_/A vssd1 vssd1 vccd1 vccd1 _5568_/B sky130_fd_sc_hd__o2bb2a_1
XANTENNA__5731__A1 _5740_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold131 _5962_/X vssd1 vssd1 vccd1 vccd1 _6409_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold120 _6112_/Q vssd1 vssd1 vccd1 vccd1 hold120/X sky130_fd_sc_hd__dlygate4sd3_1
X_4518_ _4205_/X hold122/X _4518_/S vssd1 vssd1 vccd1 vccd1 _4518_/X sky130_fd_sc_hd__mux2_1
Xhold142 _4489_/X vssd1 vssd1 vccd1 vccd1 _6189_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5498_ _5478_/A _5478_/B _5490_/Y _5497_/X vssd1 vssd1 vccd1 vccd1 _5503_/A sky130_fd_sc_hd__a31o_1
Xhold153 _6213_/Q vssd1 vssd1 vccd1 vccd1 hold153/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold186 _4431_/X vssd1 vssd1 vccd1 vccd1 _6137_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold164 _4356_/X vssd1 vssd1 vccd1 vccd1 _6111_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4449_ _3923_/X hold203/X _4455_/S vssd1 vssd1 vccd1 vccd1 _4449_/X sky130_fd_sc_hd__mux2_1
Xhold175 _6070_/Q vssd1 vssd1 vccd1 vccd1 hold175/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4917__S0 _5052_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold197 _6074_/Q vssd1 vssd1 vccd1 vccd1 hold197/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_95_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6119_ _6399_/CLK _6119_/D fanout173/X vssd1 vssd1 vccd1 vccd1 _6119_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__4926__S _5060_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5798__A1 _6323_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout59_A _5815_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3785__B _3862_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3041__A _6297_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4213__A1 _5258_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3820_ _6164_/Q _3784_/X _3786_/X _6172_/Q vssd1 vssd1 vccd1 vccd1 _3820_/X sky130_fd_sc_hd__a22o_1
X_3751_ _3952_/A _4070_/A vssd1 vssd1 vccd1 vccd1 _3751_/X sky130_fd_sc_hd__or2_1
XFILLER_0_15_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3682_ _3682_/A _5991_/A _3680_/X vssd1 vssd1 vccd1 vccd1 _3682_/X sky130_fd_sc_hd__or3b_2
XFILLER_0_30_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5421_ _6437_/Q _4843_/X _5518_/S vssd1 vssd1 vccd1 vccd1 _5422_/C sky130_fd_sc_hd__mux2_1
X_5352_ _3484_/B _3482_/X _3484_/C _3365_/A vssd1 vssd1 vccd1 vccd1 _5353_/B sky130_fd_sc_hd__o31a_1
XFILLER_0_23_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4303_ _6064_/S _4299_/A _4302_/X vssd1 vssd1 vccd1 vccd1 _4303_/X sky130_fd_sc_hd__o21a_1
X_5283_ _5283_/A vssd1 vssd1 vccd1 vccd1 _5283_/Y sky130_fd_sc_hd__inv_2
X_4234_ _3656_/A _4229_/X _5343_/B _4233_/X vssd1 vssd1 vccd1 vccd1 _4234_/X sky130_fd_sc_hd__a211o_1
XANTENNA__3650__S input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4165_ _5217_/A _6343_/Q vssd1 vssd1 vccd1 vccd1 _4166_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_4_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3116_ _3116_/A _3285_/B _3116_/C vssd1 vssd1 vccd1 vccd1 _3116_/X sky130_fd_sc_hd__and3_1
X_4096_ _4096_/A vssd1 vssd1 vccd1 vccd1 _4098_/A sky130_fd_sc_hd__inv_2
X_3047_ _5981_/A vssd1 vssd1 vccd1 vccd1 _3047_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_77_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4204__A1 _5690_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4481__S _4482_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4998_ _6445_/Q _5056_/A2 _4997_/X vssd1 vssd1 vccd1 vccd1 _4998_/X sky130_fd_sc_hd__a21o_1
X_3949_ _6338_/Q _6342_/Q _6301_/Q vssd1 vssd1 vccd1 vccd1 _5216_/C sky130_fd_sc_hd__mux2_1
XFILLER_0_73_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5619_ _6380_/Q _5600_/X _5602_/X _6417_/Q _5618_/X vssd1 vssd1 vccd1 vccd1 _5620_/B
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4510__A _4510_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold642_A _6421_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout70 _4636_/B vssd1 vssd1 vccd1 vccd1 _4673_/B sky130_fd_sc_hd__buf_4
Xfanout92 _5029_/S vssd1 vssd1 vccd1 vccd1 _5371_/A sky130_fd_sc_hd__clkbuf_8
Xfanout81 _4321_/A vssd1 vssd1 vccd1 vccd1 _6057_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3036__A _5226_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5459__A0 _6422_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5970_ input6/X hold631/X _5975_/S vssd1 vssd1 vccd1 vccd1 _6418_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_35_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4921_ _6267_/Q _4758_/X _4920_/B _4757_/Y vssd1 vssd1 vccd1 vccd1 _4921_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_74_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4852_ _4852_/A _4852_/B _4852_/C vssd1 vssd1 vccd1 vccd1 _4852_/X sky130_fd_sc_hd__or3_1
XFILLER_0_74_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3803_ hold276/X _3715_/X _3794_/X _6214_/Q _3802_/X vssd1 vssd1 vccd1 vccd1 _3804_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_74_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4783_ _6320_/Q _4752_/X _4751_/B vssd1 vssd1 vccd1 vccd1 _4783_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_7_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3734_ _6301_/Q _5088_/B vssd1 vssd1 vccd1 vccd1 _3757_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_7_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3665_ _5158_/A _4346_/B vssd1 vssd1 vccd1 vccd1 _3666_/A sky130_fd_sc_hd__or2_1
XFILLER_0_70_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5404_ _6418_/Q _5403_/X _5471_/S vssd1 vssd1 vccd1 vccd1 _5404_/X sky130_fd_sc_hd__mux2_1
X_3596_ _4768_/A _3596_/B vssd1 vssd1 vccd1 vccd1 _3597_/A sky130_fd_sc_hd__and2_1
XANTENNA_fanout109_A _4732_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6384_ _6384_/CLK _6384_/D fanout167/X vssd1 vssd1 vccd1 vccd1 _6384_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_0_23_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5335_ _5725_/A _5332_/Y _5977_/S vssd1 vssd1 vccd1 vccd1 _5335_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__4370__B1 _5673_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5266_ _5266_/A _5266_/B _5266_/C _5266_/D vssd1 vssd1 vccd1 vccd1 _5266_/X sky130_fd_sc_hd__or4_1
XFILLER_0_55_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4217_ _5315_/B _5314_/A vssd1 vssd1 vccd1 vccd1 _4217_/X sky130_fd_sc_hd__or2_1
XANTENNA__4476__S _4482_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5197_ _6341_/Q _3502_/A _4188_/C _4079_/Y vssd1 vssd1 vccd1 vccd1 _5197_/X sky130_fd_sc_hd__a31o_1
XANTENNA__5161__A _6423_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3476__A2 _6425_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4148_ _4145_/X _4146_/X _4147_/X _4427_/S vssd1 vssd1 vccd1 vccd1 _4148_/X sky130_fd_sc_hd__a22o_2
X_4079_ _4079_/A vssd1 vssd1 vccd1 vccd1 _4079_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_93_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold592_A _6324_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4664__A1 _6341_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5071__A _5243_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5613__B1 _5676_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3927__B1 _3791_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3450_ hold69/X _3449_/X _3465_/A vssd1 vssd1 vccd1 vccd1 hold70/A sky130_fd_sc_hd__a21o_1
X_3381_ _4210_/A _6389_/Q vssd1 vssd1 vccd1 vccd1 _5480_/D sky130_fd_sc_hd__nand2_2
X_5120_ _5120_/A _5219_/C vssd1 vssd1 vccd1 vccd1 _5121_/B sky130_fd_sc_hd__xor2_1
XANTENNA__4104__B1 _3781_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5051_ _6115_/Q _6106_/Q _6098_/Q _6143_/Q _5051_/S0 _5052_/S1 vssd1 vssd1 vccd1
+ vccd1 _5051_/X sky130_fd_sc_hd__mux4_1
XANTENNA__4655__A1 _6343_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5852__A0 _6416_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4002_ _4111_/A _3930_/B _3935_/A vssd1 vssd1 vccd1 vccd1 _4003_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5953_ _3081_/Y _6396_/Q _5937_/B _5952_/A vssd1 vssd1 vccd1 vccd1 _5953_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_62_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5884_ _5878_/Y _5883_/X _5932_/S vssd1 vssd1 vccd1 vccd1 _5884_/X sky130_fd_sc_hd__mux2_1
X_4904_ _6323_/Q _6324_/Q _6325_/Q _6326_/Q vssd1 vssd1 vccd1 vccd1 _4905_/D sky130_fd_sc_hd__and4_1
X_4835_ _6322_/Q _4834_/X _5849_/S vssd1 vssd1 vccd1 vccd1 _4835_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_90_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4766_ _5272_/C vssd1 vssd1 vccd1 vccd1 _4766_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_7_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5855__S _5933_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3883__B _6337_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3717_ _4510_/A _4474_/A vssd1 vssd1 vccd1 vccd1 _4206_/S sky130_fd_sc_hd__or2_4
XFILLER_0_15_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4697_ hold416/X _3073_/A _4727_/S vssd1 vssd1 vccd1 vccd1 _4697_/X sky130_fd_sc_hd__mux2_1
X_3648_ _6121_/Q _6124_/Q input1/X vssd1 vssd1 vccd1 vccd1 _3648_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_3_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6436_ _6440_/CLK _6436_/D fanout171/X vssd1 vssd1 vccd1 vccd1 _6436_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_0_101_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3579_ _4734_/B _3579_/B vssd1 vssd1 vccd1 vccd1 _3580_/A sky130_fd_sc_hd__nand2_4
X_6367_ _6376_/CLK _6367_/D fanout166/X vssd1 vssd1 vccd1 vccd1 _6367_/Q sky130_fd_sc_hd__dfrtp_1
X_5318_ _3530_/D _5315_/X _5317_/X _5584_/A1 _5313_/X vssd1 vssd1 vccd1 vccd1 _5318_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_87_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6298_ _6343_/CLK _6298_/D fanout170/X vssd1 vssd1 vccd1 vccd1 _6298_/Q sky130_fd_sc_hd__dfstp_2
XANTENNA__5603__B _5603_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold13 hold13/A vssd1 vssd1 vccd1 vccd1 hold13/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 hold35/A vssd1 vssd1 vccd1 vccd1 hold35/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 hold46/A vssd1 vssd1 vccd1 vccd1 hold46/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 hold24/A vssd1 vssd1 vccd1 vccd1 hold24/X sky130_fd_sc_hd__dlygate4sd3_1
X_5249_ _5249_/A _5249_/B _5249_/C _5249_/D vssd1 vssd1 vccd1 vccd1 _5250_/C sky130_fd_sc_hd__or4_1
Xclkbuf_leaf_2_wb_clk_i clkbuf_leaf_6_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6410_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold57 hold57/A vssd1 vssd1 vccd1 vccd1 hold57/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold68 hold68/A vssd1 vssd1 vccd1 vccd1 hold68/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 hold79/A vssd1 vssd1 vccd1 vccd1 hold79/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6020__B1 _6057_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6425__RESET_B fanout173/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3845__C1 _3850_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xci2406_z80_203 vssd1 vssd1 vccd1 vccd1 ci2406_z80_203/HI io_oeb[32] sky130_fd_sc_hd__conb_1
XFILLER_0_76_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output22_A _6487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5062__A1 _6386_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5598__C1 _5691_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3612__A2 _5715_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4620_ _4744_/A _4615_/X _4617_/Y _4619_/X vssd1 vssd1 vccd1 vccd1 _4620_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_72_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_17_wb_clk_i_A _6404_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4551_ _4541_/A _4541_/C _4550_/C vssd1 vssd1 vccd1 vccd1 _4551_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_13_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3502_ _3502_/A _3725_/B vssd1 vssd1 vccd1 vccd1 _3537_/B sky130_fd_sc_hd__nor2_1
Xhold516 _6401_/Q vssd1 vssd1 vccd1 vccd1 _3645_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold527 _5559_/X vssd1 vssd1 vccd1 vccd1 _6334_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold505 _5830_/X vssd1 vssd1 vccd1 vccd1 _6377_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4482_ _4427_/X hold276/X _4482_/S vssd1 vssd1 vccd1 vccd1 _4482_/X sky130_fd_sc_hd__mux2_1
X_3433_ _5265_/A _3405_/Y _3406_/Y _3432_/X _4637_/A vssd1 vssd1 vccd1 vccd1 _3433_/X
+ sky130_fd_sc_hd__a221o_1
Xhold549 _6243_/Q vssd1 vssd1 vccd1 vccd1 hold549/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4325__A0 _5053_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold538 _6378_/Q vssd1 vssd1 vccd1 vccd1 hold538/X sky130_fd_sc_hd__dlygate4sd3_1
X_6221_ _6221_/CLK hold84/X vssd1 vssd1 vccd1 vccd1 hold83/A sky130_fd_sc_hd__dfxtp_1
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6152_ _6194_/CLK _6152_/D vssd1 vssd1 vccd1 vccd1 _6152_/Q sky130_fd_sc_hd__dfxtp_1
X_5103_ _6292_/Q _5083_/Y _5101_/X _5740_/A vssd1 vssd1 vccd1 vccd1 _5103_/X sky130_fd_sc_hd__o22a_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3364_ _6317_/Q _6316_/Q vssd1 vssd1 vccd1 vccd1 _4762_/S sky130_fd_sc_hd__or2_1
XFILLER_0_0_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4628__A1 _3952_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3295_ _5270_/A _3339_/A _5360_/B _3295_/D vssd1 vssd1 vccd1 vccd1 _3318_/D sky130_fd_sc_hd__and4b_1
XANTENNA__3224__A _3369_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6083_ _6271_/CLK _6083_/D fanout169/X vssd1 vssd1 vccd1 vccd1 _6083_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5034_ _5054_/A _6057_/C vssd1 vssd1 vccd1 vccd1 _5034_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_79_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3138__D_N _3183_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout176_A fanout177/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5936_ _5949_/C _5936_/B vssd1 vssd1 vccd1 vccd1 _5936_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__4800__A1 _5054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5867_ _5847_/X _5858_/A _5866_/X vssd1 vssd1 vccd1 vccd1 _5869_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_16_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5798_ _6323_/Q _5825_/S _5850_/B1 _5797_/X vssd1 vssd1 vccd1 vccd1 _5798_/X sky130_fd_sc_hd__a22o_1
X_4818_ _5773_/A _4818_/B vssd1 vssd1 vccd1 vccd1 _4818_/Y sky130_fd_sc_hd__nand2_1
X_4749_ _5077_/A _3597_/A _3771_/Y _4748_/X _4746_/Y vssd1 vssd1 vccd1 vccd1 _5772_/S
+ sky130_fd_sc_hd__a41o_2
XFILLER_0_71_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5761__C1 _5747_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3118__B _3183_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6419_ _6423_/CLK _6419_/D fanout175/X vssd1 vssd1 vccd1 vccd1 _6419_/Q sky130_fd_sc_hd__dfrtp_4
Xoutput25 _6280_/Q vssd1 vssd1 vccd1 vccd1 io_out[11] sky130_fd_sc_hd__buf_12
XFILLER_0_101_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput47 _3650_/X vssd1 vssd1 vccd1 vccd1 io_out[33] sky130_fd_sc_hd__buf_12
Xoutput36 _6290_/Q vssd1 vssd1 vccd1 vccd1 io_out[21] sky130_fd_sc_hd__buf_12
XANTENNA__3833__S _3838_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4411__S0 _5676_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4664__S _4674_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5831__A3 _3580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5044__A1 _6385_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3044__A _5553_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3080_ _3080_/A vssd1 vssd1 vccd1 vccd1 _3080_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3979__A _6243_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5035__A1 _6273_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3982_ _6292_/Q _4073_/C _3978_/Y _3981_/Y vssd1 vssd1 vccd1 vccd1 _5123_/B sky130_fd_sc_hd__a31o_1
XFILLER_0_57_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5721_ _6272_/Q hold534/X _5723_/S vssd1 vssd1 vccd1 vccd1 _5721_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_72_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5652_ _5651_/X _5648_/X _4053_/X _4404_/X _5691_/S _5690_/S vssd1 vssd1 vccd1 vccd1
+ _5652_/X sky130_fd_sc_hd__mux4_1
X_5583_ _5096_/A _5291_/A _5580_/X _5582_/X vssd1 vssd1 vccd1 vccd1 _5583_/X sky130_fd_sc_hd__a211o_1
X_4603_ _5695_/A1 hold532/X _4546_/Y _4602_/X vssd1 vssd1 vccd1 vccd1 _4603_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4546__B1 _5339_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3219__A _4228_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4534_ hold464/X _6293_/Q _4539_/S vssd1 vssd1 vccd1 vccd1 _4534_/X sky130_fd_sc_hd__mux2_1
Xhold302 _6407_/Q vssd1 vssd1 vccd1 vccd1 hold302/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold335 _4672_/X vssd1 vssd1 vccd1 vccd1 _6265_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold313 _4647_/X vssd1 vssd1 vccd1 vccd1 _6260_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold324 _4303_/X vssd1 vssd1 vccd1 vccd1 _6081_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold368 _4610_/X vssd1 vssd1 vccd1 vccd1 _6250_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold357 _6299_/Q vssd1 vssd1 vccd1 vccd1 hold357/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_7_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4465_ _4465_/A _5959_/B vssd1 vssd1 vccd1 vccd1 _4473_/S sky130_fd_sc_hd__or2_4
Xhold346 _6282_/Q vssd1 vssd1 vccd1 vccd1 hold346/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5434__A _5715_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6204_ _6204_/CLK _6204_/D fanout174/X vssd1 vssd1 vccd1 vccd1 _6204_/Q sky130_fd_sc_hd__dfrtp_1
X_3416_ _3396_/Y _3401_/A _3415_/X _5935_/A vssd1 vssd1 vccd1 vccd1 _3439_/S sky130_fd_sc_hd__a31o_1
X_4396_ _4424_/A _4396_/B vssd1 vssd1 vccd1 vccd1 _4396_/Y sky130_fd_sc_hd__nor2_1
Xhold379 _6373_/Q vssd1 vssd1 vccd1 vccd1 _5765_/A sky130_fd_sc_hd__dlygate4sd3_1
X_3347_ _5574_/A _3336_/A _3336_/B _3336_/C _3309_/Y vssd1 vssd1 vccd1 vccd1 _3657_/B
+ sky130_fd_sc_hd__o41a_2
X_6135_ _6410_/CLK _6135_/D vssd1 vssd1 vccd1 vccd1 _6135_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3278_ _3278_/A _5303_/A vssd1 vssd1 vccd1 vccd1 _5322_/D sky130_fd_sc_hd__nor2_4
XFILLER_0_84_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4484__S _4491_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5017_ _6272_/Q _4758_/X _5016_/B _4757_/Y vssd1 vssd1 vccd1 vccd1 _5017_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5468__A2_N _5377_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5919_ _6333_/Q _5928_/A2 _5928_/B1 _5918_/X vssd1 vssd1 vccd1 vccd1 _5919_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4880__S0 _5358_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6088__RESET_B fanout174/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4659__S _4674_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4935__S1 _5052_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3790__C _3838_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4068__A2 _6248_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3815__A2 _3789_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5017__A1 _6272_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4776__B1 _4867_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4250_ _4214_/A _5291_/A _5324_/C _3337_/A _4249_/X vssd1 vssd1 vccd1 vccd1 _4273_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_10_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3503__B2 _6118_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3201_ _3278_/A _3628_/B vssd1 vssd1 vccd1 vccd1 _5322_/B sky130_fd_sc_hd__nor2_1
X_4181_ _6292_/Q _4172_/X _4173_/Y _4180_/X vssd1 vssd1 vccd1 vccd1 _5219_/C sky130_fd_sc_hd__o31a_1
X_3132_ _4214_/B _3132_/B vssd1 vssd1 vccd1 vccd1 _3237_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_38_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3063_ _3063_/A vssd1 vssd1 vccd1 vccd1 _3063_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3806__A2 _3784_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3502__A _3502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3221__B _3566_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3648__S input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3965_ _3963_/X _3964_/X _4427_/S vssd1 vssd1 vccd1 vccd1 _3965_/X sky130_fd_sc_hd__mux2_2
X_3896_ _3748_/Y _4188_/C _3896_/S vssd1 vssd1 vccd1 vccd1 _3896_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_70_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5704_ hold3/X _3811_/Y _6060_/S vssd1 vssd1 vccd1 vccd1 hold4/A sky130_fd_sc_hd__mux2_1
XANTENNA_fanout139_A _6256_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5635_ _5635_/A _5635_/B vssd1 vssd1 vccd1 vccd1 _5635_/X sky130_fd_sc_hd__or2_1
XFILLER_0_85_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5566_ _4541_/C _4258_/X _5565_/X vssd1 vssd1 vccd1 vccd1 _5566_/Y sky130_fd_sc_hd__a21oi_1
Xhold110 _4355_/X vssd1 vssd1 vccd1 vccd1 _6110_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5731__A2 _5729_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold143 _6104_/Q vssd1 vssd1 vccd1 vccd1 hold143/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold121 _4357_/X vssd1 vssd1 vccd1 vccd1 _6112_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4517_ _4148_/X hold83/X _4518_/S vssd1 vssd1 vccd1 vccd1 hold84/A sky130_fd_sc_hd__mux2_1
XANTENNA__4479__S _4482_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5497_ _5476_/B _5489_/B _5554_/A vssd1 vssd1 vccd1 vccd1 _5497_/X sky130_fd_sc_hd__o21a_1
Xhold132 _6134_/Q vssd1 vssd1 vccd1 vccd1 hold132/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold176 _3966_/X vssd1 vssd1 vccd1 vccd1 _6070_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4448_ _3881_/X hold233/X _4455_/S vssd1 vssd1 vccd1 vccd1 _4448_/X sky130_fd_sc_hd__mux2_1
Xhold165 _6143_/Q vssd1 vssd1 vccd1 vccd1 hold165/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold154 _4508_/X vssd1 vssd1 vccd1 vccd1 _6213_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold187 _6128_/Q vssd1 vssd1 vccd1 vccd1 hold187/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold198 _6142_/Q vssd1 vssd1 vccd1 vccd1 hold198/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4917__S1 _5051_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5495__A1 _6417_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4379_ _3080_/Y _3700_/B _4382_/C vssd1 vssd1 vccd1 vccd1 _4379_/Y sky130_fd_sc_hd__a21oi_1
X_6118_ _6399_/CLK _6118_/D fanout173/X vssd1 vssd1 vccd1 vccd1 _6118_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6049_ _3046_/A _6047_/X _6048_/Y hold399/X _6029_/Y vssd1 vssd1 vccd1 vccd1 _6049_/X
+ sky130_fd_sc_hd__o32a_1
XANTENNA__4942__S _5058_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold420_A _6246_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold518_A _6385_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5339__A _5339_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3785__C _3838_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5486__A1 _5553_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5238__A1 _6298_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3750_ _6303_/Q _3757_/B _6304_/Q vssd1 vssd1 vccd1 vccd1 _3985_/A sky130_fd_sc_hd__and3b_4
XFILLER_0_82_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3681_ _3611_/A _5739_/A _3611_/Y vssd1 vssd1 vccd1 vccd1 _3682_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5420_ _5715_/A _6420_/Q vssd1 vssd1 vccd1 vccd1 _5422_/B sky130_fd_sc_hd__or2_1
XFILLER_0_42_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5351_ hold433/X _5603_/B _5727_/S vssd1 vssd1 vccd1 vccd1 _5351_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_10_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4921__B1 _4920_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5282_ _5077_/A _5279_/X _5281_/X vssd1 vssd1 vccd1 vccd1 _5283_/A sky130_fd_sc_hd__a21oi_1
X_4302_ _6270_/Q _4316_/B _4297_/X _4301_/X vssd1 vssd1 vccd1 vccd1 _4302_/X sky130_fd_sc_hd__a22o_1
X_4233_ _3132_/B _5733_/A _3770_/A _4232_/X vssd1 vssd1 vccd1 vccd1 _4233_/X sky130_fd_sc_hd__a31o_1
X_4164_ _5217_/A _6343_/Q vssd1 vssd1 vccd1 vccd1 _4164_/X sky130_fd_sc_hd__or2_1
X_3115_ _3289_/A _6254_/Q _3534_/A vssd1 vssd1 vccd1 vccd1 _3116_/C sky130_fd_sc_hd__or3_2
XFILLER_0_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4328__A _4510_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4095_ _4394_/A _4095_/B vssd1 vssd1 vccd1 vccd1 _4096_/A sky130_fd_sc_hd__xnor2_1
X_3046_ _3046_/A vssd1 vssd1 vccd1 vccd1 _3046_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_77_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3660__B1 _3309_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5159__A _6421_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5401__B2 _5441_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4997_ _6271_/Q _4758_/X _4996_/B _4757_/Y vssd1 vssd1 vccd1 vccd1 _4997_/X sky130_fd_sc_hd__a22o_1
X_3948_ _3948_/A _3948_/B vssd1 vssd1 vccd1 vccd1 _5209_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_73_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3879_ _3724_/A _5250_/A _3768_/Y vssd1 vssd1 vccd1 vccd1 _3879_/X sky130_fd_sc_hd__a21o_1
X_5618_ _6292_/Q _5587_/X _5594_/Y _5617_/X vssd1 vssd1 vccd1 vccd1 _5618_/X sky130_fd_sc_hd__a22o_1
X_5549_ _6057_/A _5547_/X _5548_/Y _5558_/S vssd1 vssd1 vccd1 vccd1 _5549_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_14_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3407__A _6389_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5468__B2 _5377_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4937__S _5053_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout71_A _3721_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5640__A1 _6294_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3651__B1 _4541_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5640__B2 _6419_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout71 _3721_/Y vssd1 vssd1 vccd1 vccd1 _5675_/C1 sky130_fd_sc_hd__clkbuf_8
Xfanout60 _5850_/B1 vssd1 vssd1 vccd1 vccd1 _5928_/B1 sky130_fd_sc_hd__buf_4
Xfanout82 _3687_/Y vssd1 vssd1 vccd1 vccd1 _4425_/A2 sky130_fd_sc_hd__buf_4
XFILLER_0_91_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout93 _3476_/Y vssd1 vssd1 vccd1 vccd1 _5029_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_0_101_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4903__B1 _6326_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_26_wb_clk_i _6404_/CLK vssd1 vssd1 vccd1 vccd1 _6297_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_99_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4920_ _5054_/A _4920_/B vssd1 vssd1 vccd1 vccd1 _4920_/Y sky130_fd_sc_hd__nand2_1
X_4851_ _6420_/Q _4758_/X _4849_/X _5061_/A1 vssd1 vssd1 vccd1 vccd1 _4852_/C sky130_fd_sc_hd__a22o_1
XFILLER_0_74_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3802_ _6135_/Q _3789_/X _3791_/X _6414_/Q vssd1 vssd1 vccd1 vccd1 _3802_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_27_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4782_ hold330/X _4781_/X _5068_/S vssd1 vssd1 vccd1 vccd1 _4782_/X sky130_fd_sc_hd__mux2_1
X_3733_ _6303_/Q _4070_/A vssd1 vssd1 vccd1 vccd1 _3736_/S sky130_fd_sc_hd__and2b_1
XFILLER_0_70_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3664_ _3164_/Y _3431_/A _3553_/Y vssd1 vssd1 vccd1 vccd1 _3668_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5403_ _5401_/X _5402_/X _5560_/D vssd1 vssd1 vccd1 vccd1 _5403_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_30_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3173__A2 _3502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3595_ _4772_/A _5481_/C _4767_/C _3595_/D vssd1 vssd1 vccd1 vccd1 _3596_/B sky130_fd_sc_hd__and4bb_1
X_6383_ _6383_/CLK _6383_/D fanout168/X vssd1 vssd1 vccd1 vccd1 _6383_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_0_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5334_ _5989_/A _5333_/X _5727_/S vssd1 vssd1 vccd1 vccd1 _6307_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_11_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5265_ _5265_/A _5265_/B vssd1 vssd1 vccd1 vccd1 _5266_/D sky130_fd_sc_hd__nor2_1
X_4216_ _4216_/A _4216_/B vssd1 vssd1 vccd1 vccd1 _5314_/A sky130_fd_sc_hd__or2_1
X_5196_ _6341_/Q _5206_/B _5196_/S vssd1 vssd1 vccd1 vccd1 _5196_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5161__B _6422_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3476__A3 _3473_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5870__A1 _6381_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4147_ hold140/X hold79/X hold83/X hold99/X _5676_/C1 _5676_/B1 vssd1 vssd1 vccd1
+ vccd1 _4147_/X sky130_fd_sc_hd__mux4_1
XANTENNA__4058__A _6247_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4078_ _3758_/Y _5219_/B _3761_/Y _4075_/A vssd1 vssd1 vccd1 vccd1 _4079_/A sky130_fd_sc_hd__o2bb2a_1
XANTENNA__5622__A1 _6418_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4521__A _5447_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3380_ _4214_/A _5574_/A vssd1 vssd1 vccd1 vccd1 _4734_/B sky130_fd_sc_hd__nor2_8
X_5050_ hold409/X _5049_/X _5068_/S vssd1 vssd1 vccd1 vccd1 _5050_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_46_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4001_ _4111_/A _4001_/B vssd1 vssd1 vccd1 vccd1 _4009_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5952_ _5952_/A _5952_/B vssd1 vssd1 vccd1 vccd1 _5952_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_87_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_46_wb_clk_i_A clkbuf_leaf_6_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_4903_ _6324_/Q _6325_/Q _4866_/B _6326_/Q vssd1 vssd1 vccd1 vccd1 _4903_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_75_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5883_ _5882_/X _5876_/A _5931_/S vssd1 vssd1 vccd1 vccd1 _5883_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_7_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4834_ _6374_/Q _4796_/B _4832_/X _4833_/X vssd1 vssd1 vccd1 vccd1 _4834_/X sky130_fd_sc_hd__o22a_1
X_4765_ _4765_/A _5481_/C vssd1 vssd1 vccd1 vccd1 _5272_/C sky130_fd_sc_hd__or2_1
XFILLER_0_55_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout121_A _5560_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3716_ _3850_/A _3850_/B _3861_/S vssd1 vssd1 vccd1 vccd1 _4474_/A sky130_fd_sc_hd__or3_1
XFILLER_0_70_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4696_ hold653/X _4695_/X _5447_/S vssd1 vssd1 vccd1 vccd1 _4696_/X sky130_fd_sc_hd__mux2_1
X_3647_ _6120_/Q _6125_/Q input1/X vssd1 vssd1 vccd1 vccd1 _3647_/X sky130_fd_sc_hd__mux2_2
X_6435_ _6440_/CLK _6435_/D fanout171/X vssd1 vssd1 vccd1 vccd1 _6435_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_0_3_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3578_ _4541_/B _3426_/A _3386_/B vssd1 vssd1 vccd1 vccd1 _3579_/B sky130_fd_sc_hd__a21o_2
X_6366_ _6376_/CLK _6366_/D fanout166/X vssd1 vssd1 vccd1 vccd1 _6366_/Q sky130_fd_sc_hd__dfrtp_1
X_5317_ _5317_/A _5317_/B _5316_/X vssd1 vssd1 vccd1 vccd1 _5317_/X sky130_fd_sc_hd__or3b_1
XFILLER_0_11_362 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4487__S _4491_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6297_ _6297_/CLK _6297_/D fanout176/X vssd1 vssd1 vccd1 vccd1 _6297_/Q sky130_fd_sc_hd__dfstp_4
Xhold14 hold14/A vssd1 vssd1 vccd1 vccd1 hold14/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 hold47/A vssd1 vssd1 vccd1 vccd1 hold47/X sky130_fd_sc_hd__dlygate4sd3_1
X_5248_ _5249_/D _5247_/X _5560_/B vssd1 vssd1 vccd1 vccd1 _5255_/S sky130_fd_sc_hd__a21oi_1
Xhold36 hold36/A vssd1 vssd1 vccd1 vccd1 hold36/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 hold25/A vssd1 vssd1 vccd1 vccd1 hold25/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5322__D _5322_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold69 hold69/A vssd1 vssd1 vccd1 vccd1 hold69/X sky130_fd_sc_hd__dlygate4sd3_1
X_5179_ _3990_/X _5178_/A _5173_/X _5178_/Y vssd1 vssd1 vccd1 vccd1 _5179_/X sky130_fd_sc_hd__a22o_1
Xhold58 hold58/A vssd1 vssd1 vccd1 vccd1 hold58/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold500_A _6247_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6020__B2 _4882_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5347__A _5347_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xci2406_z80_204 vssd1 vssd1 vccd1 vccd1 ci2406_z80_204/HI io_oeb[33] sky130_fd_sc_hd__conb_1
XFILLER_0_8_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4573__A1 _5695_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4550_ _5578_/A _4550_/B _4550_/C vssd1 vssd1 vccd1 vccd1 _4550_/Y sky130_fd_sc_hd__nor3_1
Xhold517 _3646_/X vssd1 vssd1 vccd1 vccd1 _6398_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3501_ _4637_/A _3501_/B vssd1 vssd1 vccd1 vccd1 _3501_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_12_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold506 _6078_/Q vssd1 vssd1 vccd1 vccd1 _4287_/A sky130_fd_sc_hd__buf_1
X_4481_ _4420_/X hold193/X _4482_/S vssd1 vssd1 vccd1 vccd1 _4481_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5691__S _5691_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3432_ _5265_/A _3224_/X _4734_/B _3431_/Y _3308_/X vssd1 vssd1 vccd1 vccd1 _3432_/X
+ sky130_fd_sc_hd__o311a_1
Xhold528 _6234_/Q vssd1 vssd1 vccd1 vccd1 hold528/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold539 _5844_/X vssd1 vssd1 vccd1 vccd1 _6378_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6220_ _6444_/CLK _6220_/D vssd1 vssd1 vccd1 vccd1 _6220_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3363_ _3363_/A _3363_/B vssd1 vssd1 vccd1 vccd1 _3365_/B sky130_fd_sc_hd__nor2_4
XFILLER_0_0_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_41_wb_clk_i clkbuf_leaf_6_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6448_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_6151_ _6414_/CLK hold66/X vssd1 vssd1 vccd1 vccd1 hold65/A sky130_fd_sc_hd__dfxtp_1
X_5102_ _5102_/A _5102_/B vssd1 vssd1 vccd1 vccd1 _5102_/Y sky130_fd_sc_hd__nor2_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4628__A2 _4615_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3294_ _4255_/B _3654_/A _4747_/D vssd1 vssd1 vccd1 vccd1 _3295_/D sky130_fd_sc_hd__a21o_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4089__B1 _3781_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5825__A1 _6325_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6082_ _6376_/CLK _6082_/D fanout169/X vssd1 vssd1 vccd1 vccd1 _6082_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__3224__B _3566_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5033_ _5032_/X _5031_/X _5053_/S vssd1 vssd1 vccd1 vccd1 _6057_/C sky130_fd_sc_hd__mux2_2
XANTENNA_clkbuf_leaf_2_wb_clk_i_A clkbuf_leaf_6_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_73_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout169_A fanout181/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5935_ _5935_/A _5937_/B vssd1 vssd1 vccd1 vccd1 _5949_/B sky130_fd_sc_hd__and2_1
X_5866_ _6379_/Q _6380_/Q _5926_/A vssd1 vssd1 vccd1 vccd1 _5866_/X sky130_fd_sc_hd__o21a_1
XANTENNA__4800__A2 _4788_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4817_ _4816_/X _6321_/Q _5825_/S vssd1 vssd1 vccd1 vccd1 _4818_/B sky130_fd_sc_hd__mux2_1
XANTENNA__4013__B1 _3781_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5797_ _6323_/Q _6375_/Q _5849_/S vssd1 vssd1 vccd1 vccd1 _5797_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4071__A _6246_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4748_ _3600_/C _3386_/B _4748_/C _4748_/D vssd1 vssd1 vccd1 vccd1 _4748_/X sky130_fd_sc_hd__and4bb_1
XFILLER_0_7_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4679_ _4679_/A _5560_/A _4679_/C _4679_/D vssd1 vssd1 vccd1 vccd1 _5192_/S sky130_fd_sc_hd__or4_4
XFILLER_0_71_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6418_ _6423_/CLK _6418_/D fanout175/X vssd1 vssd1 vccd1 vccd1 _6418_/Q sky130_fd_sc_hd__dfrtp_4
Xoutput15 _6481_/X vssd1 vssd1 vccd1 vccd1 io_oeb[22] sky130_fd_sc_hd__buf_12
XFILLER_0_31_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput48 _3649_/X vssd1 vssd1 vccd1 vccd1 io_out[34] sky130_fd_sc_hd__buf_12
Xoutput37 _6263_/Q vssd1 vssd1 vccd1 vccd1 io_out[22] sky130_fd_sc_hd__buf_12
XANTENNA__4411__S1 _5676_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput26 _6281_/Q vssd1 vssd1 vccd1 vccd1 io_out[12] sky130_fd_sc_hd__buf_12
XANTENNA__5106__S _5447_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3415__A _4637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6349_ _6355_/CLK hold6/X vssd1 vssd1 vccd1 vccd1 hold5/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__3827__B1 _3786_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3922__S0 _5676_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5077__A _5077_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4858__A2 _4313_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3279__D1 _5322_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3979__B _6244_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3294__A1 _4255_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3060__A _6248_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3981_ _3981_/A _3981_/B vssd1 vssd1 vccd1 vccd1 _3981_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_69_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5720_ _6271_/Q hold502/X _5723_/S vssd1 vssd1 vccd1 vccd1 _5720_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_57_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4794__B2 _4788_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5651_ _5651_/A _5651_/B vssd1 vssd1 vccd1 vccd1 _5651_/X sky130_fd_sc_hd__or2_1
X_5582_ _5480_/D _5577_/X _5581_/X _3337_/A vssd1 vssd1 vccd1 vccd1 _5582_/X sky130_fd_sc_hd__a2bb2o_1
XANTENNA__5743__B1 _5735_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4602_ hold414/X _4567_/Y _4568_/X _6447_/Q _4601_/X vssd1 vssd1 vccd1 vccd1 _4602_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3219__B _3566_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4533_ hold528/X _6292_/Q _4539_/S vssd1 vssd1 vccd1 vccd1 _4533_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_80_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold325 _6391_/Q vssd1 vssd1 vccd1 vccd1 _3466_/B sky130_fd_sc_hd__buf_1
XANTENNA__5715__A _5715_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold314 _6310_/Q vssd1 vssd1 vccd1 vccd1 _3070_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold303 _5960_/X vssd1 vssd1 vccd1 vccd1 _6407_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6203_ _6397_/CLK hold32/X fanout174/X vssd1 vssd1 vccd1 vccd1 hold31/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold358 _5255_/X vssd1 vssd1 vccd1 vccd1 _6299_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold336 _6335_/Q vssd1 vssd1 vccd1 vccd1 _5561_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold369 _6083_/Q vssd1 vssd1 vccd1 vccd1 _4313_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_0_7_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5434__B _6421_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold347 _4916_/X vssd1 vssd1 vccd1 vccd1 _6282_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4464_ _4427_/X hold283/X _4464_/S vssd1 vssd1 vccd1 vccd1 _6167_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_68_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3415_ _4637_/A _3415_/B vssd1 vssd1 vccd1 vccd1 _3415_/X sky130_fd_sc_hd__or2_1
XFILLER_0_0_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4395_ _4395_/A _4395_/B vssd1 vssd1 vccd1 vccd1 _4396_/B sky130_fd_sc_hd__xnor2_1
X_3346_ _4558_/A _3581_/A _3343_/Y _5481_/A _3345_/X vssd1 vssd1 vccd1 vccd1 _3346_/Y
+ sky130_fd_sc_hd__a311oi_1
X_6134_ _6413_/CLK _6134_/D vssd1 vssd1 vccd1 vccd1 _6134_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6316__RESET_B fanout173/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3277_ _3277_/A _3520_/A vssd1 vssd1 vccd1 vccd1 _3386_/B sky130_fd_sc_hd__or2_2
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5016_ _5054_/A _5016_/B vssd1 vssd1 vccd1 vccd1 _5016_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3809__B1 _3794_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5918_ _6366_/Q _6385_/Q _5927_/S vssd1 vssd1 vccd1 vccd1 _5918_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_75_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5329__A3 _4734_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5849_ _6360_/Q _6379_/Q _5849_/S vssd1 vssd1 vccd1 vccd1 _5849_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4880__S1 _4326_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4537__A1 _6296_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3129__B _3656_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5973__A0 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4776__A1 _5061_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5513__A2_N _5377_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4528__A1 _6271_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3055__A _6244_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4180_ _4172_/C _4178_/Y _4179_/X _4178_/A _3064_/Y vssd1 vssd1 vccd1 vccd1 _4180_/X
+ sky130_fd_sc_hd__a221o_1
X_3200_ _3483_/A _4318_/B vssd1 vssd1 vccd1 vccd1 _5480_/C sky130_fd_sc_hd__or2_1
X_3131_ _3290_/B _3374_/A vssd1 vssd1 vccd1 vccd1 _3683_/C sky130_fd_sc_hd__nor2_4
X_3062_ _3062_/A vssd1 vssd1 vccd1 vccd1 _4029_/B sky130_fd_sc_hd__inv_2
XANTENNA__3502__B _3725_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5639__S0 _5691_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3964_ hold183/X hold63/X hold288/X hold109/X _5676_/C1 _4200_/S vssd1 vssd1 vccd1
+ vccd1 _3964_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_18_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3895_ _3761_/A _5216_/B _5130_/B _3985_/A vssd1 vssd1 vccd1 vccd1 _3895_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_45_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5703_ hold5/X _3818_/Y _6060_/S vssd1 vssd1 vccd1 vccd1 hold6/A sky130_fd_sc_hd__mux2_1
XFILLER_0_70_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5716__A0 _6267_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5634_ _6131_/Q _4382_/B _4384_/S _6210_/Q _5673_/C1 vssd1 vssd1 vccd1 vccd1 _5635_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_33_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5192__A1 _6296_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5565_ _3656_/A _3100_/B _4257_/Y _3226_/Y _5578_/A vssd1 vssd1 vccd1 vccd1 _5565_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_79_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold100 _4359_/X vssd1 vssd1 vccd1 vccd1 _6114_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold111 _6162_/Q vssd1 vssd1 vccd1 vccd1 hold111/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold144 _4343_/X vssd1 vssd1 vccd1 vccd1 _6104_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4516_ _4102_/X hold103/X _4518_/S vssd1 vssd1 vccd1 vccd1 _4516_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_13_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold122 _6222_/Q vssd1 vssd1 vccd1 vccd1 hold122/X sky130_fd_sc_hd__dlygate4sd3_1
X_5496_ hold383/X _5495_/X _6060_/S vssd1 vssd1 vccd1 vccd1 _5496_/X sky130_fd_sc_hd__mux2_1
Xhold133 _4421_/X vssd1 vssd1 vccd1 vccd1 _6134_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold155 _6178_/Q vssd1 vssd1 vccd1 vccd1 hold155/X sky130_fd_sc_hd__dlygate4sd3_1
X_4447_ _4510_/A _4465_/A vssd1 vssd1 vccd1 vccd1 _4455_/S sky130_fd_sc_hd__or2_4
Xhold166 _4437_/X vssd1 vssd1 vccd1 vccd1 _6143_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold177 _6211_/Q vssd1 vssd1 vccd1 vccd1 hold177/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold188 _4368_/X vssd1 vssd1 vccd1 vccd1 _6128_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold199 _6092_/Q vssd1 vssd1 vccd1 vccd1 hold199/X sky130_fd_sc_hd__dlygate4sd3_1
X_6117_ _6399_/CLK _6117_/D fanout173/X vssd1 vssd1 vccd1 vccd1 _6117_/Q sky130_fd_sc_hd__dfrtp_1
X_4378_ _4376_/Y _4377_/X _3910_/Y vssd1 vssd1 vccd1 vccd1 _4378_/X sky130_fd_sc_hd__a21o_1
XANTENNA__4495__S _4500_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3329_ _6293_/Q _4081_/S _3328_/Y _3323_/X _3324_/Y vssd1 vssd1 vccd1 vccd1 _3336_/A
+ sky130_fd_sc_hd__a2111o_1
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6048_ _6048_/A _6063_/S vssd1 vssd1 vccd1 vccd1 _6048_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_95_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6448__SET_B fanout181/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3839__S _3862_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5339__B _5977_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3497__A1 _4070_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4997__A1 _6271_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4749__A1 _5077_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3680_ _5096_/B _3675_/X _3679_/X vssd1 vssd1 vccd1 vccd1 _3680_/X sky130_fd_sc_hd__o21a_1
X_5350_ _4382_/B _5349_/Y _5727_/S vssd1 vssd1 vccd1 vccd1 _5350_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4921__A1 _6267_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5281_ _3656_/A _6118_/Q _5277_/Y _5280_/X _5584_/A1 vssd1 vssd1 vccd1 vccd1 _5281_/X
+ sky130_fd_sc_hd__a32o_1
X_4301_ _4305_/S _4304_/B _5695_/A1 vssd1 vssd1 vccd1 vccd1 _4301_/X sky130_fd_sc_hd__a21o_1
X_4232_ _3656_/A _4541_/A _3952_/B _3109_/B _5315_/A vssd1 vssd1 vccd1 vccd1 _4232_/X
+ sky130_fd_sc_hd__a41o_1
X_4163_ _4163_/A _5107_/B vssd1 vssd1 vccd1 vccd1 _4163_/Y sky130_fd_sc_hd__nand2_1
X_3114_ _4744_/B _6254_/Q vssd1 vssd1 vccd1 vccd1 _3233_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_65_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4094_ _4095_/B vssd1 vssd1 vccd1 vccd1 _4094_/Y sky130_fd_sc_hd__inv_2
X_3045_ _6425_/Q vssd1 vssd1 vccd1 vccd1 _5097_/A sky130_fd_sc_hd__inv_2
XANTENNA__5634__C1 _5673_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout151_A _3566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4996_ _5054_/A _4996_/B vssd1 vssd1 vccd1 vccd1 _4996_/Y sky130_fd_sc_hd__nand2_1
X_3947_ _6243_/Q _6244_/Q vssd1 vssd1 vccd1 vccd1 _3948_/B sky130_fd_sc_hd__xor2_1
XANTENNA__5159__B _6420_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5401__A2 _5377_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3878_ _3878_/A _3878_/B vssd1 vssd1 vccd1 vccd1 _5250_/A sky130_fd_sc_hd__nor2_1
X_5617_ _5616_/X _4375_/X _5691_/S vssd1 vssd1 vccd1 vccd1 _5617_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_45_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5548_ _5548_/A _6057_/A vssd1 vssd1 vccd1 vccd1 _5548_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__4912__A1 _6326_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4373__C1 _5675_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6331__RESET_B fanout171/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5479_ _4313_/C _5377_/X hold522/X vssd1 vssd1 vccd1 vccd1 _5479_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_1_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4953__S _5557_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5625__C1 _5676_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3651__A1 _5715_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold628_A _6392_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout83 _3687_/Y vssd1 vssd1 vccd1 vccd1 _4391_/A2 sky130_fd_sc_hd__clkbuf_4
Xfanout72 _5673_/C1 vssd1 vssd1 vccd1 vccd1 _5676_/C1 sky130_fd_sc_hd__buf_6
XANTENNA__5784__S _5784_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout61 _4751_/Y vssd1 vssd1 vccd1 vccd1 _5850_/B1 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_91_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout94 _4313_/C vssd1 vssd1 vccd1 vccd1 _6057_/A sky130_fd_sc_hd__buf_4
XFILLER_0_36_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4903__A1 _6324_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4429__A _4510_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output45_A _3648_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_36_wb_clk_i_A clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__4164__A _5217_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4850_ _6437_/Q _4756_/Y _4757_/Y _4843_/X _4754_/X vssd1 vssd1 vccd1 vccd1 _4852_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3801_ hold283/X _3784_/X _3786_/X hold241/X vssd1 vssd1 vccd1 vccd1 _3804_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_7_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4781_ _6078_/Q _5557_/S _4780_/X vssd1 vssd1 vccd1 vccd1 _4781_/X sky130_fd_sc_hd__o21a_1
X_3732_ _6242_/Q _3732_/B vssd1 vssd1 vccd1 vccd1 _3738_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5147__A1 _6343_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3663_ _3656_/X _3661_/X _3662_/X _3655_/Y vssd1 vssd1 vccd1 vccd1 _3663_/X sky130_fd_sc_hd__o31a_1
XFILLER_0_70_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5402_ hold585/X input6/X _5469_/S vssd1 vssd1 vccd1 vccd1 _5402_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_2_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6382_ _6383_/CLK _6382_/D fanout168/X vssd1 vssd1 vccd1 vccd1 _6382_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_11_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3227__B _3566_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3594_ _3594_/A _5733_/A vssd1 vssd1 vccd1 vccd1 _4767_/C sky130_fd_sc_hd__nand2_1
X_5333_ _4604_/S _5339_/D _5979_/A vssd1 vssd1 vccd1 vccd1 _5333_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3173__A3 _4222_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5264_ _5317_/A _5264_/B vssd1 vssd1 vccd1 vccd1 _5266_/C sky130_fd_sc_hd__nor2_1
X_4215_ _3334_/C _5715_/C _4679_/D _5303_/A vssd1 vssd1 vccd1 vccd1 _4216_/B sky130_fd_sc_hd__a211oi_2
X_5195_ _6296_/Q _5082_/X _5194_/X _5371_/A _5102_/B vssd1 vssd1 vccd1 vccd1 _5195_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3243__A _4685_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3330__A0 _5715_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4146_ hold29/X _4425_/A2 _5597_/B vssd1 vssd1 vccd1 vccd1 _4146_/X sky130_fd_sc_hd__o21a_1
XANTENNA__3881__A1 _4427_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4077_ _4172_/C _4077_/B vssd1 vssd1 vccd1 vccd1 _5219_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4074__A _6247_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4979_ _6382_/Q _6330_/Q _6315_/Q vssd1 vssd1 vccd1 vccd1 _4979_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_61_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4521__B _5371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5310__B2 _5560_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5310__A1 _4221_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5613__A2 _4198_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3388__B1 _6389_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3927__A2 _3789_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6253__RESET_B fanout174/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5019__S _6315_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5301__A1 _5317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4104__A2 _3779_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4000_ _4000_/A _4000_/B vssd1 vssd1 vccd1 vccd1 _4001_/B sky130_fd_sc_hd__or2_2
X_5951_ _3625_/B _5950_/Y _4323_/A _5952_/B vssd1 vssd1 vccd1 vccd1 _5951_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_1_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4902_ _4900_/B _4901_/X _5058_/S vssd1 vssd1 vccd1 vccd1 _4902_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_75_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5882_ _6419_/Q _5881_/X _5930_/S vssd1 vssd1 vccd1 vccd1 _5882_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_75_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5368__A1 _5715_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4833_ _6419_/Q _4758_/X _4867_/B _4828_/Y _4831_/X vssd1 vssd1 vccd1 vccd1 _4833_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_83_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4764_ _3216_/A _3600_/B _5272_/B _4745_/C _3600_/A vssd1 vssd1 vccd1 vccd1 _4772_/B
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3715_ _3863_/A _3862_/S _3838_/S vssd1 vssd1 vccd1 vccd1 _3715_/X sky130_fd_sc_hd__and3_4
XANTENNA__6012__A2_N _6054_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4695_ _3909_/Y _4694_/X _4731_/S vssd1 vssd1 vccd1 vccd1 _4695_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_31_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6434_ _6440_/CLK _6434_/D fanout171/X vssd1 vssd1 vccd1 vccd1 _6434_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA_fanout114_A _4679_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3646_ _3424_/X _3645_/Y _5931_/S vssd1 vssd1 vccd1 vccd1 _3646_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_3_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3577_ _3577_/A _5956_/B vssd1 vssd1 vccd1 vccd1 _3605_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_60_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4974__S0 _5051_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6365_ _6384_/CLK _6365_/D fanout167/X vssd1 vssd1 vccd1 vccd1 _6365_/Q sky130_fd_sc_hd__dfrtp_2
X_5316_ _4541_/B _5265_/B _3573_/B _5480_/D _3572_/Y vssd1 vssd1 vccd1 vccd1 _5316_/X
+ sky130_fd_sc_hd__o221a_1
X_6296_ _6297_/CLK _6296_/D fanout176/X vssd1 vssd1 vccd1 vccd1 _6296_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_0_11_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4069__A _4070_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5247_ _5247_/A _5247_/B vssd1 vssd1 vccd1 vccd1 _5247_/X sky130_fd_sc_hd__or2_1
Xhold37 hold37/A vssd1 vssd1 vccd1 vccd1 hold37/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5603__D _5603_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold26 hold26/A vssd1 vssd1 vccd1 vccd1 hold26/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold15 hold15/A vssd1 vssd1 vccd1 vccd1 hold15/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold48 hold48/A vssd1 vssd1 vccd1 vccd1 hold48/X sky130_fd_sc_hd__dlygate4sd3_1
X_5178_ _5178_/A _5178_/B vssd1 vssd1 vccd1 vccd1 _5178_/Y sky130_fd_sc_hd__nor2_1
Xhold59 hold59/A vssd1 vssd1 vccd1 vccd1 hold59/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4129_ _4179_/A _4172_/B _4127_/X _3064_/Y vssd1 vssd1 vccd1 vccd1 _4129_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_97_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3611__A _3611_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xci2406_z80_205 vssd1 vssd1 vccd1 vccd1 ci2406_z80_205/HI io_oeb[34] sky130_fd_sc_hd__conb_1
XFILLER_0_16_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4161__B _6343_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3058__A _6246_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3500_ _4214_/A _3497_/X _3499_/X vssd1 vssd1 vccd1 vccd1 _3500_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_80_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5972__S _5975_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold518 _6385_/Q vssd1 vssd1 vccd1 vccd1 _5914_/A sky130_fd_sc_hd__dlygate4sd3_1
X_4480_ _4412_/X hold210/X _4482_/S vssd1 vssd1 vccd1 vccd1 _4480_/X sky130_fd_sc_hd__mux2_1
Xhold507 _4289_/X vssd1 vssd1 vccd1 vccd1 _6078_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3431_ _3431_/A _4284_/C vssd1 vssd1 vccd1 vccd1 _3431_/Y sky130_fd_sc_hd__nor2_1
Xhold529 _4533_/X vssd1 vssd1 vccd1 vccd1 _6234_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4956__S0 _5051_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3362_ _3611_/A _3362_/B vssd1 vssd1 vccd1 vccd1 _3362_/X sky130_fd_sc_hd__and2_1
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6150_ _6408_/CLK _6150_/D vssd1 vssd1 vccd1 vccd1 _6150_/Q sky130_fd_sc_hd__dfxtp_1
X_5101_ _6234_/Q _4520_/Y _5076_/A _5100_/Y vssd1 vssd1 vccd1 vccd1 _5101_/X sky130_fd_sc_hd__o22a_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3293_ _4744_/A _3293_/B _5303_/A vssd1 vssd1 vccd1 vccd1 _4747_/D sky130_fd_sc_hd__or3_4
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6081_ _6368_/CLK _6081_/D fanout169/X vssd1 vssd1 vccd1 vccd1 _6081_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3836__A1 _3850_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5032_ hold83/A _6158_/Q _6198_/Q _6074_/Q _5051_/S0 _5052_/S1 vssd1 vssd1 vccd1
+ vccd1 _5032_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_10_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6430_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__5038__A0 _6057_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4261__B2 _4228_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5934_ _5949_/C _6396_/Q vssd1 vssd1 vccd1 vccd1 _5934_/X sky130_fd_sc_hd__and2_1
X_5865_ _5865_/A _5926_/A vssd1 vssd1 vccd1 vccd1 _5889_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4352__A _4510_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5448__A _5715_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4816_ _5849_/S _4815_/X _4804_/X vssd1 vssd1 vccd1 vccd1 _4816_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_35_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5796_ _5813_/B _5796_/B vssd1 vssd1 vccd1 vccd1 _5796_/X sky130_fd_sc_hd__and2b_1
XANTENNA__4071__B _6247_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4747_ _3600_/A _3600_/B _4747_/C _4747_/D vssd1 vssd1 vccd1 vccd1 _4748_/D sky130_fd_sc_hd__and4bb_1
XFILLER_0_43_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4678_ _5989_/A _4678_/B vssd1 vssd1 vccd1 vccd1 _4731_/S sky130_fd_sc_hd__nand2_4
XFILLER_0_101_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3629_ _3683_/B _3629_/B vssd1 vssd1 vccd1 vccd1 _3634_/B sky130_fd_sc_hd__nand2_1
X_6417_ _6421_/CLK _6417_/D fanout175/X vssd1 vssd1 vccd1 vccd1 _6417_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__4498__S _4500_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5513__B2 _5377_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput38 _6262_/Q vssd1 vssd1 vccd1 vccd1 io_out[23] sky130_fd_sc_hd__buf_12
Xoutput49 _3647_/X vssd1 vssd1 vccd1 vccd1 io_out[3] sky130_fd_sc_hd__buf_12
Xoutput16 _6482_/X vssd1 vssd1 vccd1 vccd1 io_oeb[23] sky130_fd_sc_hd__buf_12
X_6348_ _6350_/CLK hold12/X vssd1 vssd1 vccd1 vccd1 hold11/A sky130_fd_sc_hd__dfxtp_1
Xoutput27 _6282_/Q vssd1 vssd1 vccd1 vccd1 io_out[13] sky130_fd_sc_hd__buf_12
XANTENNA__5277__B1 _3400_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6279_ _6376_/CLK _6279_/D fanout166/X vssd1 vssd1 vccd1 vccd1 _6279_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__3922__S1 _5676_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4252__A1 _4228_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4961__S _6315_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_hold610_A _6293_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3445__A_N _3473_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3325__B _4685_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3979__C _6245_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3294__A2 _3654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3980_ _4066_/B _3979_/X _6292_/Q vssd1 vssd1 vccd1 vccd1 _3981_/B sky130_fd_sc_hd__a21o_1
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4779__C1 _5054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5650_ _6095_/Q _4382_/B _4200_/S _6140_/Q _5673_/C1 vssd1 vssd1 vccd1 vccd1 _5651_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_45_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6059__A1_N _6022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4601_ _6422_/Q _4569_/X _4570_/X _6273_/Q _4600_/X vssd1 vssd1 vccd1 vccd1 _4601_/X
+ sky130_fd_sc_hd__a221o_1
X_5581_ _5270_/A _5728_/B _5324_/C _3599_/A vssd1 vssd1 vccd1 vccd1 _5581_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_72_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5743__A1 _5236_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4532_ hold490/X _4070_/A _4539_/S vssd1 vssd1 vccd1 vccd1 _4532_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_13_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4900__A _5054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold326 _3545_/B vssd1 vssd1 vccd1 vccd1 hold326/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold304 _6107_/Q vssd1 vssd1 vccd1 vccd1 hold304/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5715__B _5715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold315 _5340_/Y vssd1 vssd1 vccd1 vccd1 _6310_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4463_ _4420_/X hold89/X _4464_/S vssd1 vssd1 vccd1 vccd1 hold90/A sky130_fd_sc_hd__mux2_1
Xhold359 _6223_/Q vssd1 vssd1 vccd1 vccd1 hold359/X sky130_fd_sc_hd__dlygate4sd3_1
X_6202_ _6397_/CLK hold70/X fanout172/X vssd1 vssd1 vccd1 vccd1 hold69/A sky130_fd_sc_hd__dfrtp_1
X_3414_ _5265_/A _4284_/C _3414_/C _3414_/D vssd1 vssd1 vccd1 vccd1 _3415_/B sky130_fd_sc_hd__or4_1
XFILLER_0_68_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold348 _6262_/Q vssd1 vssd1 vccd1 vccd1 hold348/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold337 _5561_/Y vssd1 vssd1 vccd1 vccd1 _6335_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4394_ _4394_/A _4394_/B vssd1 vssd1 vccd1 vccd1 _4395_/B sky130_fd_sc_hd__xnor2_1
X_3345_ _5560_/A _3373_/A _5324_/A _5360_/C vssd1 vssd1 vccd1 vccd1 _3345_/X sky130_fd_sc_hd__or4b_1
XFILLER_0_68_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6133_ _6412_/CLK _6133_/D vssd1 vssd1 vccd1 vccd1 _6133_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3276_ _5270_/C _4734_/C vssd1 vssd1 vccd1 vccd1 _3600_/C sky130_fd_sc_hd__or2_2
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6064_ hold594/X _6063_/X _6064_/S vssd1 vssd1 vccd1 vccd1 _6448_/D sky130_fd_sc_hd__mux2_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5015_ _5014_/X _5013_/X _5053_/S vssd1 vssd1 vccd1 vccd1 _5016_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_84_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout181_A input14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4234__A1 _3656_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5917_ _5917_/A _5917_/B vssd1 vssd1 vccd1 vccd1 _5917_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_91_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5982__A1 _3577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5848_ _5848_/A _5848_/B vssd1 vssd1 vccd1 vccd1 _5848_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_90_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5734__B2 _3770_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5779_ _6374_/Q _5779_/B vssd1 vssd1 vccd1 vccd1 _5780_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_44_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout94_A _4313_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold658_A _6272_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4257__A _4541_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4225__A1 _3594_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3984__A0 _6244_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3433__C1 _4637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3671__A1_N _5097_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3130_ _5226_/A _3952_/A vssd1 vssd1 vccd1 vccd1 _3374_/A sky130_fd_sc_hd__nand2b_4
X_3061_ _3061_/A vssd1 vssd1 vccd1 vccd1 _3061_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_89_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5639__S1 _5690_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3963_ hold19/X _4425_/A2 _3962_/X vssd1 vssd1 vccd1 vccd1 _3963_/X sky130_fd_sc_hd__o21a_1
X_3894_ _6242_/Q _6244_/Q _4135_/S vssd1 vssd1 vccd1 vccd1 _5130_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_70_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5702_ hold11/X _3826_/B _6060_/S vssd1 vssd1 vccd1 vccd1 hold12/A sky130_fd_sc_hd__mux2_1
X_5633_ _6410_/Q _4382_/B _4384_/S _6179_/Q _5675_/C1 vssd1 vssd1 vccd1 vccd1 _5635_/A
+ sky130_fd_sc_hd__o221a_1
X_5564_ _4541_/C _5562_/X _5563_/X _4274_/A vssd1 vssd1 vccd1 vccd1 _5564_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_60_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold101 _6089_/Q vssd1 vssd1 vccd1 vccd1 hold101/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4515_ _4054_/X hold212/X _4518_/S vssd1 vssd1 vccd1 vccd1 _4515_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_13_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold112 _4459_/X vssd1 vssd1 vccd1 vccd1 _6162_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold123 _4518_/X vssd1 vssd1 vccd1 vccd1 _6222_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5495_ _6417_/Q _5558_/S _5494_/X vssd1 vssd1 vccd1 vccd1 _5495_/X sky130_fd_sc_hd__o21ba_1
Xhold134 _6115_/Q vssd1 vssd1 vccd1 vccd1 hold134/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold167 _6161_/Q vssd1 vssd1 vccd1 vccd1 hold167/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold156 _4477_/X vssd1 vssd1 vccd1 vccd1 _6178_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold145 _6096_/Q vssd1 vssd1 vccd1 vccd1 hold145/X sky130_fd_sc_hd__dlygate4sd3_1
X_4446_ hold65/X _4427_/X _4446_/S vssd1 vssd1 vccd1 vccd1 hold66/A sky130_fd_sc_hd__mux2_1
X_4377_ _5249_/A _5249_/B _3723_/X vssd1 vssd1 vccd1 vccd1 _4377_/X sky130_fd_sc_hd__o21a_1
XANTENNA__4152__B1 _3781_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold189 _6212_/Q vssd1 vssd1 vccd1 vccd1 hold189/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold178 _4506_/X vssd1 vssd1 vccd1 vccd1 _6211_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_95_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3328_ _3525_/A _3525_/B _6293_/Q _3334_/C vssd1 vssd1 vccd1 vccd1 _3328_/Y sky130_fd_sc_hd__nor4b_1
X_6116_ _6432_/CLK _6116_/D fanout173/X vssd1 vssd1 vccd1 vccd1 _6116_/Q sky130_fd_sc_hd__dfstp_1
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3259_ _5096_/A _6389_/Q vssd1 vssd1 vccd1 vccd1 _3770_/A sky130_fd_sc_hd__or2_4
X_6047_ _6057_/A _6046_/X _6063_/S vssd1 vssd1 vccd1 vccd1 _6047_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_95_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5404__A0 _6418_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5339__C _5339_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4391__B1 _5597_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4686__S _4727_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5486__A3 _5484_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5371__A _5371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_26_wb_clk_i_A _6404_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5280_ _3656_/A _5278_/X _3357_/C vssd1 vssd1 vccd1 vccd1 _5280_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_2_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4300_ _4313_/C _4307_/B vssd1 vssd1 vccd1 vccd1 _4304_/B sky130_fd_sc_hd__nand2_1
X_4231_ _4224_/A _3511_/A _4224_/C _4230_/X vssd1 vssd1 vccd1 vccd1 _5343_/B sky130_fd_sc_hd__a31o_1
XFILLER_0_49_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5882__A0 _6419_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4162_ _4163_/A _5107_/B vssd1 vssd1 vccd1 vccd1 _4162_/X sky130_fd_sc_hd__or2_1
XFILLER_0_65_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3113_ _4744_/A _3289_/A _6254_/Q _3183_/B vssd1 vssd1 vccd1 vccd1 _3285_/B sky130_fd_sc_hd__or4b_4
X_4093_ _4093_/A _4093_/B vssd1 vssd1 vccd1 vccd1 _4095_/B sky130_fd_sc_hd__nor2_2
X_3044_ _5553_/S vssd1 vssd1 vccd1 vccd1 _5715_/A sky130_fd_sc_hd__inv_4
XANTENNA__4625__A input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3660__A2 _3654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4995_ _4994_/X _4993_/X _5053_/S vssd1 vssd1 vccd1 vccd1 _4996_/B sky130_fd_sc_hd__mux2_2
XANTENNA_fanout144_A _3482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3946_ _6292_/Q _3886_/A _4073_/B vssd1 vssd1 vccd1 vccd1 _3948_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_45_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3877_ _3877_/A _3877_/B _3877_/C vssd1 vssd1 vccd1 vccd1 _3878_/B sky130_fd_sc_hd__and3_1
X_5616_ _5615_/X _3922_/X _5690_/S vssd1 vssd1 vccd1 vccd1 _5616_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_26_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5547_ _6333_/Q _5377_/X _5546_/X _5377_/A vssd1 vssd1 vccd1 vccd1 _5547_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_5_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5478_ _5478_/A _5478_/B vssd1 vssd1 vccd1 vccd1 _5478_/Y sky130_fd_sc_hd__xnor2_1
X_4429_ _4510_/A _4501_/A vssd1 vssd1 vccd1 vccd1 _4437_/S sky130_fd_sc_hd__nor2_4
XANTENNA__5873__A0 _6418_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4519__B _4520_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6300__RESET_B fanout179/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5625__B1 _5676_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3651__A2 _5975_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout73 _3720_/X vssd1 vssd1 vccd1 vccd1 _5673_/C1 sky130_fd_sc_hd__buf_6
XFILLER_0_9_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout62 _5825_/S vssd1 vssd1 vccd1 vccd1 _5928_/A2 sky130_fd_sc_hd__buf_4
XANTENNA__3585__S _4309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout84 _4197_/B vssd1 vssd1 vccd1 vccd1 _5597_/B sky130_fd_sc_hd__buf_4
XFILLER_0_24_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout95 _3475_/X vssd1 vssd1 vccd1 vccd1 _4313_/C sky130_fd_sc_hd__buf_4
XFILLER_0_101_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5084__A1_N _4070_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4903__A2 _6325_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4667__A1 _5715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4164__B _6343_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5975__S _5975_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3800_ hold71/X _3779_/X _3781_/X hold65/X vssd1 vssd1 vccd1 vccd1 _3804_/A sky130_fd_sc_hd__a22o_1
X_4780_ _6319_/Q _5728_/D _4742_/X _4779_/X _5740_/A vssd1 vssd1 vccd1 vccd1 _4780_/X
+ sky130_fd_sc_hd__a221o_1
X_3731_ _6242_/Q _6336_/Q _3938_/A vssd1 vssd1 vccd1 vccd1 _3731_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_51_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_35_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6376_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_27_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3662_ _3657_/A _3657_/B _3553_/Y _3287_/Y _3658_/Y vssd1 vssd1 vccd1 vccd1 _3662_/X
+ sky130_fd_sc_hd__a221o_1
X_3593_ _4520_/B _3686_/C _5323_/C _4541_/D vssd1 vssd1 vccd1 vccd1 _5481_/C sky130_fd_sc_hd__or4_1
X_5401_ hold585/X _5377_/X _5400_/Y _5441_/A vssd1 vssd1 vccd1 vccd1 _5401_/X sky130_fd_sc_hd__a22o_1
X_6381_ _6386_/CLK _6381_/D fanout167/X vssd1 vssd1 vccd1 vccd1 _6381_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_2_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5332_ _5339_/D vssd1 vssd1 vccd1 vccd1 _5332_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_11_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4107__B1 _3794_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5263_ _5257_/X _5262_/X _6118_/Q vssd1 vssd1 vccd1 vccd1 _5263_/X sky130_fd_sc_hd__o21a_1
XANTENNA__3524__A _6118_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4214_ _4214_/A _4214_/B _5258_/B vssd1 vssd1 vccd1 vccd1 _4216_/A sky130_fd_sc_hd__and3_1
XFILLER_0_76_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5194_ _6238_/Q _5075_/B _5076_/Y _5193_/X vssd1 vssd1 vccd1 vccd1 _5194_/X sky130_fd_sc_hd__a22o_1
X_4145_ _3724_/A _4115_/X _4144_/X vssd1 vssd1 vccd1 vccd1 _4145_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_92_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4076_ _4128_/A _4177_/A _6292_/Q vssd1 vssd1 vccd1 vccd1 _4077_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_78_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5885__S _5933_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4978_ _6444_/Q _5056_/A2 _4977_/X vssd1 vssd1 vccd1 vccd1 _4978_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_18_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3929_ _3929_/A _3929_/B vssd1 vssd1 vccd1 vccd1 _3930_/B sky130_fd_sc_hd__or2_2
XANTENNA__4521__C _5075_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4649__A1 _6342_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3434__A _5935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4964__S _5060_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3085__B1 _5935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5096__A _5096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4888__B2 _4882_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3560__A1 _3502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3312__A1 _4214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5950_ _5952_/A _3466_/B _3620_/B _5949_/X vssd1 vssd1 vccd1 vccd1 _5950_/Y sky130_fd_sc_hd__a31oi_1
XFILLER_0_87_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4901_ _6378_/Q _6326_/Q _4901_/S vssd1 vssd1 vccd1 vccd1 _4901_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4812__B2 _4807_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5881_ _5929_/A1 _5880_/X _4976_/Y vssd1 vssd1 vccd1 vccd1 _5881_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_75_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5368__A2 _6416_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4832_ _6436_/Q _4756_/Y _4757_/Y _4830_/B _4754_/X vssd1 vssd1 vccd1 vccd1 _4832_/X
+ sky130_fd_sc_hd__a221o_1
X_4763_ _3361_/A _4763_/B vssd1 vssd1 vccd1 vccd1 _4867_/B sky130_fd_sc_hd__and2b_4
XFILLER_0_43_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3519__A _5733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3714_ _3699_/Y _3704_/S _3711_/Y _3712_/X vssd1 vssd1 vccd1 vccd1 _3838_/S sky130_fd_sc_hd__a31oi_4
X_4694_ _4692_/X _4693_/X _5102_/A vssd1 vssd1 vccd1 vccd1 _4694_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_43_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6433_ _6433_/CLK _6433_/D fanout171/X vssd1 vssd1 vccd1 vccd1 _6433_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_0_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3645_ _3645_/A _3645_/B vssd1 vssd1 vccd1 vccd1 _3645_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_3_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3576_ _3459_/Y _3575_/X _5313_/A vssd1 vssd1 vccd1 vccd1 _3583_/B sky130_fd_sc_hd__a21oi_2
XANTENNA_fanout107_A _4732_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4974__S1 _5052_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6364_ _6376_/CLK _6364_/D fanout166/X vssd1 vssd1 vccd1 vccd1 _6364_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_0_23_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5315_ _5315_/A _5315_/B _5343_/C vssd1 vssd1 vccd1 vccd1 _5315_/X sky130_fd_sc_hd__or3_1
X_6295_ _6295_/CLK _6295_/D fanout177/X vssd1 vssd1 vccd1 vccd1 _6295_/Q sky130_fd_sc_hd__dfstp_2
XANTENNA__3254__A _3254_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5246_ _5249_/D vssd1 vssd1 vccd1 vccd1 _5246_/Y sky130_fd_sc_hd__inv_2
Xhold38 hold38/A vssd1 vssd1 vccd1 vccd1 hold38/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold27 hold27/A vssd1 vssd1 vccd1 vccd1 hold27/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold16 hold16/A vssd1 vssd1 vccd1 vccd1 hold16/X sky130_fd_sc_hd__dlygate4sd3_1
X_5177_ _3759_/A _5174_/X _5176_/X vssd1 vssd1 vccd1 vccd1 _5178_/B sky130_fd_sc_hd__a21oi_1
Xhold49 hold49/A vssd1 vssd1 vccd1 vccd1 hold49/X sky130_fd_sc_hd__dlygate4sd3_1
X_4128_ _4128_/A _4128_/B vssd1 vssd1 vccd1 vccd1 _4172_/B sky130_fd_sc_hd__nand2_1
X_4059_ _4059_/A _4059_/B vssd1 vssd1 vccd1 vccd1 _4061_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_78_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold590_A _6326_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3542__B2 _5313_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5295__B2 _4228_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3845__A2 _3838_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3611__B _5715_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xci2406_z80_206 vssd1 vssd1 vccd1 vccd1 ci2406_z80_206/HI io_out[4] sky130_fd_sc_hd__conb_1
XFILLER_0_16_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5598__A2 _5690_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3230__B1 _3566_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6403__RESET_B fanout180/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold508 _6446_/Q vssd1 vssd1 vccd1 vccd1 hold508/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4869__S _5058_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3430_ _3394_/C _3392_/Y _3428_/X _3429_/X _3686_/A vssd1 vssd1 vccd1 vccd1 _3434_/C
+ sky130_fd_sc_hd__o41a_1
XANTENNA__4956__S1 _5052_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold519 _5923_/X vssd1 vssd1 vccd1 vccd1 _6385_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3533__B2 _6390_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3361_ _3361_/A _4763_/B vssd1 vssd1 vccd1 vccd1 _3361_/X sky130_fd_sc_hd__and2_1
X_5100_ _3064_/Y _5192_/S _5193_/S vssd1 vssd1 vccd1 vccd1 _5100_/Y sky130_fd_sc_hd__a21boi_1
XANTENNA__3074__A _6270_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6080_ _6368_/CLK _6080_/D fanout169/X vssd1 vssd1 vccd1 vccd1 _6080_/Q sky130_fd_sc_hd__dfrtp_1
X_3292_ _4744_/A _4744_/B _3292_/C vssd1 vssd1 vccd1 vccd1 _5324_/A sky130_fd_sc_hd__and3b_2
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4089__A2 _3779_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5031_ hold99/A hold79/A _6097_/Q _6142_/Q _5051_/S0 _5052_/S1 vssd1 vssd1 vccd1
+ vccd1 _5031_/X sky130_fd_sc_hd__mux4_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4261__A2 _3654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_50_wb_clk_i clkbuf_leaf_6_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6217_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_5933_ _5925_/A _5932_/X _5933_/S vssd1 vssd1 vccd1 vccd1 _5933_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_8_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5864_ _5856_/A _5742_/Y _5863_/X _5933_/S vssd1 vssd1 vccd1 vccd1 _5864_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5448__B _6422_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4815_ _6373_/Q _4796_/B _4812_/X _4814_/X vssd1 vssd1 vccd1 vccd1 _4815_/X sky130_fd_sc_hd__o22a_1
XANTENNA__3249__A _5313_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4013__A2 _3779_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5795_ _5795_/A _5795_/B _5793_/X vssd1 vssd1 vccd1 vccd1 _5796_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_90_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4746_ _5376_/B vssd1 vssd1 vccd1 vccd1 _4746_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_71_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5761__A2 _5728_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4677_ _5715_/B _4673_/Y _4676_/X hold332/X _4635_/Y vssd1 vssd1 vccd1 vccd1 _4677_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_0_31_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3628_ _5560_/A _3628_/B vssd1 vssd1 vccd1 vccd1 _3629_/B sky130_fd_sc_hd__nor2_1
X_6416_ _6423_/CLK _6416_/D fanout175/X vssd1 vssd1 vccd1 vccd1 _6416_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_31_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput39 _6264_/Q vssd1 vssd1 vccd1 vccd1 io_out[24] sky130_fd_sc_hd__buf_12
Xoutput17 _6483_/X vssd1 vssd1 vccd1 vccd1 io_oeb[24] sky130_fd_sc_hd__buf_12
X_6347_ _6350_/CLK hold16/X vssd1 vssd1 vccd1 vccd1 hold15/A sky130_fd_sc_hd__dfxtp_1
Xoutput28 _6283_/Q vssd1 vssd1 vccd1 vccd1 io_out[14] sky130_fd_sc_hd__buf_12
X_3559_ _3559_/A _3559_/B _3559_/C _3551_/X vssd1 vssd1 vccd1 vccd1 _3561_/B sky130_fd_sc_hd__or4b_1
XANTENNA__5277__A1 _3337_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6278_ _6376_/CLK _6278_/D fanout166/X vssd1 vssd1 vccd1 vccd1 _6278_/Q sky130_fd_sc_hd__dfrtp_1
X_5229_ _6417_/Q _6416_/Q _6421_/Q _6420_/Q vssd1 vssd1 vccd1 vccd1 _5229_/X sky130_fd_sc_hd__or4_1
XANTENNA__5403__S _5560_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3827__A2 _3784_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3431__B _4284_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4252__A2 _3654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5737__C1 _6392_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold603_A _6380_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3763__A1 _6242_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5268__A1 _4224_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4600_ _4111_/B _4604_/S _4564_/A _4599_/Y vssd1 vssd1 vccd1 vccd1 _4600_/X sky130_fd_sc_hd__o211a_1
X_5580_ _3183_/B _3373_/A _3661_/A _4208_/B _5579_/X vssd1 vssd1 vccd1 vccd1 _5580_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_72_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4531_ hold445/X _6274_/Q _4539_/S vssd1 vssd1 vccd1 vccd1 _4531_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_4_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4900__B _4900_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5284__A _6389_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5715__C _5715_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold316 _6249_/Q vssd1 vssd1 vccd1 vccd1 hold316/X sky130_fd_sc_hd__dlygate4sd3_1
X_4462_ _4412_/X hold228/X _4464_/S vssd1 vssd1 vccd1 vccd1 _6165_/D sky130_fd_sc_hd__mux2_1
Xhold305 _6414_/Q vssd1 vssd1 vccd1 vccd1 hold305/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold327 _3508_/X vssd1 vssd1 vccd1 vccd1 _6397_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6201_ _6397_/CLK hold34/X fanout172/X vssd1 vssd1 vccd1 vccd1 hold33/A sky130_fd_sc_hd__dfrtp_1
X_3413_ _3572_/A _3654_/A _4767_/B _3431_/A _4260_/A vssd1 vssd1 vccd1 vccd1 _3414_/D
+ sky130_fd_sc_hd__a221o_1
Xhold349 _4657_/X vssd1 vssd1 vccd1 vccd1 _6262_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold338 _6277_/Q vssd1 vssd1 vccd1 vccd1 hold338/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5051__S0 _5051_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4703__B1 _5075_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4393_ hold45/X _4392_/X _4428_/S vssd1 vssd1 vccd1 vccd1 hold46/A sky130_fd_sc_hd__mux2_1
X_3344_ _3344_/A _5256_/A vssd1 vssd1 vccd1 vccd1 _5481_/A sky130_fd_sc_hd__nand2_2
X_6132_ _6410_/CLK _6132_/D vssd1 vssd1 vccd1 vccd1 _6132_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3275_ _3290_/B _3369_/B vssd1 vssd1 vccd1 vccd1 _4734_/C sky130_fd_sc_hd__nor2_1
X_6063_ _4193_/Y _6062_/X _6063_/S vssd1 vssd1 vccd1 vccd1 _6063_/X sky130_fd_sc_hd__mux2_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5014_ _6220_/Q hold85/A _6197_/Q _6073_/Q _5358_/A0 _4326_/B vssd1 vssd1 vccd1 vccd1
+ _5014_/X sky130_fd_sc_hd__mux4_1
XANTENNA__3809__A2 _3715_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3251__B _3725_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout174_A fanout181/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5431__B2 _5740_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5916_ _5906_/A _5909_/B _5907_/A vssd1 vssd1 vccd1 vccd1 _5917_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_75_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6396__RESET_B fanout173/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6325__RESET_B fanout174/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5847_ _5846_/A _5846_/B _5848_/A vssd1 vssd1 vccd1 vccd1 _5847_/X sky130_fd_sc_hd__o21ba_1
XANTENNA__5734__A2 _4767_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5778_ _5778_/A _5779_/B vssd1 vssd1 vccd1 vccd1 _5795_/A sky130_fd_sc_hd__and2_1
XANTENNA__4942__A0 _4938_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4729_ _6274_/Q _4681_/X _4728_/X _5371_/A vssd1 vssd1 vccd1 vccd1 _4729_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_31_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3442__A _5931_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_16_wb_clk_i_A _6404_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5369__A _6392_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3984__A1 _6246_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6126__SET_B fanout180/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5832__A _6378_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3060_ _6248_/Q vssd1 vssd1 vccd1 vccd1 _4130_/A sky130_fd_sc_hd__inv_2
XFILLER_0_89_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4183__A _4679_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5701_ hold15/X _4394_/B _6060_/S vssd1 vssd1 vccd1 vccd1 hold16/A sky130_fd_sc_hd__mux2_1
X_3962_ _3724_/A _5252_/B _3961_/Y vssd1 vssd1 vccd1 vccd1 _3962_/X sky130_fd_sc_hd__a21o_1
X_3893_ _6337_/Q _6341_/Q _6301_/Q vssd1 vssd1 vccd1 vccd1 _5216_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_73_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5632_ _5695_/A1 _3061_/A _5571_/Y _5631_/X vssd1 vssd1 vccd1 vccd1 _5632_/X sky130_fd_sc_hd__a22o_1
X_5563_ _5563_/A _5563_/B _5563_/C vssd1 vssd1 vccd1 vccd1 _5563_/X sky130_fd_sc_hd__or3_1
XFILLER_0_72_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4924__A0 _4920_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4514_ _4007_/X hold231/X _4518_/S vssd1 vssd1 vccd1 vccd1 _4514_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold113 _6300_/Q vssd1 vssd1 vccd1 vccd1 hold113/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold102 _3527_/X vssd1 vssd1 vccd1 vccd1 _6089_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold124 _6207_/Q vssd1 vssd1 vccd1 vccd1 hold124/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold135 _4360_/X vssd1 vssd1 vccd1 vccd1 _6115_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5494_ _6057_/A _5377_/A _5492_/Y _5493_/Y _5558_/S vssd1 vssd1 vccd1 vccd1 _5494_/X
+ sky130_fd_sc_hd__o311a_1
Xhold168 _4458_/X vssd1 vssd1 vccd1 vccd1 _6161_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold146 _4334_/X vssd1 vssd1 vccd1 vccd1 _6096_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold157 _6368_/Q vssd1 vssd1 vccd1 vccd1 hold157/X sky130_fd_sc_hd__dlygate4sd3_1
X_4445_ hold136/X _4420_/X _4446_/S vssd1 vssd1 vccd1 vccd1 _4445_/X sky130_fd_sc_hd__mux2_1
X_4376_ _5249_/A _5249_/B vssd1 vssd1 vccd1 vccd1 _4376_/Y sky130_fd_sc_hd__nand2_1
Xhold179 _6215_/Q vssd1 vssd1 vccd1 vccd1 hold179/X sky130_fd_sc_hd__dlygate4sd3_1
X_3327_ _3525_/A _3374_/A vssd1 vssd1 vccd1 vccd1 _4042_/A sky130_fd_sc_hd__nor2_1
X_6115_ _6444_/CLK _6115_/D vssd1 vssd1 vccd1 vccd1 _6115_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3258_ _5096_/A _6389_/Q vssd1 vssd1 vccd1 vccd1 _3581_/A sky130_fd_sc_hd__nor2_4
X_6046_ _5524_/X _6054_/B _6057_/B _4996_/B vssd1 vssd1 vccd1 vccd1 _6046_/X sky130_fd_sc_hd__o2bb2a_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3189_ _4520_/B _3189_/B _3189_/C vssd1 vssd1 vccd1 vccd1 _3196_/A sky130_fd_sc_hd__or3_1
XFILLER_0_76_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5955__A2 _3639_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5168__B1 _5447_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold670_A _6118_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold680 _6311_/Q vssd1 vssd1 vccd1 vccd1 hold680/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5371__B _5441_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3172__A _5935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5643__A1 _6270_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6483__A _6487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6404__CLK _6404_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5038__S _5058_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4877__S _5029_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4230_ _5096_/A _3409_/B _3343_/Y vssd1 vssd1 vccd1 vccd1 _4230_/X sky130_fd_sc_hd__o21a_1
X_4161_ _5088_/B _6343_/Q vssd1 vssd1 vccd1 vccd1 _5107_/B sky130_fd_sc_hd__xor2_1
XANTENNA__3893__A0 _6337_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3112_ _3254_/A _3136_/B _3289_/A vssd1 vssd1 vccd1 vccd1 _4257_/B sky130_fd_sc_hd__or3_2
X_4092_ _6073_/Q _3715_/X _3794_/X _6141_/Q _4091_/X vssd1 vssd1 vccd1 vccd1 _4093_/B
+ sky130_fd_sc_hd__a221o_1
X_3043_ _3043_/A vssd1 vssd1 vccd1 vccd1 _4558_/A sky130_fd_sc_hd__inv_2
XANTENNA__4625__B _4631_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4994_ _6219_/Q _6156_/Q _6196_/Q _6072_/Q _5051_/S0 _4326_/B vssd1 vssd1 vccd1 vccd1
+ _4994_/X sky130_fd_sc_hd__mux4_1
X_3945_ _3938_/A _3939_/A _3061_/Y _3760_/B _3944_/Y vssd1 vssd1 vccd1 vccd1 _5112_/A
+ sky130_fd_sc_hd__a41o_1
XFILLER_0_73_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5615_ _5615_/A _5615_/B vssd1 vssd1 vccd1 vccd1 _5615_/X sky130_fd_sc_hd__or2_1
XFILLER_0_33_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3876_ _3877_/B _3877_/C _3877_/A vssd1 vssd1 vccd1 vccd1 _3876_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_83_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5570__B1 _5339_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5546_ _5546_/A _5546_/B vssd1 vssd1 vccd1 vccd1 _5546_/X sky130_fd_sc_hd__xor2_1
XANTENNA__4787__S _4901_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5477_ _5477_/A _5477_/B vssd1 vssd1 vccd1 vccd1 _5478_/B sky130_fd_sc_hd__nor2_1
X_4428_ hold259/X _4427_/X _4428_/S vssd1 vssd1 vccd1 vccd1 _4428_/X sky130_fd_sc_hd__mux2_1
X_4359_ hold99/X _4148_/X _4360_/S vssd1 vssd1 vccd1 vccd1 _4359_/X sky130_fd_sc_hd__mux2_1
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6029_ _5994_/A _6063_/S _3046_/A vssd1 vssd1 vccd1 vccd1 _6029_/Y sky130_fd_sc_hd__a21oi_4
Xclkbuf_leaf_5_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6408_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_96_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6050__A1 _6057_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout74 _5989_/X vssd1 vssd1 vccd1 vccd1 _6026_/B sky130_fd_sc_hd__buf_4
Xfanout63 _5772_/S vssd1 vssd1 vccd1 vccd1 _5825_/S sky130_fd_sc_hd__buf_4
XFILLER_0_9_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4600__A2 _4604_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout96 _5740_/A vssd1 vssd1 vccd1 vccd1 _5560_/D sky130_fd_sc_hd__buf_4
Xfanout85 _3684_/X vssd1 vssd1 vccd1 vccd1 _4427_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_0_9_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3167__A _3482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4697__S _4727_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5864__B2 _5933_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6081__RESET_B fanout169/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3722__S0 _5676_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4052__B1 _5597_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3730_ _3938_/A _6336_/Q vssd1 vssd1 vccd1 vccd1 _3732_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3130__A_N _5226_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3661_ _3661_/A _5563_/A vssd1 vssd1 vccd1 vccd1 _3661_/X sky130_fd_sc_hd__or2_1
X_3592_ _3592_/A _3592_/B vssd1 vssd1 vccd1 vccd1 _4768_/A sky130_fd_sc_hd__nor2_1
X_5400_ _5400_/A vssd1 vssd1 vccd1 vccd1 _5400_/Y sky130_fd_sc_hd__inv_2
X_6380_ _6384_/CLK _6380_/D fanout167/X vssd1 vssd1 vccd1 vccd1 _6380_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_2_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5331_ _5317_/A _5096_/B _5330_/X _3686_/A vssd1 vssd1 vccd1 vccd1 _5339_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_100_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4400__S _4428_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5262_ _3549_/A _5578_/A _5258_/Y _5261_/Y vssd1 vssd1 vccd1 vccd1 _5262_/X sky130_fd_sc_hd__o22a_1
XANTENNA__3524__B _5258_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4213_ _5258_/B _4346_/B _3233_/D vssd1 vssd1 vccd1 vccd1 _5315_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_76_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5193_ _6272_/Q _5192_/X _5193_/S vssd1 vssd1 vccd1 vccd1 _5193_/X sky130_fd_sc_hd__mux2_1
X_4144_ _3724_/A _6022_/A _4425_/A2 vssd1 vssd1 vccd1 vccd1 _4144_/X sky130_fd_sc_hd__o21a_1
XANTENNA__5607__A1 _6416_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4075_ _4075_/A _4075_/B vssd1 vssd1 vccd1 vccd1 _4177_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__4636__A _6032_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3618__B1 _4750_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4291__B1 _4316_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4977_ _6270_/Q _4758_/X _4976_/B _4757_/Y vssd1 vssd1 vccd1 vccd1 _4977_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_18_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3928_ _6070_/Q _3715_/X _3794_/X _6138_/Q _3927_/X vssd1 vssd1 vccd1 vccd1 _3929_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_73_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3859_ _3850_/B _3856_/X _3858_/X vssd1 vssd1 vccd1 vccd1 _3864_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_6_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5529_ _5526_/A _5528_/X _6060_/S vssd1 vssd1 vccd1 vccd1 _5529_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_5_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5074__A2 _5247_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4980__S _5058_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4821__A2 _5557_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5377__A _5377_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4585__A1 _6419_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4585__B2 _6270_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5096__B _5096_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3328__C _6293_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6262__RESET_B fanout177/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5880_ _6330_/Q _5928_/A2 _5928_/B1 _5879_/X vssd1 vssd1 vccd1 vccd1 _5880_/X sky130_fd_sc_hd__a22o_1
X_4900_ _5054_/A _4900_/B vssd1 vssd1 vccd1 vccd1 _4900_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_75_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4831_ _3365_/B _4829_/X _4830_/X _5061_/A1 vssd1 vssd1 vccd1 vccd1 _4831_/X sky130_fd_sc_hd__o211a_1
XANTENNA__5368__A3 _5365_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4762_ _5365_/C _4761_/X _4762_/S vssd1 vssd1 vccd1 vccd1 _4762_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4576__B2 _6268_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4576__A1 _6417_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3713_ _3699_/Y _3704_/S _3711_/Y _3712_/X vssd1 vssd1 vccd1 vccd1 _3861_/S sky130_fd_sc_hd__a31o_4
X_4693_ hold377/X _4298_/B _4727_/S vssd1 vssd1 vccd1 vccd1 _4693_/X sky130_fd_sc_hd__mux2_1
X_3644_ _3048_/Y _5728_/B _3643_/X vssd1 vssd1 vccd1 vccd1 _3644_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_70_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6432_ _6432_/CLK _6432_/D fanout178/X vssd1 vssd1 vccd1 vccd1 _6432_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3535__A _4685_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3575_ _3570_/X _3571_/X _3572_/Y _3574_/Y _3686_/A vssd1 vssd1 vccd1 vccd1 _3575_/X
+ sky130_fd_sc_hd__a41o_1
X_6363_ _6384_/CLK _6363_/D fanout167/X vssd1 vssd1 vccd1 vccd1 _6363_/Q sky130_fd_sc_hd__dfrtp_2
X_5314_ _5314_/A _5563_/B vssd1 vssd1 vccd1 vccd1 _5343_/C sky130_fd_sc_hd__or2_1
X_6294_ _6295_/CLK _6294_/D fanout177/X vssd1 vssd1 vccd1 vccd1 _6294_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_0_11_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3254__B _3566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5245_ _3473_/A _3697_/X _3680_/X _3674_/B _3674_/A vssd1 vssd1 vccd1 vccd1 _5249_/D
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_0_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold28 hold28/A vssd1 vssd1 vccd1 vccd1 hold28/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold17 hold17/A vssd1 vssd1 vccd1 vccd1 hold17/X sky130_fd_sc_hd__dlygate4sd3_1
X_5176_ _6294_/Q _5149_/X _5175_/X _3986_/X _5241_/S vssd1 vssd1 vccd1 vccd1 _5176_/X
+ sky130_fd_sc_hd__a2111o_1
Xhold39 hold39/A vssd1 vssd1 vccd1 vccd1 hold39/X sky130_fd_sc_hd__dlygate4sd3_1
X_4127_ _4172_/C _4128_/A _4128_/B vssd1 vssd1 vccd1 vccd1 _4127_/X sky130_fd_sc_hd__a21o_1
X_4058_ _6247_/Q _4058_/B vssd1 vssd1 vccd1 vccd1 _4061_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6005__A1 _5560_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4016__B1 _3794_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4305__S _4305_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5764__B1 _5735_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold583_A _6381_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6291__SET_B fanout177/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4975__S _5053_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5295__A2 _3400_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xci2406_z80_207 vssd1 vssd1 vccd1 vccd1 ci2406_z80_207/HI io_out[30] sky130_fd_sc_hd__conb_1
XANTENNA__5678__S0 _5691_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5507__A0 _6418_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold509 _6053_/X vssd1 vssd1 vccd1 vccd1 _6446_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3360_ _4755_/A _4757_/B vssd1 vssd1 vccd1 vccd1 _4763_/B sky130_fd_sc_hd__and2b_1
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4885__S _5058_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3291_ _3386_/A _3657_/A vssd1 vssd1 vccd1 vccd1 _5360_/B sky130_fd_sc_hd__nor2_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5030_ hold403/X _5029_/X _5068_/S vssd1 vssd1 vccd1 vccd1 _5030_/X sky130_fd_sc_hd__mux2_1
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5932_ _5926_/X _5931_/X _5932_/S vssd1 vssd1 vccd1 vccd1 _5932_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_87_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5863_ _5932_/S _5858_/Y _5862_/X _5747_/Y vssd1 vssd1 vccd1 vccd1 _5863_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_75_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5794_ _5795_/A _5795_/B _5793_/X vssd1 vssd1 vccd1 vccd1 _5813_/B sky130_fd_sc_hd__o21ba_1
X_4814_ _4867_/B _4808_/X _4828_/B _4813_/X vssd1 vssd1 vccd1 vccd1 _4814_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_90_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4745_ _5560_/A _4745_/B _4745_/C _4744_/X vssd1 vssd1 vccd1 vccd1 _5376_/B sky130_fd_sc_hd__or4b_2
XFILLER_0_56_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4676_ _3691_/B _4675_/X _4673_/B vssd1 vssd1 vccd1 vccd1 _4676_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_31_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3627_ _3639_/B _3639_/C vssd1 vssd1 vccd1 vccd1 _3627_/Y sky130_fd_sc_hd__nor2_1
X_6415_ _6423_/CLK _6415_/D fanout175/X vssd1 vssd1 vccd1 vccd1 _6415_/Q sky130_fd_sc_hd__dfstp_2
X_3558_ _3553_/Y _3554_/X _3555_/Y _4224_/C _3557_/Y vssd1 vssd1 vccd1 vccd1 _3559_/B
+ sky130_fd_sc_hd__a221o_1
X_6346_ _6351_/CLK hold24/X vssd1 vssd1 vccd1 vccd1 hold23/A sky130_fd_sc_hd__dfxtp_1
Xoutput29 _6284_/Q vssd1 vssd1 vccd1 vccd1 io_out[15] sky130_fd_sc_hd__buf_12
Xoutput18 _6484_/X vssd1 vssd1 vccd1 vccd1 io_oeb[25] sky130_fd_sc_hd__buf_12
XFILLER_0_11_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5277__A2 _3502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5480__A _5560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3489_ _3611_/A _5472_/S _5739_/A vssd1 vssd1 vccd1 vccd1 _3505_/B sky130_fd_sc_hd__and3_1
X_6277_ _6376_/CLK _6277_/D fanout166/X vssd1 vssd1 vccd1 vccd1 _6277_/Q sky130_fd_sc_hd__dfrtp_1
X_5228_ _5221_/X _5227_/X _5241_/S vssd1 vssd1 vccd1 vccd1 _5228_/X sky130_fd_sc_hd__mux2_1
X_5159_ _6421_/Q _6420_/Q vssd1 vssd1 vccd1 vccd1 _5165_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3460__A1 _5560_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_hold429_A _6242_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_45_wb_clk_i_A clkbuf_leaf_6_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_30_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6486__A _6487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3622__B _5956_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5673__C1 _5673_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5743__A3 _3580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4530_ hold443/X _6273_/Q _4539_/S vssd1 vssd1 vccd1 vccd1 _4530_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_4_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold306 _6430_/Q vssd1 vssd1 vccd1 vccd1 hold306/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold317 _4608_/X vssd1 vssd1 vccd1 vccd1 _6249_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4461_ _4405_/X hold266/X _4464_/S vssd1 vssd1 vccd1 vccd1 _6164_/D sky130_fd_sc_hd__mux2_1
X_6200_ _6204_/CLK hold38/X fanout174/X vssd1 vssd1 vccd1 vccd1 hold37/A sky130_fd_sc_hd__dfrtp_1
Xhold328 _6261_/Q vssd1 vssd1 vccd1 vccd1 hold328/X sky130_fd_sc_hd__dlygate4sd3_1
X_3412_ _3573_/B _5480_/D vssd1 vssd1 vccd1 vccd1 _4260_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_7_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold339 _4822_/X vssd1 vssd1 vccd1 vccd1 _6277_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5051__S1 _5052_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4392_ _4427_/S _4388_/X _4390_/X _4391_/X vssd1 vssd1 vccd1 vccd1 _4392_/X sky130_fd_sc_hd__a22o_2
XFILLER_0_21_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6131_ _6410_/CLK _6131_/D vssd1 vssd1 vccd1 vccd1 _6131_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3343_ _5265_/A _5325_/A vssd1 vssd1 vccd1 vccd1 _3343_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_0_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3274_ _3426_/A _4520_/B _5291_/B _3274_/D vssd1 vssd1 vccd1 vccd1 _3280_/A sky130_fd_sc_hd__or4_1
XANTENNA__6437__SET_B fanout171/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6062_ hold594/X _5994_/Y _6061_/X _4313_/C vssd1 vssd1 vccd1 vccd1 _6062_/X sky130_fd_sc_hd__o22a_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5013_ _6113_/Q _6104_/Q _6096_/Q _6141_/Q _5358_/A0 _4326_/B vssd1 vssd1 vccd1 vccd1
+ _5013_/X sky130_fd_sc_hd__mux4_1
XANTENNA__3251__C _4679_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout167_A fanout168/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5915_ _5915_/A _5915_/B vssd1 vssd1 vccd1 vccd1 _5917_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_91_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5719__A0 _6270_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5846_ _5846_/A _5846_/B vssd1 vssd1 vccd1 vccd1 _5848_/B sky130_fd_sc_hd__or2_1
XFILLER_0_75_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5195__A1 _6296_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5195__B2 _5371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5777_ _5236_/S _6419_/Q _3580_/A _5735_/X vssd1 vssd1 vccd1 vccd1 _5779_/B sky130_fd_sc_hd__o31a_1
XFILLER_0_90_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4728_ _6274_/Q _4680_/X _5075_/B hold445/X vssd1 vssd1 vccd1 vccd1 _4728_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_71_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4659_ _6336_/Q _6340_/Q _4674_/S vssd1 vssd1 vccd1 vccd1 _4659_/X sky130_fd_sc_hd__mux2_1
X_6329_ _6383_/CLK _6329_/D fanout168/X vssd1 vssd1 vccd1 vccd1 _6329_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_98_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3681__A1 _3611_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5369__B _6427_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4630__B1 _4617_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5186__A1 _3573_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_1_wb_clk_i_A clkbuf_leaf_6_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_10_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3633__A _5715_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5646__C1 _5675_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3672__A1 _3482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_29_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6326_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_58_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3961_ _3723_/X _6040_/A _4391_/A2 vssd1 vssd1 vccd1 vccd1 _3961_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_97_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5700_ hold23/X _3841_/Y _6060_/S vssd1 vssd1 vccd1 vccd1 hold24/A sky130_fd_sc_hd__mux2_1
X_3892_ _5087_/A _6243_/Q _6337_/Q _3740_/Y _3891_/X vssd1 vssd1 vccd1 vccd1 _5111_/B
+ sky130_fd_sc_hd__o41a_1
XFILLER_0_85_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5631_ _5631_/A _5631_/B vssd1 vssd1 vccd1 vccd1 _5631_/X sky130_fd_sc_hd__or2_1
X_5562_ _5323_/C _4208_/B _5315_/A vssd1 vssd1 vccd1 vccd1 _5562_/X sky130_fd_sc_hd__a21o_1
XANTENNA__4385__C1 _5673_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4513_ _3965_/X hold288/X _4518_/S vssd1 vssd1 vccd1 vccd1 _6217_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_13_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold114 _5285_/X vssd1 vssd1 vccd1 vccd1 _6300_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold125 _4502_/X vssd1 vssd1 vccd1 vccd1 _6207_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold103 _6220_/Q vssd1 vssd1 vccd1 vccd1 hold103/X sky130_fd_sc_hd__dlygate4sd3_1
X_5493_ _6057_/A _5377_/X hold383/X vssd1 vssd1 vccd1 vccd1 _5493_/Y sky130_fd_sc_hd__o21ai_1
Xhold147 _6097_/Q vssd1 vssd1 vccd1 vccd1 hold147/X sky130_fd_sc_hd__dlygate4sd3_1
X_4444_ hold49/X _4412_/X _4446_/S vssd1 vssd1 vccd1 vccd1 hold50/A sky130_fd_sc_hd__mux2_1
Xhold158 _5724_/X vssd1 vssd1 vccd1 vccd1 _6368_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold136 _6150_/Q vssd1 vssd1 vccd1 vccd1 hold136/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4639__A _4679_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4375_ _5690_/S _4372_/X _4373_/X _4374_/X vssd1 vssd1 vccd1 vccd1 _4375_/X sky130_fd_sc_hd__o31a_1
XANTENNA__5234__S _5447_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold169 _6098_/Q vssd1 vssd1 vccd1 vccd1 hold169/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4152__A2 _3779_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3326_ _3525_/B _3334_/C _3525_/A vssd1 vssd1 vccd1 vccd1 _4081_/S sky130_fd_sc_hd__and3b_2
XANTENNA__3543__A _4541_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6114_ _6194_/CLK _6114_/D vssd1 vssd1 vccd1 vccd1 hold99/A sky130_fd_sc_hd__dfxtp_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3262__B _5578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5637__C1 _5673_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6045_ _3046_/A _6043_/X _6044_/Y hold411/X _6029_/Y vssd1 vssd1 vccd1 vccd1 _6045_/X
+ sky130_fd_sc_hd__o32a_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3257_ _3403_/B _3501_/B _3546_/B _3632_/B vssd1 vssd1 vccd1 vccd1 _3257_/X sky130_fd_sc_hd__and4b_1
XANTENNA__4691__A1_N _6268_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3188_ _5733_/A _3386_/A _3520_/A _3686_/C vssd1 vssd1 vccd1 vccd1 _3189_/C sky130_fd_sc_hd__or4_1
XFILLER_0_88_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5168__A1 _6040_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5829_ _5836_/B _5823_/X _5828_/X _5932_/S vssd1 vssd1 vccd1 vccd1 _5829_/X sky130_fd_sc_hd__a2bb2o_1
XANTENNA__3718__A _6313_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold496_A _6336_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold670 _6118_/Q vssd1 vssd1 vccd1 vccd1 hold670/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold681 _6307_/Q vssd1 vssd1 vccd1 vccd1 hold681/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_hold663_A _6318_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4284__A _4284_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3628__A _5560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5331__A1 _5317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4160_ _5217_/A _4160_/B vssd1 vssd1 vccd1 vccd1 _4163_/A sky130_fd_sc_hd__xor2_1
XANTENNA__3342__B1 _3309_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3111_ _4744_/A _3293_/B _6254_/Q vssd1 vssd1 vccd1 vccd1 _3116_/A sky130_fd_sc_hd__or3_4
XANTENNA__3893__A1 _6341_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5095__A0 _4070_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4091_ _6096_/Q _3789_/X _3791_/X _6197_/Q vssd1 vssd1 vccd1 vccd1 _4091_/X sky130_fd_sc_hd__a22o_1
X_3042_ _6389_/Q vssd1 vssd1 vccd1 vccd1 _5574_/A sky130_fd_sc_hd__clkinv_4
XANTENNA__5634__A2 _4382_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4993_ _6112_/Q hold77/A _6095_/Q _6140_/Q _5051_/S0 _4326_/B vssd1 vssd1 vccd1 vccd1
+ _4993_/X sky130_fd_sc_hd__mux4_1
X_3944_ _3740_/Y _3942_/X _3943_/X vssd1 vssd1 vccd1 vccd1 _3944_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_85_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3875_ _3877_/B _3877_/C _3877_/A vssd1 vssd1 vccd1 vccd1 _3878_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_73_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5614_ _6092_/Q _4198_/B _5676_/B1 _6137_/Q _5676_/C1 vssd1 vssd1 vccd1 vccd1 _5615_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_26_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4373__A2 _4382_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5545_ _5533_/B _5535_/B _5531_/X vssd1 vssd1 vccd1 vccd1 _5546_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_41_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5476_ _5554_/A _5476_/B vssd1 vssd1 vccd1 vccd1 _5477_/B sky130_fd_sc_hd__nor2_1
XANTENNA__4125__A2 _6248_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3402__A_N _4679_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4427_ _4425_/X _4426_/X _4427_/S vssd1 vssd1 vccd1 vccd1 _4427_/X sky130_fd_sc_hd__mux2_2
X_4358_ hold246/X _4102_/X _4360_/S vssd1 vssd1 vccd1 vccd1 _6113_/D sky130_fd_sc_hd__mux2_1
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5899__S _5933_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3309_ _5574_/A _4558_/A _4541_/A vssd1 vssd1 vccd1 vccd1 _3309_/Y sky130_fd_sc_hd__a21oi_4
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4289_ _4287_/A _4288_/X _6064_/S vssd1 vssd1 vccd1 vccd1 _4289_/X sky130_fd_sc_hd__mux2_1
X_6028_ _6028_/A _6028_/B vssd1 vssd1 vccd1 vccd1 _6063_/S sky130_fd_sc_hd__or2_4
XANTENNA__5625__A2 _4198_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4833__B1 _4867_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5312__A1_N _3502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5389__A1 input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout64 _5833_/B vssd1 vssd1 vccd1 vccd1 _5926_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_91_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout97 _3475_/X vssd1 vssd1 vccd1 vccd1 _5740_/A sky130_fd_sc_hd__clkbuf_8
Xfanout86 _3684_/X vssd1 vssd1 vccd1 vccd1 _4382_/C sky130_fd_sc_hd__buf_4
Xfanout75 _3718_/Y vssd1 vssd1 vccd1 vccd1 _5676_/B1 sky130_fd_sc_hd__buf_4
XFILLER_0_36_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3167__B _3656_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5010__A0 _6420_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3630__B _6404_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3722__S1 _5676_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5049__S _5557_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3660_ _3510_/B _3654_/A _5728_/B _3309_/Y _3386_/A vssd1 vssd1 vccd1 vccd1 _5563_/A
+ sky130_fd_sc_hd__a32o_2
XFILLER_0_82_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3591_ _5322_/B _3591_/B _5481_/A _5077_/B vssd1 vssd1 vccd1 vccd1 _3592_/B sky130_fd_sc_hd__or4_1
XFILLER_0_23_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5330_ _4214_/A _5329_/X _5330_/S vssd1 vssd1 vccd1 vccd1 _5330_/X sky130_fd_sc_hd__mux2_1
X_5261_ _5258_/B _5256_/A _5260_/Y vssd1 vssd1 vccd1 vccd1 _5261_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__5304__A1 _3482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4107__A2 _3715_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4212_ _4207_/X _4209_/Y _5343_/A _4228_/A vssd1 vssd1 vccd1 vccd1 _4212_/X sky130_fd_sc_hd__o31a_1
XFILLER_0_11_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5192_ _3075_/Y _6296_/Q _5192_/S vssd1 vssd1 vccd1 vccd1 _5192_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_44_wb_clk_i clkbuf_leaf_6_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6355_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_76_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4143_ _6022_/A vssd1 vssd1 vccd1 vccd1 _4143_/Y sky130_fd_sc_hd__inv_2
X_4074_ _6247_/Q _4075_/B vssd1 vssd1 vccd1 vccd1 _4174_/C sky130_fd_sc_hd__or2_1
XANTENNA__4636__B _4636_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3618__A1 _4214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5240__A0 hold560/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4976_ _5054_/A _4976_/B vssd1 vssd1 vccd1 vccd1 _4976_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__3268__A _4255_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3927_ _6093_/Q _3789_/X _3791_/X _6194_/Q vssd1 vssd1 vccd1 vccd1 _3927_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_6_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3858_ _3862_/S _3857_/X _3850_/A vssd1 vssd1 vccd1 vccd1 _3858_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_61_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3789_ _3850_/A _3862_/S _3861_/S vssd1 vssd1 vccd1 vccd1 _3789_/X sky130_fd_sc_hd__and3_4
X_5528_ _6420_/Q _5558_/S _5527_/X vssd1 vssd1 vccd1 vccd1 _5528_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_14_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3715__B _3862_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5459_ _6422_/Q _5458_/Y _5471_/S vssd1 vssd1 vccd1 vccd1 _5459_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_10_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4562__A _5725_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5231__B1 _5242_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5393__A _6427_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5568__A _5935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4830_ _5058_/S _4830_/B vssd1 vssd1 vccd1 vccd1 _4830_/X sky130_fd_sc_hd__or2_1
XFILLER_0_28_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3088__A _5226_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4761_ _6371_/Q _6319_/Q _6315_/Q vssd1 vssd1 vccd1 vccd1 _4761_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_28_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3712_ _3473_/A _3697_/X _3674_/B _3365_/B vssd1 vssd1 vccd1 vccd1 _3712_/X sky130_fd_sc_hd__o211a_2
X_4692_ _6268_/Q _4681_/X _4691_/X _5029_/S vssd1 vssd1 vccd1 vccd1 _4692_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_43_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3643_ _5931_/S _5978_/A _5728_/C vssd1 vssd1 vccd1 vccd1 _3643_/X sky130_fd_sc_hd__or3b_1
X_6431_ _6432_/CLK _6431_/D fanout178/X vssd1 vssd1 vccd1 vccd1 _6431_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__5525__B2 _5377_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6362_ _6376_/CLK _6362_/D fanout167/X vssd1 vssd1 vccd1 vccd1 _6362_/Q sky130_fd_sc_hd__dfrtp_2
X_5313_ _5313_/A _5313_/B vssd1 vssd1 vccd1 vccd1 _5313_/X sky130_fd_sc_hd__and2_1
XANTENNA__3535__B _6256_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3574_ _5096_/A _3574_/B vssd1 vssd1 vccd1 vccd1 _3574_/Y sky130_fd_sc_hd__nand2_1
X_6293_ _6423_/CLK _6293_/D fanout175/X vssd1 vssd1 vccd1 vccd1 _6293_/Q sky130_fd_sc_hd__dfstp_4
X_5244_ hold617/X _5243_/X _5347_/A vssd1 vssd1 vccd1 vccd1 _5244_/X sky130_fd_sc_hd__mux2_1
X_5175_ _6339_/Q _3502_/A _4188_/C _3985_/X vssd1 vssd1 vccd1 vccd1 _5175_/X sky130_fd_sc_hd__a31o_1
Xhold18 hold18/A vssd1 vssd1 vccd1 vccd1 hold18/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 hold29/A vssd1 vssd1 vccd1 vccd1 hold29/X sky130_fd_sc_hd__dlygate4sd3_1
X_4126_ _6248_/Q _4171_/S vssd1 vssd1 vccd1 vccd1 _4128_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__3551__A _5096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5242__S _5242_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4057_ _5088_/B _6341_/Q vssd1 vssd1 vccd1 vccd1 _4058_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5213__B1 _5560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4959_ _6269_/Q _4758_/X _4958_/B _4757_/Y vssd1 vssd1 vccd1 vccd1 _4959_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5764__A1 _5236_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5516__A1 _6419_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3445__B _3473_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_35_wb_clk_i_A clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_14_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xci2406_z80_208 vssd1 vssd1 vccd1 vccd1 ci2406_z80_208/HI io_out[31] sky130_fd_sc_hd__conb_1
XANTENNA__4991__S _5557_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5678__S1 _5690_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4007__B2 _4427_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4191__A0 _6423_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3290_ _3293_/B _3290_/B _3289_/C vssd1 vssd1 vccd1 vccd1 _3418_/A sky130_fd_sc_hd__or3b_2
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5443__B1 _5371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5931_ _5930_/X _5925_/A _5931_/S vssd1 vssd1 vccd1 vccd1 _5931_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4633__C _4633_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4406__S _4428_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5862_ _6417_/Q _5861_/X _5930_/S vssd1 vssd1 vccd1 vccd1 _5862_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4549__A2 _5578_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5793_ _5813_/A _5793_/B vssd1 vssd1 vccd1 vccd1 _5793_/X sky130_fd_sc_hd__or2_1
X_4813_ _6418_/Q _4758_/X _4811_/X _5061_/A1 vssd1 vssd1 vccd1 vccd1 _4813_/X sky130_fd_sc_hd__a22o_1
X_4744_ _4744_/A _4744_/B _6258_/Q vssd1 vssd1 vccd1 vccd1 _4744_/X sky130_fd_sc_hd__and3_1
XFILLER_0_16_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3546__A _4224_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4675_ _4674_/X _6245_/Q _4675_/S vssd1 vssd1 vccd1 vccd1 _4675_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_71_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3626_ _6415_/Q _4287_/B _3639_/C _3047_/Y vssd1 vssd1 vccd1 vccd1 _3626_/X sky130_fd_sc_hd__o211a_1
X_6414_ _6414_/CLK _6414_/D vssd1 vssd1 vccd1 vccd1 _6414_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3557_ _3116_/C _3556_/X _5256_/A vssd1 vssd1 vccd1 vccd1 _3557_/Y sky130_fd_sc_hd__o21ai_1
X_6345_ _6351_/CLK _6345_/D vssd1 vssd1 vccd1 vccd1 _6345_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput19 _6485_/X vssd1 vssd1 vccd1 vccd1 io_oeb[26] sky130_fd_sc_hd__buf_12
X_6276_ _6368_/CLK _6276_/D fanout169/X vssd1 vssd1 vccd1 vccd1 _6276_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__5480__B _5733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3488_ _4541_/B _5975_/S vssd1 vssd1 vccd1 vccd1 _4287_/B sky130_fd_sc_hd__nor2_4
X_5227_ _5240_/S _5222_/X _5226_/X vssd1 vssd1 vccd1 vccd1 _5227_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_98_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5158_ _5158_/A _5158_/B vssd1 vssd1 vccd1 vccd1 _5158_/Y sky130_fd_sc_hd__nor2_1
X_5089_ _5150_/B _5182_/B _5089_/S vssd1 vssd1 vccd1 vccd1 _5089_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_79_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4109_ _4110_/B vssd1 vssd1 vccd1 vccd1 _4111_/B sky130_fd_sc_hd__inv_2
XANTENNA__5700__S _6060_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5985__B2 _5518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3460__A2 _3443_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3996__B1 _3781_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5737__A1 _4639_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3515__A3 _4734_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4734__B _4734_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5525__A2_N _5377_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5057__S _6315_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5284__C _5347_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold307 _5980_/X vssd1 vssd1 vccd1 vccd1 _6424_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4460_ _4399_/X hold285/X _4464_/S vssd1 vssd1 vccd1 vccd1 _6163_/D sky130_fd_sc_hd__mux2_1
Xhold329 _4652_/X vssd1 vssd1 vccd1 vccd1 _6261_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3411_ _5158_/A _3224_/X _4268_/A vssd1 vssd1 vccd1 vccd1 _3414_/C sky130_fd_sc_hd__a21oi_1
Xhold318 hold680/X vssd1 vssd1 vccd1 vccd1 _4633_/B sky130_fd_sc_hd__buf_1
X_4391_ hold23/X _4391_/A2 _5597_/B vssd1 vssd1 vccd1 vccd1 _4391_/X sky130_fd_sc_hd__o21a_1
XANTENNA__5900__A1 _6384_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3342_ _3337_/A _3549_/B _3309_/Y _3427_/B _3341_/X vssd1 vssd1 vccd1 vccd1 _3342_/X
+ sky130_fd_sc_hd__o221a_1
X_6130_ _6209_/CLK hold46/X vssd1 vssd1 vccd1 vccd1 hold45/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__3911__B1 _3786_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3273_ _3591_/B _3373_/B _3273_/C vssd1 vssd1 vccd1 vccd1 _3274_/D sky130_fd_sc_hd__or3_1
X_6061_ _6057_/B _5054_/B _5555_/Y _5992_/Y vssd1 vssd1 vccd1 vccd1 _6061_/X sky130_fd_sc_hd__o22a_1
XANTENNA__4197__A _6314_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5012_ hold401/X _5011_/X _5068_/S vssd1 vssd1 vccd1 vccd1 _5012_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_30_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4219__A1 _3254_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5914_ _5914_/A _5926_/A vssd1 vssd1 vccd1 vccd1 _5915_/B sky130_fd_sc_hd__or2_1
XFILLER_0_48_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5845_ _5845_/A _5926_/A vssd1 vssd1 vccd1 vccd1 _5848_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_29_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5776_ _5765_/A _5742_/A _5775_/X _5731_/X vssd1 vssd1 vccd1 vccd1 _5776_/X sky130_fd_sc_hd__o22a_1
X_4727_ hold560/X hold157/X _4727_/S vssd1 vssd1 vccd1 vccd1 _4727_/X sky130_fd_sc_hd__mux2_1
X_4658_ _6048_/A _4673_/B vssd1 vssd1 vccd1 vccd1 _4658_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3609_ _3607_/X _3608_/Y _4309_/A vssd1 vssd1 vccd1 vccd1 _6127_/D sky130_fd_sc_hd__mux2_2
XFILLER_0_31_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4589_ _4020_/B _3826_/B _4604_/S vssd1 vssd1 vccd1 vccd1 _4589_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6334__RESET_B fanout168/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6328_ _6448_/CLK _6328_/D fanout168/X vssd1 vssd1 vccd1 vccd1 _6328_/Q sky130_fd_sc_hd__dfrtp_1
X_6259_ _6266_/CLK _6259_/D fanout177/X vssd1 vssd1 vccd1 vccd1 _6259_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__3681__A2 _5739_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold441_A _6244_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5186__A2 _5193_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4570__A _4604_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5591__C1 _5675_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6443__SET_B fanout171/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4146__B1 _5597_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5646__B1 _5676_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4745__A _5560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3672__A2 _5322_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3960_ _6040_/A vssd1 vssd1 vccd1 vccd1 _3960_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_85_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3891_ _3740_/Y _3889_/X _3890_/X vssd1 vssd1 vccd1 vccd1 _3891_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_72_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5630_ _6435_/Q _5588_/X _5610_/X _6443_/Q _5629_/X vssd1 vssd1 vccd1 vccd1 _5631_/B
+ sky130_fd_sc_hd__a221o_1
X_5561_ _5561_/A _5561_/B vssd1 vssd1 vccd1 vccd1 _5561_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__4385__B1 _3718_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4512_ _3923_/X hold209/X _4518_/S vssd1 vssd1 vccd1 vccd1 _6216_/D sky130_fd_sc_hd__mux2_1
X_5492_ _5492_/A _5492_/B vssd1 vssd1 vccd1 vccd1 _5492_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold126 _6109_/Q vssd1 vssd1 vccd1 vccd1 hold126/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold104 _4516_/X vssd1 vssd1 vccd1 vccd1 _6220_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold115 _6177_/Q vssd1 vssd1 vccd1 vccd1 hold115/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3695__C_N _4633_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold148 _4335_/X vssd1 vssd1 vccd1 vccd1 _6097_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4443_ hold61/X _4405_/X _4446_/S vssd1 vssd1 vccd1 vccd1 hold62/A sky130_fd_sc_hd__mux2_1
Xhold159 _6190_/Q vssd1 vssd1 vccd1 vccd1 hold159/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold137 _4445_/X vssd1 vssd1 vccd1 vccd1 _6150_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4639__B _4639_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4374_ _6314_/Q _4197_/B _5675_/C1 _4371_/X _4370_/X vssd1 vssd1 vccd1 vccd1 _4374_/X
+ sky130_fd_sc_hd__a221o_1
X_3325_ _3525_/A _4685_/A vssd1 vssd1 vccd1 vccd1 _3494_/B sky130_fd_sc_hd__nand2_1
XANTENNA__3543__B _4734_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6113_ _6331_/CLK _6113_/D vssd1 vssd1 vccd1 vccd1 _6113_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3256_ _3278_/A _5256_/A vssd1 vssd1 vccd1 vccd1 _3546_/B sky130_fd_sc_hd__or2_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6044_ _6044_/A _6063_/S vssd1 vssd1 vccd1 vccd1 _6044_/Y sky130_fd_sc_hd__nor2_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3187_ _3683_/B _3683_/C vssd1 vssd1 vccd1 vccd1 _3686_/C sky130_fd_sc_hd__and2_1
XFILLER_0_95_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5168__A2 _5243_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5828_ _5827_/X hold504/X _5931_/S vssd1 vssd1 vccd1 vccd1 _5828_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_29_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5759_ _5758_/X _6320_/Q _5825_/S vssd1 vssd1 vccd1 vccd1 _5760_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_8_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3718__B _4382_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold671 _6256_/Q vssd1 vssd1 vccd1 vccd1 hold671/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold660 _4620_/X vssd1 vssd1 vccd1 vccd1 _6252_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout92_A _5029_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold682 _6406_/Q vssd1 vssd1 vccd1 vccd1 hold682/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_hold656_A _6090_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4851__A1 _6420_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4284__B _4639_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4851__B2 _5061_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4603__A1 _5695_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3909__A _6036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4504__S _4509_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6256__RESET_B fanout179/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5331__A2 _5096_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3342__A1 _3337_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3110_ _3483_/A _3451_/C vssd1 vssd1 vccd1 vccd1 _3362_/B sky130_fd_sc_hd__or2_1
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4090_ _6220_/Q _3784_/X _3786_/X hold85/A _4089_/X vssd1 vssd1 vccd1 vccd1 _4093_/A
+ sky130_fd_sc_hd__a221o_1
X_3041_ _6297_/Q vssd1 vssd1 vccd1 vccd1 _3333_/S sky130_fd_sc_hd__inv_2
X_4992_ hold389/X _4991_/X _5068_/S vssd1 vssd1 vccd1 vccd1 _4992_/X sky130_fd_sc_hd__mux2_1
X_3943_ _5087_/B _3938_/X _3942_/A _3741_/X vssd1 vssd1 vccd1 vccd1 _3943_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_18_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3874_ _3805_/B _3811_/Y _3818_/Y _3826_/B _4111_/A vssd1 vssd1 vccd1 vccd1 _3877_/C
+ sky130_fd_sc_hd__o41ai_2
X_5613_ _6193_/Q _4198_/B _5676_/B1 _6069_/Q _5675_/C1 vssd1 vssd1 vccd1 vccd1 _5615_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_60_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5570__A2 _5603_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5544_ _5542_/X _5544_/B vssd1 vssd1 vccd1 vccd1 _5546_/A sky130_fd_sc_hd__nand2b_1
X_5475_ _5475_/A _5476_/B vssd1 vssd1 vccd1 vccd1 _5477_/A sky130_fd_sc_hd__and2_1
XFILLER_0_30_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4125__A3 _6342_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4426_ hold241/X hold65/X hold283/X hold71/X _5673_/C1 _4384_/S vssd1 vssd1 vccd1
+ vccd1 _4426_/X sky130_fd_sc_hd__mux4_1
XANTENNA__4369__B _4382_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4357_ hold120/X _4054_/X _4360_/S vssd1 vssd1 vccd1 vccd1 _4357_/X sky130_fd_sc_hd__mux2_1
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5086__A1 _5217_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3308_ _3611_/A _5158_/A vssd1 vssd1 vccd1 vccd1 _3308_/X sky130_fd_sc_hd__or2_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4288_ _6267_/Q _4287_/X _4305_/S vssd1 vssd1 vccd1 vccd1 _4288_/X sky130_fd_sc_hd__mux2_1
X_3239_ _3683_/C _3238_/C _3591_/B vssd1 vssd1 vccd1 vccd1 _3479_/B sky130_fd_sc_hd__a21o_1
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6027_ _3046_/A _6025_/X _6026_/Y hold536/X _5995_/Y vssd1 vssd1 vccd1 vccd1 _6027_/X
+ sky130_fd_sc_hd__o32a_1
XANTENNA__4833__A1 _6419_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6035__B1 _6063_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout65 _5475_/A vssd1 vssd1 vccd1 vccd1 _5554_/A sky130_fd_sc_hd__buf_4
Xfanout98 _4762_/S vssd1 vssd1 vccd1 vccd1 _5058_/S sky130_fd_sc_hd__clkbuf_8
Xfanout76 _3718_/Y vssd1 vssd1 vccd1 vccd1 _4200_/S sky130_fd_sc_hd__buf_4
XFILLER_0_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3183__B _3183_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold490 _6233_/Q vssd1 vssd1 vccd1 vccd1 hold490/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4279__B _5603_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6274__SET_B fanout169/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3590_ _4679_/D _3590_/B vssd1 vssd1 vccd1 vccd1 _5077_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_70_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5260_ _5294_/A _5294_/B _5294_/C vssd1 vssd1 vccd1 vccd1 _5260_/Y sky130_fd_sc_hd__nor3_1
XFILLER_0_50_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4211_ _4223_/B _4222_/B _4211_/C vssd1 vssd1 vccd1 vccd1 _5343_/A sky130_fd_sc_hd__and3_1
XANTENNA__3315__A1 _3573_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5191_ hold613/X _5190_/X _5347_/A vssd1 vssd1 vccd1 vccd1 _6295_/D sky130_fd_sc_hd__mux2_1
X_4142_ _3063_/Y _4141_/Y _4142_/S vssd1 vssd1 vccd1 vccd1 _6022_/A sky130_fd_sc_hd__mux2_4
X_4073_ _6246_/Q _4073_/B _4073_/C vssd1 vssd1 vccd1 vccd1 _4075_/B sky130_fd_sc_hd__or3_1
XFILLER_0_92_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_13_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6397_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_78_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4975_ _4974_/X _4973_/X _5053_/S vssd1 vssd1 vccd1 vccd1 _4976_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_25_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout142_A _3482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3926_ _6110_/Q _3779_/X _3781_/X hold63/A _3925_/X vssd1 vssd1 vccd1 vccd1 _3929_/A
+ sky130_fd_sc_hd__a221o_1
XANTENNA__6024__A2_N _6054_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3268__B _5258_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6107__RESET_B fanout177/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3857_ _6176_/Q _6407_/Q _3861_/S vssd1 vssd1 vccd1 vccd1 _3857_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_6_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4426__S0 _5673_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3788_ hold179/X _4510_/B _4465_/A hold233/X _3783_/X vssd1 vssd1 vccd1 vccd1 _3797_/A
+ sky130_fd_sc_hd__o221a_1
X_5527_ _6057_/A _5525_/X _5526_/Y _5558_/S vssd1 vssd1 vccd1 vccd1 _5527_/X sky130_fd_sc_hd__o211a_1
XANTENNA_clkbuf_leaf_25_wb_clk_i_A _6404_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3715__C _3838_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5458_ _5560_/D _5455_/X _5457_/Y vssd1 vssd1 vccd1 vccd1 _5458_/Y sky130_fd_sc_hd__o21ai_1
X_5389_ hold579/X input8/X _5469_/S vssd1 vssd1 vccd1 vccd1 _5389_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5703__S _6060_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4409_ _4424_/A _4409_/B vssd1 vssd1 vccd1 vccd1 _4409_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__4827__B _6322_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4562__B _4568_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold619_A _6274_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3459__A _5935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4990__A0 _6419_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5298__A1 _3482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output36_A _6290_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4753__A _6389_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5222__A1 _6297_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3088__B _3952_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4760_ _6433_/Q _4756_/Y _4759_/X vssd1 vssd1 vccd1 vccd1 _4760_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_83_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6200__RESET_B fanout174/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3711_ hold35/A _3700_/B _4197_/B vssd1 vssd1 vccd1 vccd1 _3711_/Y sky130_fd_sc_hd__o21ai_2
X_4691_ _6268_/Q _4680_/X _5075_/B hold453/X vssd1 vssd1 vccd1 vccd1 _4691_/X sky130_fd_sc_hd__a2bb2o_1
XANTENNA__4899__S _6085_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3642_ _5077_/A _4255_/B _3642_/C _4222_/B vssd1 vssd1 vccd1 vccd1 _5728_/C sky130_fd_sc_hd__and4_1
X_6430_ _6430_/CLK _6430_/D fanout172/X vssd1 vssd1 vccd1 vccd1 _6430_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3536__A1 _4224_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4733__B1 _3477_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6361_ _6376_/CLK _6361_/D fanout167/X vssd1 vssd1 vccd1 vccd1 _6361_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5312_ _3502_/A _5256_/Y _5311_/Y _5578_/A vssd1 vssd1 vccd1 vccd1 _5313_/B sky130_fd_sc_hd__a2bb2o_1
X_3573_ _3573_/A _3573_/B vssd1 vssd1 vccd1 vccd1 _3574_/B sky130_fd_sc_hd__nor2_1
XANTENNA__3535__C _3725_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6292_ _6295_/CLK _6292_/D fanout177/X vssd1 vssd1 vccd1 vccd1 _6292_/Q sky130_fd_sc_hd__dfstp_4
X_5243_ _4193_/Y _5242_/X _5243_/S vssd1 vssd1 vccd1 vccd1 _5243_/X sky130_fd_sc_hd__mux2_1
X_5174_ _3992_/A _5205_/B _5196_/S vssd1 vssd1 vccd1 vccd1 _5174_/X sky130_fd_sc_hd__mux2_1
Xhold19 hold19/A vssd1 vssd1 vccd1 vccd1 hold19/X sky130_fd_sc_hd__dlygate4sd3_1
X_4125_ _5087_/A _6248_/Q _6342_/Q _3740_/Y _4124_/X vssd1 vssd1 vccd1 vccd1 _5109_/A
+ sky130_fd_sc_hd__o41a_2
XANTENNA__3551__B _5578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4056_ _4056_/A _4158_/B vssd1 vssd1 vccd1 vccd1 _4056_/X sky130_fd_sc_hd__and2_1
XANTENNA__4663__A _6052_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5749__C1 _4319_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4382__B _4382_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4016__A2 _3715_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4958_ _5054_/A _4958_/B vssd1 vssd1 vccd1 vccd1 _4958_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_19_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5764__A2 _6418_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3775__A1 _4224_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3909_ _6036_/A vssd1 vssd1 vccd1 vccd1 _3909_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4889_ _6422_/Q _4758_/X _4885_/X _5061_/A1 vssd1 vssd1 vccd1 vccd1 _4889_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_34_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3527__B2 _5472_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5433__S _5472_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4557__B _5578_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_1__f_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xci2406_z80_209 vssd1 vssd1 vccd1 vccd1 ci2406_z80_209/HI io_out[35] sky130_fd_sc_hd__conb_1
XFILLER_0_97_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3189__A _4520_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3230__A3 _4679_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4512__S _4518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4715__B1 _5075_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3652__A _4309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5443__A1 _5441_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5930_ _6423_/Q _5929_/X _5930_/S vssd1 vssd1 vccd1 vccd1 _5930_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_87_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5861_ _5929_/A1 _5860_/X _4938_/Y vssd1 vssd1 vccd1 vccd1 _5861_/X sky130_fd_sc_hd__a21bo_1
X_5792_ _6375_/Q _5792_/B vssd1 vssd1 vccd1 vccd1 _5793_/B sky130_fd_sc_hd__nor2_1
X_4812_ _6435_/Q _5056_/A2 _4757_/Y _4807_/X _4754_/X vssd1 vssd1 vccd1 vccd1 _4812_/X
+ sky130_fd_sc_hd__a221o_1
X_4743_ _5324_/A _5324_/B _4743_/C _5326_/C vssd1 vssd1 vccd1 vccd1 _4745_/C sky130_fd_sc_hd__or4_1
XFILLER_0_56_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5518__S _5518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4674_ _6339_/Q _6343_/Q _4674_/S vssd1 vssd1 vccd1 vccd1 _4674_/X sky130_fd_sc_hd__mux2_1
X_6413_ _6413_/CLK _6413_/D vssd1 vssd1 vccd1 vccd1 _6413_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3625_ _3625_/A _3625_/B vssd1 vssd1 vccd1 vccd1 _3639_/C sky130_fd_sc_hd__nand2_2
XFILLER_0_3_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3556_ _3186_/B _4346_/B _4637_/B _3590_/B vssd1 vssd1 vccd1 vccd1 _3556_/X sky130_fd_sc_hd__o22a_1
XANTENNA__4182__A1 _5217_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6344_ _6344_/CLK _6344_/D vssd1 vssd1 vccd1 vccd1 _6344_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout105_A _4732_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4658__A _6048_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6275_ _6368_/CLK _6275_/D fanout166/X vssd1 vssd1 vccd1 vccd1 _6275_/Q sky130_fd_sc_hd__dfrtp_1
X_5226_ _5226_/A _6427_/Q _5226_/C _5226_/D vssd1 vssd1 vccd1 vccd1 _5226_/X sky130_fd_sc_hd__and4_1
X_3487_ _3485_/A _5354_/A _3484_/B vssd1 vssd1 vccd1 vccd1 _3487_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_0_51_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5682__A1 _6273_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5157_ _5102_/B _5156_/X _5242_/S vssd1 vssd1 vccd1 vccd1 _5157_/X sky130_fd_sc_hd__o21ba_1
X_5088_ _6303_/Q _5088_/B vssd1 vssd1 vccd1 vccd1 _5182_/B sky130_fd_sc_hd__nor2_1
X_4108_ _4108_/A _4108_/B vssd1 vssd1 vccd1 vccd1 _4110_/B sky130_fd_sc_hd__nor2_1
XANTENNA__4237__A2 _6118_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4039_ _4066_/A _3760_/B _4031_/B _4038_/Y vssd1 vssd1 vccd1 vccd1 _5110_/A sky130_fd_sc_hd__a31o_1
XFILLER_0_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4332__S _4336_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4568__A _5725_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3472__A _3473_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4287__B _4287_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4507__S _4509_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4750__B _4750_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold308 _6309_/Q vssd1 vssd1 vccd1 vccd1 _5988_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3410_ _4541_/B _4637_/B vssd1 vssd1 vccd1 vccd1 _3410_/Y sky130_fd_sc_hd__nand2_1
X_4390_ _3723_/X _4389_/X _3961_/Y vssd1 vssd1 vccd1 vccd1 _4390_/X sky130_fd_sc_hd__a21o_1
Xhold319 _6279_/Q vssd1 vssd1 vccd1 vccd1 hold319/X sky130_fd_sc_hd__dlygate4sd3_1
X_3341_ _3654_/A _5728_/B _3510_/B vssd1 vssd1 vccd1 vccd1 _3341_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_0_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3272_ _5303_/A _4257_/B vssd1 vssd1 vccd1 vccd1 _3273_/C sky130_fd_sc_hd__nor2_1
X_6060_ _6054_/A _6059_/X _6060_/S vssd1 vssd1 vccd1 vccd1 _6447_/D sky130_fd_sc_hd__mux2_1
XANTENNA__4197__B _4197_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5011_ _6364_/Q _5010_/X _5557_/S vssd1 vssd1 vccd1 vccd1 _5011_/X sky130_fd_sc_hd__mux2_1
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4219__A2 _6118_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5416__A1 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3978__A1 _6243_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5913_ _5914_/A _5926_/A vssd1 vssd1 vccd1 vccd1 _5915_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_48_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5844_ hold538/X _5843_/X _5933_/S vssd1 vssd1 vccd1 vccd1 _5844_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_8_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5775_ _5932_/S _5770_/X _5774_/X _5747_/A vssd1 vssd1 vccd1 vccd1 _5775_/X sky130_fd_sc_hd__o22a_1
X_4726_ hold647/X _4725_/X _5447_/S vssd1 vssd1 vccd1 vccd1 _6273_/D sky130_fd_sc_hd__mux2_1
X_4657_ _5715_/B _4653_/Y _4656_/X hold348/X _4635_/Y vssd1 vssd1 vccd1 vccd1 _4657_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_0_44_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3608_ _3577_/A _5956_/B _4616_/A vssd1 vssd1 vccd1 vccd1 _3608_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_101_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4588_ _5695_/A1 hold470/X _4546_/Y _4587_/X vssd1 vssd1 vccd1 vccd1 _4588_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_12_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6327_ _6448_/CLK _6327_/D fanout168/X vssd1 vssd1 vccd1 vccd1 _6327_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_101_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3539_ _3100_/B _3537_/B _3528_/Y _3538_/X _4616_/B vssd1 vssd1 vccd1 vccd1 _3539_/X
+ sky130_fd_sc_hd__a32o_1
X_6258_ _6403_/CLK _6258_/D fanout179/X vssd1 vssd1 vccd1 vccd1 _6258_/Q sky130_fd_sc_hd__dfrtp_4
X_5209_ _5209_/A _5209_/B _5123_/B vssd1 vssd1 vccd1 vccd1 _5210_/C sky130_fd_sc_hd__or3b_1
X_6189_ _6221_/CLK _6189_/D vssd1 vssd1 vccd1 vccd1 _6189_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6374__RESET_B fanout169/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5711__S _6064_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6303__RESET_B fanout179/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5407__A1 _4830_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5958__A2 _3639_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4091__B1 _3791_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4630__A2 _4615_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold601_A _6325_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3467__A _5935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5591__B1 _5676_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6018__A _6052_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4082__B1 _6341_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3890_ _5087_/B _3885_/X _3889_/A _3741_/X vssd1 vssd1 vccd1 vccd1 _3890_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_57_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5560_ _5560_/A _5560_/B _5560_/C _5560_/D vssd1 vssd1 vccd1 vccd1 _5561_/B sky130_fd_sc_hd__or4_1
XFILLER_0_5_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_38_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6386_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_4511_ _3881_/X hold179/X _4518_/S vssd1 vssd1 vccd1 vccd1 _4511_/X sky130_fd_sc_hd__mux2_1
X_5491_ _5478_/A _5478_/B _5477_/A vssd1 vssd1 vccd1 vccd1 _5492_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_26_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4137__A1 _4255_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold105 _6184_/Q vssd1 vssd1 vccd1 vccd1 hold105/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4442_ hold59/X _4399_/X _4446_/S vssd1 vssd1 vccd1 vccd1 hold60/A sky130_fd_sc_hd__mux2_1
XANTENNA__4700__S _5240_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold116 _4476_/X vssd1 vssd1 vccd1 vccd1 _6177_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold127 _4354_/X vssd1 vssd1 vccd1 vccd1 _6109_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4688__A2 _5240_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold149 _6159_/Q vssd1 vssd1 vccd1 vccd1 hold149/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 _6108_/Q vssd1 vssd1 vccd1 vccd1 hold138/X sky130_fd_sc_hd__dlygate4sd3_1
X_4373_ hold239/X _4382_/B _4384_/S hold115/X _5675_/C1 vssd1 vssd1 vccd1 vccd1 _4373_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_95_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3324_ _3525_/A _3334_/C _4070_/A _3525_/B vssd1 vssd1 vccd1 vccd1 _3324_/Y sky130_fd_sc_hd__nor4b_1
X_6112_ _6331_/CLK _6112_/D vssd1 vssd1 vccd1 vccd1 _6112_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3255_ _3278_/A _5256_/A vssd1 vssd1 vccd1 vccd1 _5359_/A sky130_fd_sc_hd__nor2_2
X_6043_ _6057_/A _6042_/X _6063_/S vssd1 vssd1 vccd1 vccd1 _6043_/X sky130_fd_sc_hd__o21a_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3186_ _4522_/D _3186_/B vssd1 vssd1 vccd1 vccd1 _3520_/A sky130_fd_sc_hd__nor2_1
XANTENNA_fanout172_A fanout173/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6062__B2 _4313_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3820__B1 _3786_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5827_ _6325_/Q _5826_/X _5852_/S vssd1 vssd1 vccd1 vccd1 _5827_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_29_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5758_ _6372_/Q _5849_/S _4783_/X vssd1 vssd1 vccd1 vccd1 _5758_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_44_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4709_ _6271_/Q _4680_/X _5075_/B hold476/X vssd1 vssd1 vccd1 vccd1 _4709_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_32_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5689_ _5689_/A _5689_/B vssd1 vssd1 vccd1 vccd1 _5689_/X sky130_fd_sc_hd__or2_1
XANTENNA__5706__S _6060_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold672 _4628_/X vssd1 vssd1 vccd1 vccd1 _6256_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold650 _6388_/Q vssd1 vssd1 vccd1 vccd1 hold650/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold661 _6315_/Q vssd1 vssd1 vccd1 vccd1 _3365_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold683 _6206_/Q vssd1 vssd1 vccd1 vccd1 hold683/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4846__A _6323_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_hold551_A _6425_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold649_A _6267_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4284__C _4284_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5800__A1 _6323_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4367__A1 _4382_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5616__S _5690_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5619__B2 _6417_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5619__A1 _6380_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3040_ _4767_/A vssd1 vssd1 vccd1 vccd1 _3040_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_65_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4991_ _6363_/Q _4990_/X _5557_/S vssd1 vssd1 vccd1 vccd1 _4991_/X sky130_fd_sc_hd__mux2_1
X_3942_ _3942_/A _3942_/B vssd1 vssd1 vccd1 vccd1 _3942_/X sky130_fd_sc_hd__xor2_1
XANTENNA__3802__B1 _3791_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3819__B _4594_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3873_ _4423_/A _4416_/A _4408_/A _4407_/B vssd1 vssd1 vccd1 vccd1 _3877_/B sky130_fd_sc_hd__or4_1
XFILLER_0_73_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5612_ _6434_/Q _5588_/X _5603_/X _6372_/Q _5611_/X vssd1 vssd1 vccd1 vccd1 _5620_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5543_ _5554_/A _5543_/B vssd1 vssd1 vccd1 vccd1 _5544_/B sky130_fd_sc_hd__or2_1
XANTENNA__3257__D _3632_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_15_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_5_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4430__S _4437_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5474_ _6441_/Q _4920_/B _5518_/S vssd1 vssd1 vccd1 vccd1 _5476_/B sky130_fd_sc_hd__mux2_1
X_4425_ hold7/X _4425_/A2 _4194_/Y _4424_/Y vssd1 vssd1 vccd1 vccd1 _4425_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_41_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4369__C _4382_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3964__S0 _5676_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4356_ hold163/X _4007_/X _4360_/S vssd1 vssd1 vccd1 vccd1 _4356_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4530__A1 _6273_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3307_ _5578_/A _5158_/A vssd1 vssd1 vccd1 vccd1 _3307_/Y sky130_fd_sc_hd__nor2_1
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4287_ _4287_/A _4287_/B vssd1 vssd1 vccd1 vccd1 _4287_/X sky130_fd_sc_hd__xor2_1
X_3238_ _3525_/B _4214_/B _3238_/C vssd1 vssd1 vccd1 vccd1 _3591_/B sky130_fd_sc_hd__and3_2
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6026_ _6026_/A _6026_/B vssd1 vssd1 vccd1 vccd1 _6026_/Y sky130_fd_sc_hd__nor2_1
X_3169_ _5303_/A _3369_/B vssd1 vssd1 vccd1 vccd1 _5328_/B sky130_fd_sc_hd__nor2_2
XANTENNA__6035__A1 _4313_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout55 _4916_/S vssd1 vssd1 vccd1 vccd1 _5068_/S sky130_fd_sc_hd__clkbuf_8
Xfanout88 _3642_/C vssd1 vssd1 vccd1 vccd1 _5258_/B sky130_fd_sc_hd__buf_4
Xfanout99 _4639_/B vssd1 vssd1 vccd1 vccd1 _5096_/B sky130_fd_sc_hd__buf_6
Xfanout77 _3718_/Y vssd1 vssd1 vccd1 vccd1 _4384_/S sky130_fd_sc_hd__buf_4
XFILLER_0_9_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout66 _5852_/S vssd1 vssd1 vccd1 vccd1 _5930_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_0_36_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4340__S _4345_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold599_A _6294_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5849__A1 _6379_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold480 _6236_/Q vssd1 vssd1 vccd1 vccd1 hold480/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold491 _4532_/X vssd1 vssd1 vccd1 vccd1 _6233_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5171__S _5193_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4588__A1 _5695_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4515__S _4518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6406__RESET_B fanout180/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4210_ _4210_/A _5258_/B vssd1 vssd1 vccd1 vccd1 _4211_/C sky130_fd_sc_hd__nand2_1
XANTENNA__3315__A2 _4214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5190_ _4049_/Y _5098_/A _5098_/Y _5189_/X vssd1 vssd1 vccd1 vccd1 _5190_/X sky130_fd_sc_hd__a22o_1
X_4141_ _5247_/A _6422_/Q _4140_/X vssd1 vssd1 vccd1 vccd1 _4141_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_48_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4072_ _4072_/A _4171_/S vssd1 vssd1 vccd1 vccd1 _4128_/A sky130_fd_sc_hd__or2_1
XANTENNA__4291__A3 _4287_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6017__A1 _6057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4974_ _6218_/Q _6155_/Q _6195_/Q _6071_/Q _5051_/S0 _5052_/S1 vssd1 vssd1 vccd1
+ vccd1 _4974_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_86_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3925_ _6217_/Q _3784_/X _3786_/X _6154_/Q vssd1 vssd1 vccd1 vccd1 _3925_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_6_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3856_ hold53/A hold95/A _3861_/S vssd1 vssd1 vccd1 vccd1 _3856_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_81_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3565__A _4637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3787_ _3850_/A _3862_/S _3861_/S vssd1 vssd1 vccd1 vccd1 _4465_/A sky130_fd_sc_hd__or3_1
X_5526_ _5526_/A _6057_/A vssd1 vssd1 vccd1 vccd1 _5526_/Y sky130_fd_sc_hd__nand2_1
X_5457_ _5560_/D _5457_/B vssd1 vssd1 vccd1 vccd1 _5457_/Y sky130_fd_sc_hd__nand2_1
X_4408_ _4408_/A _4408_/B vssd1 vssd1 vccd1 vccd1 _4409_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_41_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5388_ hold579/X _5377_/X _5387_/Y _5441_/A vssd1 vssd1 vccd1 vccd1 _5388_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_10_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3504__S _5472_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4339_ hold51/X _3923_/X _4345_/S vssd1 vssd1 vccd1 vccd1 hold52/A sky130_fd_sc_hd__mux2_1
XFILLER_0_5_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6009_ _5560_/D _6008_/X _5989_/X vssd1 vssd1 vccd1 vccd1 _6009_/X sky130_fd_sc_hd__o21a_1
XANTENNA__6008__B2 _4830_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4335__S _4336_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5298__A2 _5317_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4703__A1_N _6270_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4258__B1 _3309_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6026__A _6026_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3369__B _3369_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3710_ _3700_/C _3702_/X _3707_/X _3708_/Y vssd1 vssd1 vccd1 vccd1 _3862_/S sky130_fd_sc_hd__o31a_4
XFILLER_0_43_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4690_ _3072_/A _4689_/Y _4732_/S vssd1 vssd1 vccd1 vccd1 _6267_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_83_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3641_ _3641_/A _3641_/B _3641_/C vssd1 vssd1 vccd1 vccd1 _3641_/X sky130_fd_sc_hd__and3_1
XFILLER_0_55_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3536__A2 _3725_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3385__A _4541_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3572_ _3572_/A _3770_/A vssd1 vssd1 vccd1 vccd1 _3572_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_70_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5930__A0 _6423_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6360_ _6376_/CLK _6360_/D fanout166/X vssd1 vssd1 vccd1 vccd1 _6360_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__4733__A1 _5931_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5311_ _5258_/B _4222_/B _5260_/Y vssd1 vssd1 vccd1 vccd1 _5311_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_11_302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6291_ _6291_/CLK _6291_/D fanout177/X vssd1 vssd1 vccd1 vccd1 _6291_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_0_11_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5242_ _5241_/X _6423_/Q _5242_/S vssd1 vssd1 vccd1 vccd1 _5242_/X sky130_fd_sc_hd__mux2_1
X_5173_ _6294_/Q _5082_/X _5172_/X _5371_/A _5102_/B vssd1 vssd1 vccd1 vccd1 _5173_/X
+ sky130_fd_sc_hd__a221o_1
X_4124_ _3740_/Y _4121_/X _4123_/X vssd1 vssd1 vccd1 vccd1 _4124_/X sky130_fd_sc_hd__a21o_1
Xinput1 custom_settings[0] vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__clkbuf_4
X_4055_ _4054_/X hold224/X _4206_/S vssd1 vssd1 vccd1 vccd1 _4055_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4382__C _4382_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6399__RESET_B fanout174/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4957_ _4956_/X _4955_/X _5053_/S vssd1 vssd1 vccd1 vccd1 _4958_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_19_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5764__A3 _3580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3775__A2 _3770_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3908_ _4142_/S _3906_/X _3907_/X vssd1 vssd1 vccd1 vccd1 _6036_/A sky130_fd_sc_hd__a21oi_4
X_4888_ _6439_/Q _5056_/A2 _4757_/Y _4882_/B _4754_/X vssd1 vssd1 vccd1 vccd1 _4888_/X
+ sky130_fd_sc_hd__a221o_1
X_3839_ _3837_/X _3838_/X _3862_/S vssd1 vssd1 vccd1 vccd1 _3839_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6328__RESET_B fanout168/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5921__A0 _6422_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5509_ _6444_/Q _4976_/B _5518_/S vssd1 vssd1 vccd1 vccd1 _5510_/B sky130_fd_sc_hd__mux2_1
XANTENNA__5714__S _6064_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_hold631_A _6418_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5676__C1 _5676_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5860_ hold383/X _5928_/A2 _5928_/B1 _5859_/X vssd1 vssd1 vccd1 vccd1 _5860_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_87_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3099__B _5226_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4811_ _4807_/X _4810_/X _5058_/S vssd1 vssd1 vccd1 vccd1 _4811_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_56_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5595__A _6314_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4403__B1 _5597_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5791_ _5791_/A _5792_/B vssd1 vssd1 vccd1 vccd1 _5813_/A sky130_fd_sc_hd__and2_1
X_4742_ _5773_/A _5365_/C _5852_/S vssd1 vssd1 vccd1 vccd1 _4742_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4673_ _6026_/A _4673_/B vssd1 vssd1 vccd1 vccd1 _4673_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__3509__A2 _4734_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3624_ _4901_/S _5952_/B vssd1 vssd1 vccd1 vccd1 _3625_/B sky130_fd_sc_hd__and2_2
XANTENNA__5903__A0 _6421_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6412_ _6412_/CLK _6412_/D vssd1 vssd1 vccd1 vccd1 _6412_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3555_ _4224_/A _3595_/D _5360_/B vssd1 vssd1 vccd1 vccd1 _3555_/Y sky130_fd_sc_hd__o21ai_1
X_6343_ _6343_/CLK _6343_/D vssd1 vssd1 vccd1 vccd1 _6343_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_3_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3390__B1 _3611_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3486_ _3479_/B _3486_/B vssd1 vssd1 vccd1 vccd1 _5354_/A sky130_fd_sc_hd__and2b_1
X_6274_ _6374_/CLK _6274_/D fanout169/X vssd1 vssd1 vccd1 vccd1 _6274_/Q sky130_fd_sc_hd__dfstp_2
X_5225_ _5225_/A _5225_/B vssd1 vssd1 vccd1 vccd1 _5226_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5156_ hold588/X _5155_/X _5240_/S vssd1 vssd1 vccd1 vccd1 _5156_/X sky130_fd_sc_hd__mux2_1
X_5087_ _5087_/A _5087_/B vssd1 vssd1 vccd1 vccd1 _5150_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_79_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4107_ _6074_/Q _3715_/X _3794_/X _6142_/Q _4106_/X vssd1 vssd1 vccd1 vccd1 _4108_/B
+ sky130_fd_sc_hd__a221o_1
X_4038_ _3740_/Y _4034_/X _4059_/B _4037_/X vssd1 vssd1 vccd1 vccd1 _4038_/Y sky130_fd_sc_hd__a31oi_1
XFILLER_0_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3996__A2 _3779_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5198__B2 _6296_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5737__A3 _3770_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5989_ _5989_/A _5989_/B _6028_/B _4633_/C vssd1 vssd1 vccd1 vccd1 _5989_/X sky130_fd_sc_hd__or4b_1
XANTENNA__5709__S _6060_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3472__B _3473_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4568__B _4568_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5673__A2 _6313_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4397__C1 _5597_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5361__A1 _3611_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold309 _5338_/X vssd1 vssd1 vccd1 vccd1 _6309_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3340_ _4616_/A _6405_/Q vssd1 vssd1 vccd1 vccd1 _5728_/B sky130_fd_sc_hd__or2_4
XANTENNA__3911__A2 _3784_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5649__C1 _5675_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3271_ _3290_/B _3502_/A vssd1 vssd1 vccd1 vccd1 _3373_/B sky130_fd_sc_hd__nor2_1
X_5010_ _6420_/Q _5009_/X _5930_/S vssd1 vssd1 vccd1 vccd1 _5010_/X sky130_fd_sc_hd__mux2_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3675__A1 _5322_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4624__B1 _4617_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3978__A2 _6244_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5912_ _5905_/A _5742_/Y _5911_/X _5933_/S vssd1 vssd1 vccd1 vccd1 _5912_/X sky130_fd_sc_hd__a22o_1
X_5843_ _5837_/X _5842_/X _5932_/S vssd1 vssd1 vccd1 vccd1 _5843_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_33_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5529__S _6060_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4433__S _4437_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4927__B2 _4867_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4927__A1 _5061_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5774_ _4819_/Y _5773_/Y _6321_/Q _5852_/S vssd1 vssd1 vccd1 vccd1 _5774_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_71_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4725_ _4143_/Y _4724_/X _4731_/S vssd1 vssd1 vccd1 vccd1 _4725_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_16_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4656_ _3691_/B _4655_/X _4673_/B vssd1 vssd1 vccd1 vccd1 _4656_/X sky130_fd_sc_hd__o21a_1
X_3607_ _3606_/A _3652_/B _3645_/B vssd1 vssd1 vccd1 vccd1 _3607_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_3_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4587_ _4564_/A _4584_/X _4586_/X vssd1 vssd1 vccd1 vccd1 _4587_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_101_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3538_ _3536_/X _3537_/Y _3529_/Y vssd1 vssd1 vccd1 vccd1 _3538_/X sky130_fd_sc_hd__a21o_1
XANTENNA__3573__A _3573_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6326_ _6326_/CLK _6326_/D fanout175/X vssd1 vssd1 vccd1 vccd1 _6326_/Q sky130_fd_sc_hd__dfrtp_4
X_6257_ _6403_/CLK _6257_/D fanout179/X vssd1 vssd1 vccd1 vccd1 _6257_/Q sky130_fd_sc_hd__dfrtp_4
X_3469_ _3469_/A _5978_/A _3469_/C vssd1 vssd1 vccd1 vccd1 _3471_/C sky130_fd_sc_hd__nor3_1
X_5208_ _3333_/S _6312_/Q _5207_/X _6304_/Q vssd1 vssd1 vccd1 vccd1 _5208_/X sky130_fd_sc_hd__a211o_1
X_6188_ _6412_/CLK hold94/X vssd1 vssd1 vccd1 vccd1 hold93/A sky130_fd_sc_hd__dfxtp_1
X_5139_ _5216_/A _5216_/B vssd1 vssd1 vccd1 vccd1 _5140_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_98_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_8_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6433_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_94_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4343__S _4345_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3467__B _6392_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5646__A2 _4198_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4518__S _4518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6084__RESET_B fanout169/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4909__A1 _6423_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5582__B2 _3337_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4385__A2 _4382_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5490_ _5492_/A vssd1 vssd1 vccd1 vccd1 _5490_/Y sky130_fd_sc_hd__inv_2
X_4510_ _4510_/A _4510_/B vssd1 vssd1 vccd1 vccd1 _4518_/S sky130_fd_sc_hd__or2_4
XFILLER_0_41_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold117 _6398_/Q vssd1 vssd1 vccd1 vccd1 _3690_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold106 _4484_/X vssd1 vssd1 vccd1 vccd1 _6184_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4441_ hold55/X _4392_/X _4446_/S vssd1 vssd1 vccd1 vccd1 hold56/A sky130_fd_sc_hd__mux2_1
XFILLER_0_41_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold128 _6306_/Q vssd1 vssd1 vccd1 vccd1 hold128/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold139 _4353_/X vssd1 vssd1 vccd1 vccd1 _6108_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4372_ hold75/X _4382_/B _4384_/S hold57/X _5673_/C1 vssd1 vssd1 vccd1 vccd1 _4372_/X
+ sky130_fd_sc_hd__o221a_1
X_6111_ _6218_/CLK _6111_/D vssd1 vssd1 vccd1 vccd1 _6111_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3323_ _3334_/C _4070_/A _3525_/A _3525_/B vssd1 vssd1 vccd1 vccd1 _3323_/X sky130_fd_sc_hd__and4b_1
XANTENNA__4639__D _4767_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3254_ _3254_/A _3566_/A _5256_/A vssd1 vssd1 vccd1 vccd1 _3501_/B sky130_fd_sc_hd__or3_2
XANTENNA__5637__A2 _4382_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6042_ _5512_/Y _6054_/B _6057_/B _4976_/B vssd1 vssd1 vccd1 vccd1 _6042_/X sky130_fd_sc_hd__o2bb2a_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4428__S _4428_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3185_ _3206_/A _3238_/C vssd1 vssd1 vccd1 vccd1 _3427_/B sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_leaf_44_wb_clk_i_A clkbuf_leaf_6_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_91_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5022__A0 _6421_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5826_ _5773_/A _5825_/X _4882_/Y vssd1 vssd1 vccd1 vccd1 _5826_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_36_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5757_ _5757_/A _5757_/B vssd1 vssd1 vccd1 vccd1 _5769_/B sky130_fd_sc_hd__nor2_1
X_4708_ hold662/X _4707_/X _5447_/S vssd1 vssd1 vccd1 vccd1 _6270_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_32_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5688_ _6135_/Q _6313_/Q _4384_/S _6214_/Q _3720_/X vssd1 vssd1 vccd1 vccd1 _5689_/B
+ sky130_fd_sc_hd__o221a_1
X_4639_ _4679_/A _4639_/B _4639_/C _4767_/B vssd1 vssd1 vccd1 vccd1 _4675_/S sky130_fd_sc_hd__and4_4
Xhold651 _5942_/X vssd1 vssd1 vccd1 vccd1 _6388_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold640 _5944_/X vssd1 vssd1 vccd1 vccd1 _6389_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold662 _6270_/Q vssd1 vssd1 vccd1 vccd1 hold662/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold673 _6405_/Q vssd1 vssd1 vccd1 vccd1 hold673/X sky130_fd_sc_hd__dlygate4sd3_1
X_6309_ _6433_/CLK _6309_/D fanout173/X vssd1 vssd1 vccd1 vccd1 _6309_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__5722__S _5723_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4338__S _4345_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold544_A _6390_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5316__A1 _4541_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6265__RESET_B fanout177/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4990_ _6419_/Q _4989_/X _5930_/S vssd1 vssd1 vccd1 vccd1 _4990_/X sky130_fd_sc_hd__mux2_1
X_3941_ _3889_/A _3889_/B _3885_/B vssd1 vssd1 vccd1 vccd1 _3942_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_85_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3872_ _4408_/A _4407_/B vssd1 vssd1 vccd1 vccd1 _3872_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_73_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5611_ _6268_/Q _5589_/X _5610_/X _6442_/Q vssd1 vssd1 vccd1 vccd1 _5611_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5807__S _5931_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4711__S _4727_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5542_ _5554_/A _5543_/B vssd1 vssd1 vccd1 vccd1 _5542_/X sky130_fd_sc_hd__and2_1
XFILLER_0_26_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5307__A1 _5715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5473_ _5467_/A _5464_/Y _5466_/B vssd1 vssd1 vccd1 vccd1 _5478_/A sky130_fd_sc_hd__o21ai_2
X_4424_ _4424_/A _4424_/B vssd1 vssd1 vccd1 vccd1 _4424_/Y sky130_fd_sc_hd__nor2_1
X_4355_ hold109/X _3965_/X _4360_/S vssd1 vssd1 vccd1 vccd1 _4355_/X sky130_fd_sc_hd__mux2_1
X_3306_ _3359_/B _4756_/A vssd1 vssd1 vccd1 vccd1 _3361_/A sky130_fd_sc_hd__or2_1
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4286_ _5226_/A _5715_/A _4727_/S vssd1 vssd1 vccd1 vccd1 _4305_/S sky130_fd_sc_hd__or3b_4
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3237_ _3237_/A _3379_/B vssd1 vssd1 vccd1 vccd1 _4320_/B sky130_fd_sc_hd__nor2_2
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6025_ _6057_/A _6024_/X _6026_/B vssd1 vssd1 vccd1 vccd1 _6025_/X sky130_fd_sc_hd__o21a_1
X_3168_ _3293_/B _3232_/A vssd1 vssd1 vccd1 vccd1 _4679_/D sky130_fd_sc_hd__or2_4
XANTENNA_clkbuf_leaf_0_wb_clk_i_A clkbuf_leaf_6_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_3099_ _4284_/A _5226_/A _3952_/A vssd1 vssd1 vccd1 vccd1 _4255_/B sky130_fd_sc_hd__and3b_4
XFILLER_0_49_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5243__A0 _4193_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xci2406_z80_190 vssd1 vssd1 vccd1 vccd1 ci2406_z80_190/HI io_oeb[9] sky130_fd_sc_hd__conb_1
Xfanout56 _5977_/S vssd1 vssd1 vccd1 vccd1 _5931_/S sky130_fd_sc_hd__buf_8
XFILLER_0_9_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout78 _5773_/A vssd1 vssd1 vccd1 vccd1 _5929_/A1 sky130_fd_sc_hd__buf_4
X_5809_ _6376_/Q _5810_/B vssd1 vssd1 vccd1 vccd1 _5821_/A sky130_fd_sc_hd__and2_1
XFILLER_0_29_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout89 _5849_/S vssd1 vssd1 vccd1 vccd1 _5927_/S sky130_fd_sc_hd__clkbuf_8
Xfanout67 _4738_/Y vssd1 vssd1 vccd1 vccd1 _5852_/S sky130_fd_sc_hd__buf_4
XFILLER_0_91_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5717__S _5723_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4350__A1_N _4639_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold481 _4535_/X vssd1 vssd1 vccd1 vccd1 _6236_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold470 _6245_/Q vssd1 vssd1 vccd1 vccd1 hold470/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold661_A _6315_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold492 _6371_/Q vssd1 vssd1 vccd1 vccd1 _5745_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_35_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5785__A1 _6322_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3639__C _3639_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5537__B2 _5441_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5627__S _5690_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4140_ _3727_/X _5109_/A _4139_/X _6305_/Q vssd1 vssd1 vccd1 vccd1 _4140_/X sky130_fd_sc_hd__o211a_1
X_4071_ _6246_/Q _6247_/Q _4071_/C vssd1 vssd1 vccd1 vccd1 _4171_/S sky130_fd_sc_hd__and3_1
XFILLER_0_25_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4973_ _6111_/Q _6102_/Q _6094_/Q _6139_/Q _5051_/S0 _5052_/S1 vssd1 vssd1 vccd1
+ vccd1 _4973_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_86_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3924_ _3923_/X hold205/X _4206_/S vssd1 vssd1 vccd1 vccd1 _3924_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_73_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5528__A1 _6420_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4441__S _4446_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3855_ _3855_/A _3855_/B vssd1 vssd1 vccd1 vccd1 _5249_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_6_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout128_A _3337_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3786_ _3863_/A _3850_/B _3838_/S vssd1 vssd1 vccd1 vccd1 _3786_/X sky130_fd_sc_hd__and3_4
Xclkbuf_leaf_22_wb_clk_i _6404_/CLK vssd1 vssd1 vccd1 vccd1 _6266_/CLK sky130_fd_sc_hd__clkbuf_16
X_5525_ _6331_/Q _5377_/X _5524_/X _5377_/A vssd1 vssd1 vccd1 vccd1 _5525_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_14_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5456_ hold601/X input5/X _5469_/S vssd1 vssd1 vccd1 vccd1 _5457_/B sky130_fd_sc_hd__mux2_1
X_4407_ _3825_/X _4407_/B vssd1 vssd1 vccd1 vccd1 _4408_/B sky130_fd_sc_hd__and2b_1
XANTENNA__3711__B1 _4197_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5387_ _5387_/A vssd1 vssd1 vccd1 vccd1 _5387_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_10_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4338_ hold97/X _3881_/X _4345_/S vssd1 vssd1 vccd1 vccd1 hold98/A sky130_fd_sc_hd__mux2_1
X_4269_ _4685_/A _4541_/A _5578_/A vssd1 vssd1 vccd1 vccd1 _4269_/X sky130_fd_sc_hd__a21o_1
XANTENNA__4267__A1 _3573_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6008_ _5413_/B _6054_/B _4321_/A _4830_/B vssd1 vssd1 vccd1 vccd1 _6008_/X sky130_fd_sc_hd__o2bb2a_1
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4351__S _5347_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5447__S _5447_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4742__A2 _5365_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3950__A0 _6243_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3491__A _5313_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3640_ hold422/X _3683_/B _3629_/B hold588/X vssd1 vssd1 vccd1 vccd1 _3641_/C sky130_fd_sc_hd__a31o_1
XANTENNA__3536__A3 _5578_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3571_ _5265_/A _4346_/A _4268_/A vssd1 vssd1 vccd1 vccd1 _3571_/X sky130_fd_sc_hd__or3_1
XFILLER_0_70_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4733__A2 _5029_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5310_ _4221_/X _5321_/S _5309_/X hold616/X _5560_/B vssd1 vssd1 vccd1 vccd1 _6304_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_11_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6290_ _6290_/CLK _6290_/D fanout167/X vssd1 vssd1 vccd1 vccd1 _6290_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_87_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5241_ _5238_/X _5240_/X _5241_/S vssd1 vssd1 vccd1 vccd1 _5241_/X sky130_fd_sc_hd__mux2_1
X_5172_ _6236_/Q _5075_/B _5076_/Y _5171_/X vssd1 vssd1 vccd1 vccd1 _5172_/X sky130_fd_sc_hd__a22o_1
XANTENNA__6280__RESET_B fanout169/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4123_ _3741_/X _4121_/A _4122_/X _5087_/B vssd1 vssd1 vccd1 vccd1 _4123_/X sky130_fd_sc_hd__a22o_1
Xinput2 io_in[22] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4249__A1 _4255_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5446__A0 _6421_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4054_ _4051_/Y _4052_/X _4053_/X _4427_/S vssd1 vssd1 vccd1 vccd1 _4054_/X sky130_fd_sc_hd__a22o_2
XANTENNA__5997__A1 _5560_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4436__S _4437_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4956_ _6217_/Q _6154_/Q _6194_/Q _6070_/Q _5051_/S0 _5052_/S1 vssd1 vssd1 vccd1
+ vccd1 _4956_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_19_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3907_ _3907_/A _4158_/B vssd1 vssd1 vccd1 vccd1 _3907_/X sky130_fd_sc_hd__and2_1
XFILLER_0_46_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4887_ _6325_/Q _4866_/X _4886_/Y vssd1 vssd1 vccd1 vccd1 _4887_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_61_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3838_ _6409_/Q _6178_/Q _3838_/S vssd1 vssd1 vccd1 vccd1 _3838_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_34_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3769_ _4224_/A _5322_/D vssd1 vssd1 vccd1 vccd1 _3769_/X sky130_fd_sc_hd__and2_1
X_5508_ hold558/X _5507_/X _6060_/S vssd1 vssd1 vccd1 vccd1 _5508_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6368__RESET_B fanout169/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5439_ _5424_/B _5426_/B _5422_/X vssd1 vssd1 vccd1 vccd1 _5440_/B sky130_fd_sc_hd__a21o_1
XANTENNA_hold457_A _6341_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4660__A1 _6242_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3999__B1 _3794_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4412__A1 _4427_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5912__B2 _5933_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5676__B1 _5676_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5428__A0 _5226_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4100__B1 _5597_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3099__C _3952_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4810_ _6373_/Q _6321_/Q _6315_/Q vssd1 vssd1 vccd1 vccd1 _4810_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_68_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5790_ _5236_/S _6420_/Q _3580_/A _5735_/X vssd1 vssd1 vccd1 vccd1 _5792_/B sky130_fd_sc_hd__o31a_1
XFILLER_0_90_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5595__B _5597_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4741_ _4740_/X _4739_/X _5053_/S vssd1 vssd1 vccd1 vccd1 _5365_/C sky130_fd_sc_hd__mux2_4
XFILLER_0_16_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4672_ _5715_/B _4668_/Y _4671_/X hold334/X _4635_/Y vssd1 vssd1 vccd1 vccd1 _4672_/X
+ sky130_fd_sc_hd__o32a_1
X_3623_ _3623_/A vssd1 vssd1 vccd1 vccd1 _5952_/B sky130_fd_sc_hd__inv_2
X_6411_ _6412_/CLK _6411_/D vssd1 vssd1 vccd1 vccd1 _6411_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3914__B1 _3794_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5815__S _5815_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3554_ _5270_/A _5728_/B _3658_/B vssd1 vssd1 vccd1 vccd1 _3554_/X sky130_fd_sc_hd__a21bo_1
X_6342_ _6373_/CLK _6342_/D vssd1 vssd1 vccd1 vccd1 _6342_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__3335__S _6298_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3390__A1 _3770_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3485_ _3485_/A vssd1 vssd1 vccd1 vccd1 _5353_/A sky130_fd_sc_hd__inv_2
X_6273_ _6343_/CLK _6273_/D fanout170/X vssd1 vssd1 vccd1 vccd1 _6273_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_0_11_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5224_ _6361_/Q _6360_/Q _6363_/Q _6362_/Q vssd1 vssd1 vccd1 vccd1 _5225_/B sky130_fd_sc_hd__or4_1
X_5155_ _6235_/Q _6293_/Q _5239_/S vssd1 vssd1 vccd1 vccd1 _5155_/X sky130_fd_sc_hd__mux2_1
X_5086_ _5217_/A _4160_/B _4163_/Y vssd1 vssd1 vccd1 vccd1 _5089_/S sky130_fd_sc_hd__a21bo_1
X_4106_ _6097_/Q _3789_/X _3791_/X _6198_/Q vssd1 vssd1 vccd1 vccd1 _4106_/X sky130_fd_sc_hd__a22o_1
X_4037_ _3741_/X _4035_/A _4036_/Y _5087_/B vssd1 vssd1 vccd1 vccd1 _4037_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4642__A1 _5715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5988_ _5988_/A _5988_/B _5988_/C vssd1 vssd1 vccd1 vccd1 _6028_/B sky130_fd_sc_hd__or3_1
XFILLER_0_93_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4939_ _6268_/Q _4758_/X _4938_/B _4757_/Y vssd1 vssd1 vccd1 vccd1 _4939_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_19_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5460__S _5472_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4865__A _6324_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4076__S _6292_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3270_ _3683_/B _3683_/C _5560_/C vssd1 vssd1 vccd1 vccd1 _5291_/B sky130_fd_sc_hd__a21bo_1
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_34_wb_clk_i_A clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_5911_ _5909_/Y _5910_/X _5747_/Y _5903_/X vssd1 vssd1 vccd1 vccd1 _5911_/X sky130_fd_sc_hd__a2bb2o_1
XANTENNA__3978__A3 _6245_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5842_ _5841_/X hold538/X _5931_/S vssd1 vssd1 vccd1 vccd1 _5842_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_8_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4714__S _4732_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5773_ _5773_/A _5773_/B vssd1 vssd1 vccd1 vccd1 _5773_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_90_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4724_ _4721_/X _4723_/X _5240_/S vssd1 vssd1 vccd1 vccd1 _4724_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_44_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4655_ _4654_/X _6343_/Q _4675_/S vssd1 vssd1 vccd1 vccd1 _4655_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_44_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3606_ _3606_/A _3652_/B vssd1 vssd1 vccd1 vccd1 _3606_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_24_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4586_ hold455/X _4567_/Y _4568_/X hold411/X _4585_/X vssd1 vssd1 vccd1 vccd1 _4586_/X
+ sky130_fd_sc_hd__a221o_1
X_3537_ _3537_/A _3537_/B vssd1 vssd1 vccd1 vccd1 _3537_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__4560__B1 _5096_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6325_ _6326_/CLK _6325_/D fanout174/X vssd1 vssd1 vccd1 vccd1 _6325_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_12_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6256_ _6403_/CLK _6256_/D fanout179/X vssd1 vssd1 vccd1 vccd1 _6256_/Q sky130_fd_sc_hd__dfrtp_4
X_3468_ _4210_/A _6389_/Q _3545_/B _3467_/X _3459_/B vssd1 vssd1 vccd1 vccd1 _3469_/C
+ sky130_fd_sc_hd__o41a_1
X_5207_ _5109_/A _5109_/B _5206_/X _5347_/B vssd1 vssd1 vccd1 vccd1 _5207_/X sky130_fd_sc_hd__o31a_1
X_3399_ _5265_/A _3400_/B vssd1 vssd1 vccd1 vccd1 _3399_/X sky130_fd_sc_hd__or2_1
XANTENNA__4685__A _4685_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6187_ _6413_/CLK hold42/X vssd1 vssd1 vccd1 vccd1 hold41/A sky130_fd_sc_hd__dfxtp_1
X_5138_ _5216_/C _5216_/D vssd1 vssd1 vccd1 vccd1 _5140_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_98_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5069_ _5069_/A _5989_/B _4633_/C vssd1 vssd1 vccd1 vccd1 _6028_/A sky130_fd_sc_hd__or3b_1
XFILLER_0_79_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4091__A2 _3789_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5576__C1 _5317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4379__B1 _4382_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6383__RESET_B fanout168/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5591__A2 _4198_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6312__RESET_B fanout179/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4854__A1 _6323_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4440_ hold254/X _4380_/X _4446_/S vssd1 vssd1 vccd1 vccd1 _4440_/X sky130_fd_sc_hd__mux2_1
Xhold107 _6102_/Q vssd1 vssd1 vccd1 vccd1 hold107/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold118 _6088_/Q vssd1 vssd1 vccd1 vccd1 hold118/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold129 _5321_/X vssd1 vssd1 vccd1 vccd1 _6306_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4371_ hold67/X hold167/X _4384_/S vssd1 vssd1 vccd1 vccd1 _4371_/X sky130_fd_sc_hd__mux2_1
X_6110_ _6218_/CLK _6110_/D vssd1 vssd1 vccd1 vccd1 _6110_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_95_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3322_ _3334_/C _3537_/A vssd1 vssd1 vccd1 vccd1 _3988_/B sky130_fd_sc_hd__nor2_1
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3253_ _3253_/A _4639_/C vssd1 vssd1 vccd1 vccd1 _3403_/B sky130_fd_sc_hd__or2_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6041_ _3046_/A _6039_/X _6040_/Y hold554/X _6029_/Y vssd1 vssd1 vccd1 vccd1 _6041_/X
+ sky130_fd_sc_hd__o32a_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3184_ _4214_/B _3216_/A _3238_/C vssd1 vssd1 vccd1 vccd1 _3386_/A sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_47_wb_clk_i clkbuf_leaf_6_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6218_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6047__B1 _6063_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4444__S _4446_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3820__A2 _3784_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5825_ _5824_/X _6325_/Q _5825_/S vssd1 vssd1 vccd1 vccd1 _5825_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5573__A2 _4222_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5756_ _5757_/A _5757_/B vssd1 vssd1 vccd1 vccd1 _5756_/X sky130_fd_sc_hd__and2_1
X_4707_ _3994_/Y _4706_/X _4731_/S vssd1 vssd1 vccd1 vccd1 _4707_/X sky130_fd_sc_hd__mux2_1
X_5687_ _6414_/Q _6313_/Q _4384_/S _6183_/Q _3721_/Y vssd1 vssd1 vccd1 vccd1 _5689_/A
+ sky130_fd_sc_hd__o221a_1
X_4638_ _6242_/Q _6336_/Q _4674_/S vssd1 vssd1 vccd1 vccd1 _4638_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_32_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold630 _6085_/Q vssd1 vssd1 vccd1 vccd1 hold630/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold641 _6419_/Q vssd1 vssd1 vccd1 vccd1 hold641/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold652 _6297_/Q vssd1 vssd1 vccd1 vccd1 hold652/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold663 _6318_/Q vssd1 vssd1 vccd1 vccd1 hold663/X sky130_fd_sc_hd__dlygate4sd3_1
X_4569_ _4604_/S _4570_/B vssd1 vssd1 vccd1 vccd1 _4569_/X sky130_fd_sc_hd__and2b_2
Xhold674 _6253_/Q vssd1 vssd1 vccd1 vccd1 hold674/X sky130_fd_sc_hd__dlygate4sd3_1
X_6308_ _6428_/CLK _6308_/D fanout173/X vssd1 vssd1 vccd1 vccd1 _6308_/Q sky130_fd_sc_hd__dfrtp_1
X_6239_ _6297_/CLK _6239_/D fanout176/X vssd1 vssd1 vccd1 vccd1 _6239_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA__3750__C _6304_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4836__A1 _6322_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5261__A1 _5258_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4354__S _4360_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3494__A _6297_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3940_ _3938_/B _3940_/B vssd1 vssd1 vccd1 vccd1 _3942_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_98_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5587__C _5691_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3802__A2 _3789_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5004__A1 _6420_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3871_ _3870_/A _3870_/B _3870_/C _4401_/A vssd1 vssd1 vccd1 vccd1 _4407_/B sky130_fd_sc_hd__a31o_1
X_5610_ _5610_/A _5610_/B vssd1 vssd1 vccd1 vccd1 _5610_/X sky130_fd_sc_hd__and2_2
XFILLER_0_60_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5541_ _6447_/Q _6057_/C _5553_/S vssd1 vssd1 vccd1 vccd1 _5543_/B sky130_fd_sc_hd__mux2_1
XANTENNA__5095__S _5447_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5472_ hold590/X _5471_/X _5472_/S vssd1 vssd1 vccd1 vccd1 _5472_/X sky130_fd_sc_hd__mux2_1
X_4423_ _4423_/A _4423_/B vssd1 vssd1 vccd1 vccd1 _4424_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_41_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4354_ hold126/X _3923_/X _4360_/S vssd1 vssd1 vccd1 vccd1 _4354_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4439__S _4446_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3305_ _4756_/A vssd1 vssd1 vccd1 vccd1 _4758_/B sky130_fd_sc_hd__inv_2
X_4285_ _4685_/A _5553_/S _4727_/S vssd1 vssd1 vccd1 vccd1 _4316_/B sky130_fd_sc_hd__and3_2
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6024_ _5467_/Y _6054_/B _6057_/B _4900_/B vssd1 vssd1 vccd1 vccd1 _6024_/X sky130_fd_sc_hd__o2bb2a_1
X_3236_ _3230_/X _3231_/Y _3235_/X vssd1 vssd1 vccd1 vccd1 _5294_/B sky130_fd_sc_hd__o21ai_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3167_ _3482_/A _3656_/A vssd1 vssd1 vccd1 vccd1 _5578_/B sky130_fd_sc_hd__nand2_4
X_3098_ _3573_/A _3525_/B vssd1 vssd1 vccd1 vccd1 _3952_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_89_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3579__A _4734_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xci2406_z80_191 vssd1 vssd1 vccd1 vccd1 ci2406_z80_191/HI io_oeb[10] sky130_fd_sc_hd__conb_1
XFILLER_0_36_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout57 _3361_/X vssd1 vssd1 vccd1 vccd1 _5061_/A1 sky130_fd_sc_hd__clkbuf_8
Xfanout79 _4321_/B vssd1 vssd1 vccd1 vccd1 _5773_/A sky130_fd_sc_hd__buf_4
XANTENNA__4902__S _5058_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5808_ _5236_/S _6421_/Q _3580_/A _5735_/X vssd1 vssd1 vccd1 vccd1 _5810_/B sky130_fd_sc_hd__o31a_1
Xfanout68 _4156_/A vssd1 vssd1 vccd1 vccd1 _4111_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_91_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5739_ _5739_/A _5739_/B vssd1 vssd1 vccd1 vccd1 _5746_/B sky130_fd_sc_hd__and2_1
XFILLER_0_17_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3745__C _6304_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold460 _4538_/X vssd1 vssd1 vccd1 vccd1 _6239_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold471 _4588_/X vssd1 vssd1 vccd1 vccd1 _6245_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout90_A _5784_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold482 _6237_/Q vssd1 vssd1 vccd1 vccd1 hold482/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold493 _5752_/X vssd1 vssd1 vccd1 vccd1 _6371_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5034__A _5054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3489__A _3611_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5785__A2 _5772_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5537__A2 _5377_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3936__B _6338_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3952__A _3952_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4767__B _4767_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4070_ _4070_/A _5126_/B vssd1 vssd1 vccd1 vccd1 _4172_/C sky130_fd_sc_hd__or2_2
XFILLER_0_78_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4972_ hold363/X _4971_/X _5068_/S vssd1 vssd1 vccd1 vccd1 _4972_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_25_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4984__A0 _6419_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3923_ _3920_/X _3921_/X _3922_/X _4427_/S vssd1 vssd1 vccd1 vccd1 _3923_/X sky130_fd_sc_hd__a22o_2
X_3854_ _4394_/A _4574_/A vssd1 vssd1 vccd1 vccd1 _3855_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_6_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5119__A _6242_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3785_ _3850_/A _3862_/S _3838_/S vssd1 vssd1 vccd1 vccd1 _4510_/B sky130_fd_sc_hd__or3_1
XANTENNA__4023__A _6292_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5524_ _5524_/A _5524_/B vssd1 vssd1 vccd1 vccd1 _5524_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_6_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5455_ hold601/X _5377_/X _5454_/Y _5377_/A vssd1 vssd1 vccd1 vccd1 _5455_/X sky130_fd_sc_hd__o2bb2a_1
XANTENNA__4958__A _5054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5553__S _5553_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4406_ hold222/X _4405_/X _4428_/S vssd1 vssd1 vccd1 vccd1 _4406_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5386_ _5386_/A _5386_/B vssd1 vssd1 vccd1 vccd1 _5387_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_10_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4337_ _4510_/A _4438_/A vssd1 vssd1 vccd1 vccd1 _4345_/S sky130_fd_sc_hd__nor2_4
X_4268_ _4268_/A _4268_/B vssd1 vssd1 vccd1 vccd1 _4273_/C sky130_fd_sc_hd__nor2_1
X_3219_ _4228_/A _3566_/B _3219_/C vssd1 vssd1 vccd1 vccd1 _3219_/X sky130_fd_sc_hd__or3_1
XANTENNA__3475__B1 _4309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4898__S0 _6318_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6007_ _5339_/A _6005_/X _6006_/Y hold435/X _5995_/Y vssd1 vssd1 vccd1 vccd1 _6007_/X
+ sky130_fd_sc_hd__o32a_1
X_4199_ hold173/X _4200_/S _5673_/C1 _4198_/X vssd1 vssd1 vccd1 vccd1 _4199_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_96_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4727__A0 hold560/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3950__A1 _6245_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3772__A _4309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5463__S _5518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3702__A1 _3473_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold290 _3531_/X vssd1 vssd1 vccd1 vccd1 _6086_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4258__A2 _3770_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5455__B2 _5377_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4807__S _5053_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3947__A _6243_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3536__A4 _4679_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3570_ _5097_/B _5265_/B _4637_/B _5265_/A vssd1 vssd1 vccd1 vccd1 _3570_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_70_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5391__A0 _6417_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5240_ hold560/X _5239_/X _5240_/S vssd1 vssd1 vccd1 vccd1 _5240_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_11_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5171_ _6270_/Q _5170_/X _5193_/S vssd1 vssd1 vccd1 vccd1 _5171_/X sky130_fd_sc_hd__mux2_1
X_4122_ _5088_/B _4122_/B vssd1 vssd1 vccd1 vccd1 _4122_/X sky130_fd_sc_hd__or2_1
X_4053_ hold235/X hold77/X hold212/X hold120/X _5676_/C1 _4200_/S vssd1 vssd1 vccd1
+ vccd1 _4053_/X sky130_fd_sc_hd__mux4_2
XANTENNA__4717__S _4727_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput3 io_in[23] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_78_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4955_ _6110_/Q hold63/A _6093_/Q _6138_/Q _5051_/S0 _5052_/S1 vssd1 vssd1 vccd1
+ vccd1 _4955_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_86_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3906_ _6417_/Q _3905_/X _3906_/S vssd1 vssd1 vccd1 vccd1 _3906_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_52_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4452__S _4455_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout140_A _3952_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4886_ _6325_/Q _4866_/X _4867_/B vssd1 vssd1 vccd1 vccd1 _4886_/Y sky130_fd_sc_hd__a21boi_1
X_3837_ _6162_/Q hold43/A _3838_/S vssd1 vssd1 vccd1 vccd1 _3837_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_6_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4709__B1 _5075_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4185__A1 _5217_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3768_ _3723_/X _6032_/A _4391_/A2 vssd1 vssd1 vccd1 vccd1 _3768_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_42_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5507_ _6418_/Q _5506_/X _5558_/S vssd1 vssd1 vccd1 vccd1 _5507_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_30_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3699_ _3473_/A _3697_/X _3365_/B vssd1 vssd1 vccd1 vccd1 _3699_/Y sky130_fd_sc_hd__o21ai_4
X_6487_ _6487_/A vssd1 vssd1 vccd1 vccd1 _6487_/X sky130_fd_sc_hd__buf_1
XFILLER_0_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5438_ _5436_/X _5438_/B vssd1 vssd1 vccd1 vccd1 _5440_/A sky130_fd_sc_hd__and2b_1
XANTENNA__5685__A1 _6298_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5369_ _6392_/Q _6427_/Q vssd1 vssd1 vccd1 vccd1 _5441_/A sky130_fd_sc_hd__and2_4
XANTENNA__3696__B1 _5339_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold617_A _6298_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5193__S _5193_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3923__B2 _4427_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6078__RESET_B fanout169/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5428__A1 _6323_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_24_wb_clk_i_A _6404_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output34_A _6415_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4939__B1 _4938_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4740_ hold95/A _6407_/Q hold53/A _6176_/Q _4326_/B _5358_/A0 vssd1 vssd1 vccd1 vccd1
+ _4740_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_28_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4671_ _3691_/B _4670_/X _4673_/B vssd1 vssd1 vccd1 vccd1 _4671_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_16_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3622_ _3622_/A _5956_/B vssd1 vssd1 vccd1 vccd1 _3623_/A sky130_fd_sc_hd__or2_2
X_6410_ _6410_/CLK _6410_/D vssd1 vssd1 vccd1 vccd1 _6410_/Q sky130_fd_sc_hd__dfxtp_1
X_6341_ _6373_/CLK _6341_/D vssd1 vssd1 vccd1 vccd1 _6341_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_101_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3553_ _5578_/A _3581_/A vssd1 vssd1 vccd1 vccd1 _3553_/Y sky130_fd_sc_hd__nor2_4
X_3484_ _5560_/D _3484_/B _3484_/C vssd1 vssd1 vccd1 vccd1 _3485_/A sky130_fd_sc_hd__or3_1
X_6272_ _6295_/CLK _6272_/D fanout177/X vssd1 vssd1 vccd1 vccd1 _6272_/Q sky130_fd_sc_hd__dfstp_4
X_5223_ _6365_/Q _6364_/Q _6367_/Q _6366_/Q vssd1 vssd1 vccd1 vccd1 _5225_/A sky130_fd_sc_hd__or4_1
X_5154_ _5154_/A _5154_/B _5148_/X vssd1 vssd1 vccd1 vccd1 _5154_/X sky130_fd_sc_hd__or3b_1
XFILLER_0_47_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4105_ hold83/A _3784_/X _3786_/X _6158_/Q _4104_/X vssd1 vssd1 vccd1 vccd1 _4108_/A
+ sky130_fd_sc_hd__a221o_1
X_5085_ hold304/X _5241_/S _5084_/X vssd1 vssd1 vccd1 vccd1 _5085_/Y sky130_fd_sc_hd__o21ai_1
X_4036_ _5087_/A _4059_/A vssd1 vssd1 vccd1 vccd1 _4036_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_79_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5987_ hold677/X _5982_/S _5979_/Y hold264/X vssd1 vssd1 vccd1 vccd1 _5987_/X sky130_fd_sc_hd__a22o_1
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4938_ _5054_/A _4938_/B vssd1 vssd1 vccd1 vccd1 _4938_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_74_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4869_ _4863_/B _4868_/X _5058_/S vssd1 vssd1 vccd1 vccd1 _4869_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_34_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4568__D _4604_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5658__A1 _5695_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4357__S _4360_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmax_cap87 _3510_/B vssd1 vssd1 vccd1 vccd1 _5270_/A sky130_fd_sc_hd__buf_2
XFILLER_0_85_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6259__RESET_B fanout177/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5217__A _5217_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3960__A _6040_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4857__C1 _5557_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4775__B _5060_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6048__A _6048_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4085__A0 _6421_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4624__A2 _4615_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5910_ _5909_/A _5909_/B _5932_/S vssd1 vssd1 vccd1 vccd1 _5910_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_88_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5841_ _6326_/Q _5840_/X _5930_/S vssd1 vssd1 vccd1 vccd1 _5841_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_91_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4388__A1 _5690_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5772_ _5771_/X _6321_/Q _5772_/S vssd1 vssd1 vccd1 vccd1 _5773_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_56_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4723_ _6273_/Q _4681_/X _4722_/X _5371_/A vssd1 vssd1 vccd1 vccd1 _4723_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_8_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5337__B1 _5977_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4730__S _5240_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4654_ _6245_/Q _6339_/Q _4674_/S vssd1 vssd1 vccd1 vccd1 _4654_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3899__B1 _6245_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3605_ _6487_/A _3605_/B vssd1 vssd1 vccd1 vccd1 _3652_/B sky130_fd_sc_hd__or2_1
XFILLER_0_12_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4585_ _6419_/Q _4569_/X _4570_/X _6270_/Q vssd1 vssd1 vccd1 vccd1 _4585_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4031__A _6246_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3536_ _4224_/A _3725_/B _5578_/B _4679_/D _3535_/X vssd1 vssd1 vccd1 vccd1 _3536_/X
+ sky130_fd_sc_hd__o41a_1
X_6324_ _6421_/CLK _6324_/D fanout175/X vssd1 vssd1 vccd1 vccd1 _6324_/Q sky130_fd_sc_hd__dfrtp_4
X_6255_ _6403_/CLK _6255_/D fanout179/X vssd1 vssd1 vccd1 vccd1 _6255_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5206_ _5206_/A _5206_/B _5110_/A vssd1 vssd1 vccd1 vccd1 _5206_/X sky130_fd_sc_hd__or3b_1
X_3467_ _5935_/A _6392_/Q vssd1 vssd1 vccd1 vccd1 _3467_/X sky130_fd_sc_hd__or2_1
XFILLER_0_58_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3398_ _5258_/B _5256_/B vssd1 vssd1 vccd1 vccd1 _3400_/B sky130_fd_sc_hd__and2_2
XANTENNA__4685__B _5715_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6186_ _6209_/CLK hold40/X vssd1 vssd1 vccd1 vccd1 hold39/A sky130_fd_sc_hd__dfxtp_1
X_5137_ _5560_/A _6293_/Q _5135_/Y _5136_/X vssd1 vssd1 vccd1 vccd1 _5137_/X sky130_fd_sc_hd__o22a_1
X_5068_ hold447/X _5067_/X _5068_/S vssd1 vssd1 vccd1 vccd1 _5068_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_79_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4019_ _4394_/A _4019_/B vssd1 vssd1 vccd1 vccd1 _4021_/A sky130_fd_sc_hd__nor2_1
XANTENNA__3823__B1 _3794_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3483__C _5740_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4303__A1 _6064_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4854__A2 _4752_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3814__B1 _3781_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold108 _4341_/X vssd1 vssd1 vccd1 vccd1 _6102_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold119 _3514_/X vssd1 vssd1 vccd1 vccd1 _6088_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4370_ hold254/X _4384_/S _5673_/C1 _4369_/X vssd1 vssd1 vccd1 vccd1 _4370_/X sky130_fd_sc_hd__o211a_1
X_3321_ _3525_/A _3525_/B vssd1 vssd1 vccd1 vccd1 _3537_/A sky130_fd_sc_hd__nand2_1
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3252_ _3374_/A _3725_/B _4679_/D vssd1 vssd1 vccd1 vccd1 _3573_/B sky130_fd_sc_hd__or3_2
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6040_ _6040_/A _6063_/S vssd1 vssd1 vccd1 vccd1 _6040_/Y sky130_fd_sc_hd__nor2_1
X_3183_ _4744_/A _3183_/B _4744_/B _3525_/A vssd1 vssd1 vccd1 vccd1 _3238_/C sky130_fd_sc_hd__and4b_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6047__A1 _6057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4725__S _4731_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_16_wb_clk_i _6404_/CLK vssd1 vssd1 vccd1 vccd1 _6432_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__5558__A0 _6423_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5824_ _6377_/Q _5849_/S _4883_/X vssd1 vssd1 vccd1 vccd1 _5824_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_8_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5755_ _5755_/A _5755_/B vssd1 vssd1 vccd1 vccd1 _5757_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_97_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4706_ _4704_/X _4705_/X _5102_/A vssd1 vssd1 vccd1 vccd1 _4706_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4460__S _4464_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5686_ _6274_/Q _5589_/X _5610_/X _6448_/Q vssd1 vssd1 vccd1 vccd1 _5694_/B sky130_fd_sc_hd__a22o_1
X_4637_ _4637_/A _4637_/B _3574_/B vssd1 vssd1 vccd1 vccd1 _4674_/S sky130_fd_sc_hd__or3b_4
XANTENNA__4533__A1 _6292_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold620 _6397_/Q vssd1 vssd1 vccd1 vccd1 _5937_/B sky130_fd_sc_hd__buf_1
XFILLER_0_69_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold642 _6421_/Q vssd1 vssd1 vccd1 vccd1 hold642/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold631 _6418_/Q vssd1 vssd1 vccd1 vccd1 hold631/X sky130_fd_sc_hd__dlygate4sd3_1
X_4568_ _5725_/A _4568_/B _4568_/C _4604_/S vssd1 vssd1 vccd1 vccd1 _4568_/X sky130_fd_sc_hd__and4_2
Xhold653 _6268_/Q vssd1 vssd1 vccd1 vccd1 hold653/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5730__B1 _3477_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3519_ _5733_/A _5323_/C _3519_/C _3519_/D vssd1 vssd1 vccd1 vccd1 _3521_/C sky130_fd_sc_hd__or4_1
X_6307_ _6433_/CLK _6307_/D fanout173/X vssd1 vssd1 vccd1 vccd1 _6307_/Q sky130_fd_sc_hd__dfrtp_1
Xhold675 _6307_/Q vssd1 vssd1 vccd1 vccd1 _3695_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold664 _5358_/X vssd1 vssd1 vccd1 vccd1 _6318_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4499_ _4148_/X hold243/X _4500_/S vssd1 vssd1 vccd1 vccd1 _6198_/D sky130_fd_sc_hd__mux2_1
X_6238_ _6297_/CLK _6238_/D fanout176/X vssd1 vssd1 vccd1 vccd1 _6238_/Q sky130_fd_sc_hd__dfstp_1
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6169_ _6407_/CLK hold68/X vssd1 vssd1 vccd1 vccd1 hold67/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6038__A1 _6057_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5797__A0 _6323_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5721__A0 _6272_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4524__A1 _6267_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4288__A0 _6267_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5230__A _6419_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5004__A2 _5060_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3870_ _3870_/A _3870_/B _3870_/C vssd1 vssd1 vccd1 vccd1 _4401_/B sky130_fd_sc_hd__nand3_1
XANTENNA__4212__B1 _4228_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3685__A _5518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5540_ hold577/X _5539_/X _6060_/S vssd1 vssd1 vccd1 vccd1 _5540_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6203__RESET_B fanout174/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5471_ _6423_/Q _5470_/X _5471_/S vssd1 vssd1 vccd1 vccd1 _5471_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_1_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4422_ _4156_/A _3811_/Y _4415_/X vssd1 vssd1 vccd1 vccd1 _4423_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_41_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4353_ hold138/X _3881_/X _4360_/S vssd1 vssd1 vccd1 vccd1 _4353_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_22_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3304_ _3304_/A _3304_/B _3304_/C vssd1 vssd1 vccd1 vccd1 _4756_/A sky130_fd_sc_hd__and3_2
X_4284_ _4284_/A _4639_/B _4284_/C vssd1 vssd1 vccd1 vccd1 _4727_/S sky130_fd_sc_hd__and3_4
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3235_ _3534_/B _3215_/C _3566_/B _3232_/Y _3234_/X vssd1 vssd1 vccd1 vccd1 _3235_/X
+ sky130_fd_sc_hd__o311a_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6023_ _3046_/A _6021_/X _6022_/Y hold414/X _5995_/Y vssd1 vssd1 vccd1 vccd1 _6023_/X
+ sky130_fd_sc_hd__o32a_1
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3166_ _4685_/A _3594_/A vssd1 vssd1 vccd1 vccd1 _4541_/C sky130_fd_sc_hd__nor2_2
X_3097_ _3525_/A _4685_/A vssd1 vssd1 vccd1 vccd1 _3100_/B sky130_fd_sc_hd__nor2_2
XANTENNA__4455__S _4455_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout170_A fanout181/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xci2406_z80_192 vssd1 vssd1 vccd1 vccd1 ci2406_z80_192/HI io_oeb[11] sky130_fd_sc_hd__conb_1
Xfanout69 _3723_/X vssd1 vssd1 vccd1 vccd1 _3724_/A sky130_fd_sc_hd__buf_4
XFILLER_0_9_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3999_ _6071_/Q _3715_/X _3794_/X _6139_/Q _3998_/X vssd1 vssd1 vccd1 vccd1 _4000_/B
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4203__B1 _5675_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5807_ _5806_/X hold552/X _5931_/S vssd1 vssd1 vccd1 vccd1 _5807_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5951__B1 _4323_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5738_ _4767_/A _5734_/X _5735_/X _5737_/X vssd1 vssd1 vccd1 vccd1 _5739_/B sky130_fd_sc_hd__a211o_1
XFILLER_0_9_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5669_ _6272_/Q _5589_/X _5610_/X _6446_/Q _5668_/X vssd1 vssd1 vccd1 vccd1 _5670_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_20_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold450 _5355_/X vssd1 vssd1 vccd1 vccd1 _6316_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold472 _6372_/Q vssd1 vssd1 vccd1 vccd1 _5755_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold461 _6343_/Q vssd1 vssd1 vccd1 vccd1 _4158_/A sky130_fd_sc_hd__buf_1
XANTENNA__5315__A _5315_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold483 _4536_/X vssd1 vssd1 vccd1 vccd1 _6237_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold494 _6375_/Q vssd1 vssd1 vccd1 vccd1 _5791_/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5034__B _6057_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold647_A _6273_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3489__B _5472_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3548__A2 _4767_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3952__B _3952_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5170__A1 _6294_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3720__A2 _4382_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6056__A _6057_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4681__B1 _5740_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3399__B _3400_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4971_ _6362_/Q _4970_/X _5557_/S vssd1 vssd1 vccd1 vccd1 _4971_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_25_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3922_ hold203/X hold51/X hold209/X hold126/X _5676_/C1 _5676_/B1 vssd1 vssd1 vccd1
+ vccd1 _3922_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_18_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3853_ _3852_/B _3852_/C _3852_/D _4111_/A vssd1 vssd1 vccd1 vccd1 _3853_/Y sky130_fd_sc_hd__a31oi_1
XFILLER_0_39_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6127__SET_B fanout180/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3784_ _3863_/A _3850_/B _3861_/S vssd1 vssd1 vccd1 vccd1 _3784_/X sky130_fd_sc_hd__and3_4
XANTENNA__4023__B _6295_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5523_ _5503_/A _5503_/B _5512_/A _5522_/X vssd1 vssd1 vccd1 vccd1 _5524_/B sky130_fd_sc_hd__a31o_1
XFILLER_0_14_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4958__B _4958_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5454_ _5454_/A _5454_/B vssd1 vssd1 vccd1 vccd1 _5454_/Y sky130_fd_sc_hd__xnor2_1
X_5385_ _5383_/X _5385_/B vssd1 vssd1 vccd1 vccd1 _5386_/B sky130_fd_sc_hd__nand2b_1
X_4405_ _4402_/X _4403_/X _4404_/X _4427_/S vssd1 vssd1 vccd1 vccd1 _4405_/X sky130_fd_sc_hd__a22o_2
XFILLER_0_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4336_ hold169/X _4205_/X _4336_/S vssd1 vssd1 vccd1 vccd1 _4336_/X sky130_fd_sc_hd__mux2_1
X_4267_ _3573_/A _3511_/A _3386_/A vssd1 vssd1 vccd1 vccd1 _4268_/B sky130_fd_sc_hd__a21oi_1
X_6067__4 _6270_/CLK vssd1 vssd1 vccd1 vccd1 _6125_/CLK sky130_fd_sc_hd__inv_2
X_3218_ _3183_/B _3116_/A _3534_/B _3232_/A vssd1 vssd1 vccd1 vccd1 _3219_/C sky130_fd_sc_hd__o22a_1
XANTENNA__3475__A1 _5553_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6006_ _6040_/A _6026_/B vssd1 vssd1 vccd1 vccd1 _6006_/Y sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_31_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6374_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_4198_ _6115_/Q _4198_/B _4427_/S vssd1 vssd1 vccd1 vccd1 _4198_/X sky130_fd_sc_hd__or3_1
XANTENNA__4898__S1 _6090_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3149_ _6257_/Q _6258_/Q vssd1 vssd1 vccd1 vccd1 _3373_/A sky130_fd_sc_hd__and2b_2
XFILLER_0_69_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4214__A _4214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5152__B2 _6293_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold280 _6071_/Q vssd1 vssd1 vccd1 vccd1 hold280/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold291 _6412_/Q vssd1 vssd1 vccd1 vccd1 hold291/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_14_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__3218__A1 _3183_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4966__A1 _6381_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3947__B _6244_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4194__A2 _6026_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5170_ _3074_/Y _6294_/Q _5192_/S vssd1 vssd1 vccd1 vccd1 _5170_/X sky130_fd_sc_hd__mux2_1
X_4121_ _4121_/A _4121_/B vssd1 vssd1 vccd1 vccd1 _4121_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_46_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4654__A0 _6245_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4249__A3 _4734_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4052_ hold17/X _4425_/A2 _5597_/B vssd1 vssd1 vccd1 vccd1 _4052_/X sky130_fd_sc_hd__o21a_1
Xinput4 io_in[24] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__buf_2
X_4954_ hold340/X _4953_/X _5068_/S vssd1 vssd1 vccd1 vccd1 _4954_/X sky130_fd_sc_hd__mux2_1
X_3905_ _4040_/A _5111_/B _5210_/B _3758_/Y _3898_/X vssd1 vssd1 vccd1 vccd1 _3905_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_19_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4885_ _4882_/B _4884_/X _5058_/S vssd1 vssd1 vccd1 vccd1 _4885_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_34_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3836_ _3850_/B _3835_/X _3850_/A vssd1 vssd1 vccd1 vccd1 _3836_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_34_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3767_ hold496/X _4158_/B _3766_/X vssd1 vssd1 vccd1 vccd1 _6032_/A sky130_fd_sc_hd__a21oi_4
XANTENNA__5382__A1 _4788_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5506_ hold558/X _5505_/X _5557_/S vssd1 vssd1 vccd1 vccd1 _5506_/X sky130_fd_sc_hd__mux2_1
X_3698_ _3473_/A _3697_/X _3365_/B vssd1 vssd1 vccd1 vccd1 _3700_/C sky130_fd_sc_hd__o21a_1
X_6486_ _6487_/A vssd1 vssd1 vccd1 vccd1 _6486_/X sky130_fd_sc_hd__buf_1
X_5437_ _5450_/A _5436_/B _5436_/C vssd1 vssd1 vccd1 vccd1 _5438_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_100_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5368_ _5715_/A _6416_/Q _5365_/C _5386_/A vssd1 vssd1 vccd1 vccd1 _5368_/Y sky130_fd_sc_hd__o31ai_1
XFILLER_0_10_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5299_ _4228_/A _3770_/A _5266_/A vssd1 vssd1 vccd1 vccd1 _5299_/X sky130_fd_sc_hd__o21a_1
X_4319_ _4767_/A _4320_/B vssd1 vssd1 vccd1 vccd1 _4319_/X sky130_fd_sc_hd__and2_1
XANTENNA__4740__S0 _4326_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3999__A2 _3715_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6377__RESET_B fanout168/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4643__S _4674_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4948__A1 _6380_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5373__A1 input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5474__S _5518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5676__A2 _4198_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4939__A1 _6268_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4670_ _4669_/X _6244_/Q _4675_/S vssd1 vssd1 vccd1 vccd1 _4670_/X sky130_fd_sc_hd__mux2_1
X_3621_ _3621_/A vssd1 vssd1 vccd1 vccd1 _3625_/A sky130_fd_sc_hd__inv_2
X_3552_ _4270_/B _4747_/D _3519_/C _6389_/Q vssd1 vssd1 vccd1 vccd1 _3559_/C sky130_fd_sc_hd__o211a_1
X_6340_ _6343_/CLK _6340_/D vssd1 vssd1 vccd1 vccd1 _6340_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__3914__A2 _3715_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3483_ _3483_/A _4615_/A _5740_/A _3639_/B vssd1 vssd1 vccd1 vccd1 _3484_/C sky130_fd_sc_hd__and4_1
X_6271_ _6271_/CLK _6271_/D fanout170/X vssd1 vssd1 vccd1 vccd1 _6271_/Q sky130_fd_sc_hd__dfstp_4
X_5222_ _6239_/Q _6297_/Q _5239_/S vssd1 vssd1 vccd1 vccd1 _5222_/X sky130_fd_sc_hd__mux2_1
X_5153_ _3759_/A _5118_/X _5152_/X vssd1 vssd1 vccd1 vccd1 _5154_/B sky130_fd_sc_hd__a21o_1
XANTENNA__5413__A _5441_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4104_ hold99/A _3779_/X _3781_/X hold79/A vssd1 vssd1 vccd1 vccd1 _4104_/X sky130_fd_sc_hd__a22o_1
X_5084_ _4070_/A _5083_/Y _5080_/Y _5371_/A vssd1 vssd1 vccd1 vccd1 _5084_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_47_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4035_ _4035_/A _5182_/A vssd1 vssd1 vccd1 vccd1 _4059_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_79_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5559__S _6060_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4463__S _4464_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5986_ hold264/X _5982_/S _5979_/Y hold269/X vssd1 vssd1 vccd1 vccd1 _5986_/X sky130_fd_sc_hd__a22o_1
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4937_ _4936_/X _4935_/X _5053_/S vssd1 vssd1 vccd1 vccd1 _4938_/B sky130_fd_sc_hd__mux2_2
X_4868_ _6376_/Q _6324_/Q _6315_/Q vssd1 vssd1 vccd1 vccd1 _4868_/X sky130_fd_sc_hd__mux2_1
X_3819_ _4394_/A _4594_/A vssd1 vssd1 vccd1 vccd1 _4408_/A sky130_fd_sc_hd__xnor2_1
X_4799_ _5773_/A _4799_/B vssd1 vssd1 vccd1 vccd1 _4799_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4211__B _4222_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3669__A1 _5096_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4638__S _4674_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5323__A _5733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4618__B1 _4617_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5217__B _6246_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5932__S _5932_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5649__A2 _4382_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6048__B _6063_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5840_ _5929_/A1 _5839_/X _4900_/Y vssd1 vssd1 vccd1 vccd1 _5840_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_29_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5585__A1 _3183_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5771_ _6373_/Q _5849_/S _4804_/X vssd1 vssd1 vccd1 vccd1 _5771_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_71_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4722_ _6273_/Q _4680_/X _5075_/B hold443/X vssd1 vssd1 vccd1 vccd1 _4722_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_29_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5337__A1 _4568_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4653_ _6044_/A _4673_/B vssd1 vssd1 vccd1 vccd1 _4653_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__3899__A1 _6243_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3604_ _4637_/A _3587_/X _3597_/Y _3603_/X vssd1 vssd1 vccd1 vccd1 _3645_/B sky130_fd_sc_hd__o22a_1
X_4584_ _4001_/B _4394_/B _4604_/S vssd1 vssd1 vccd1 vccd1 _4584_/X sky130_fd_sc_hd__mux2_1
X_3535_ _4685_/A _6256_/Q _3725_/B _3535_/D vssd1 vssd1 vccd1 vccd1 _3535_/X sky130_fd_sc_hd__or4_1
X_6323_ _6399_/CLK _6323_/D fanout173/X vssd1 vssd1 vccd1 vccd1 _6323_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_12_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6254_ _6403_/CLK _6254_/D fanout179/X vssd1 vssd1 vccd1 vccd1 _6254_/Q sky130_fd_sc_hd__dfrtp_4
X_3466_ _6390_/Q _3466_/B vssd1 vssd1 vccd1 vccd1 _3545_/B sky130_fd_sc_hd__or2_1
XANTENNA__5842__S _5931_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5205_ _5205_/A _5205_/B _5112_/A vssd1 vssd1 vccd1 vccd1 _5206_/A sky130_fd_sc_hd__or3b_1
X_3397_ _5096_/A _5941_/A vssd1 vssd1 vccd1 vccd1 _5256_/B sky130_fd_sc_hd__and2_1
X_6185_ _6430_/CLK _6185_/D vssd1 vssd1 vccd1 vccd1 _6185_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4458__S _4464_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5136_ _5135_/A _5135_/B _5077_/A vssd1 vssd1 vccd1 vccd1 _5136_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_98_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5067_ _6367_/Q _5066_/X _5557_/S vssd1 vssd1 vccd1 vccd1 _5067_/X sky130_fd_sc_hd__mux2_1
X_4018_ _4019_/B vssd1 vssd1 vccd1 vccd1 _4020_/B sky130_fd_sc_hd__inv_2
XFILLER_0_79_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5969_ input8/X hold632/X _5975_/S vssd1 vssd1 vccd1 vccd1 _6417_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_47_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3110__B _3451_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3780__B _3862_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4368__S _4428_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6321__RESET_B fanout181/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3301__A _3594_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4116__B _6342_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5567__B2 _4637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5319__A1 _5715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4790__A2 _5060_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4542__A2 _5733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold109 _6110_/Q vssd1 vssd1 vccd1 vccd1 hold109/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6292__SET_B fanout177/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3320_ _3359_/B _4758_/C vssd1 vssd1 vccd1 vccd1 _4755_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3251_ _3374_/A _3725_/B _4679_/D vssd1 vssd1 vccd1 vccd1 _4639_/C sky130_fd_sc_hd__nor3_4
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3182_ _5303_/A _3285_/B vssd1 vssd1 vccd1 vccd1 _5733_/A sky130_fd_sc_hd__nor2_4
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5823_ _5820_/X _5821_/Y _5932_/S vssd1 vssd1 vccd1 vccd1 _5823_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_63_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4741__S _5053_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4230__A1 _5096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5754_ _6372_/Q _5755_/B vssd1 vssd1 vccd1 vccd1 _5769_/A sky130_fd_sc_hd__and2_1
XFILLER_0_44_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4781__A2 _5557_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4705_ hold484/X _4299_/A _4727_/S vssd1 vssd1 vccd1 vccd1 _4705_/X sky130_fd_sc_hd__mux2_1
X_5685_ _6298_/Q _5587_/X _5588_/X _6440_/Q vssd1 vssd1 vccd1 vccd1 _5694_/A sky130_fd_sc_hd__a22o_1
X_4636_ _6032_/A _4636_/B vssd1 vssd1 vccd1 vccd1 _4636_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_8_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold621 _5953_/X vssd1 vssd1 vccd1 vccd1 hold621/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold610 _6293_/Q vssd1 vssd1 vccd1 vccd1 hold610/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5730__A1 _5740_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6306_ _6432_/CLK _6306_/D fanout175/X vssd1 vssd1 vccd1 vccd1 _6306_/Q sky130_fd_sc_hd__dfrtp_1
Xhold643 _6422_/Q vssd1 vssd1 vccd1 vccd1 hold643/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold632 _6417_/Q vssd1 vssd1 vccd1 vccd1 hold632/X sky130_fd_sc_hd__dlygate4sd3_1
X_4567_ _5339_/C _4567_/B _4604_/S vssd1 vssd1 vccd1 vccd1 _4567_/Y sky130_fd_sc_hd__nor3_4
Xhold654 _4696_/X vssd1 vssd1 vccd1 vccd1 _6268_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3518_ _3496_/A _3517_/X _3510_/B _6405_/Q vssd1 vssd1 vccd1 vccd1 _3519_/D sky130_fd_sc_hd__a2bb2o_1
Xhold676 _6305_/Q vssd1 vssd1 vccd1 vccd1 _4191_/S sky130_fd_sc_hd__dlygate4sd3_1
Xhold665 _6399_/Q vssd1 vssd1 vccd1 vccd1 _3619_/A sky130_fd_sc_hd__dlygate4sd3_1
X_4498_ _4102_/X hold263/X _4500_/S vssd1 vssd1 vccd1 vccd1 _6197_/D sky130_fd_sc_hd__mux2_1
X_3449_ _3469_/A _5956_/B vssd1 vssd1 vccd1 vccd1 _3449_/X sky130_fd_sc_hd__or2_4
X_6237_ _6270_/CLK _6237_/D fanout176/X vssd1 vssd1 vccd1 vccd1 _6237_/Q sky130_fd_sc_hd__dfstp_1
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6168_ _6407_/CLK hold54/X vssd1 vssd1 vccd1 vccd1 hold53/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5119_ _6242_/Q _5119_/B vssd1 vssd1 vccd1 vccd1 _5121_/A sky130_fd_sc_hd__xnor2_1
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6038__A2 _4958_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5601__A _5603_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6099_ _6221_/CLK hold98/X vssd1 vssd1 vccd1 vccd1 hold97/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5549__A1 _6057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold425_A _6342_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3980__B1 _6292_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5721__A1 hold534/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6029__A2 _6063_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5788__B2 _5747_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5788__A1 _5932_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5230__B _6418_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5470_ _5468_/Y _5469_/X _5560_/D vssd1 vssd1 vccd1 vccd1 _5470_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_26_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4421_ hold132/X _4420_/X _4428_/S vssd1 vssd1 vccd1 vccd1 _4421_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5392__S _5447_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4352_ _4510_/A _4483_/A vssd1 vssd1 vccd1 vccd1 _4360_/S sky130_fd_sc_hd__nor2_4
X_3303_ _3281_/Y _3318_/D _3302_/X _3269_/X vssd1 vssd1 vccd1 vccd1 _3304_/C sky130_fd_sc_hd__a31o_1
X_4283_ _4639_/B _4284_/C vssd1 vssd1 vccd1 vccd1 _5226_/C sky130_fd_sc_hd__and2_1
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3234_ _3573_/A _4228_/A _5303_/B _3566_/B _3233_/X vssd1 vssd1 vccd1 vccd1 _3234_/X
+ sky130_fd_sc_hd__o41a_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6022_ _6022_/A _6026_/B vssd1 vssd1 vccd1 vccd1 _6022_/Y sky130_fd_sc_hd__nor2_1
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3165_ _5303_/B _5256_/A vssd1 vssd1 vccd1 vccd1 _3632_/B sky130_fd_sc_hd__or2_2
XANTENNA__5228__A0 _5221_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3096_ _3206_/A _3683_/B vssd1 vssd1 vccd1 vccd1 _3483_/A sky130_fd_sc_hd__and2_1
XFILLER_0_89_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout163_A _4326_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xci2406_z80_193 vssd1 vssd1 vccd1 vccd1 ci2406_z80_193/HI io_oeb[12] sky130_fd_sc_hd__conb_1
Xci2406_z80_182 vssd1 vssd1 vccd1 vccd1 ci2406_z80_182/HI io_oeb[0] sky130_fd_sc_hd__conb_1
XANTENNA__4471__S _4473_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3998_ _6094_/Q _3789_/X _3791_/X _6195_/Q vssd1 vssd1 vccd1 vccd1 _3998_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4203__A1 _6314_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5806_ _6324_/Q _5805_/X _5852_/S vssd1 vssd1 vccd1 vccd1 _5806_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_29_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout59 _5815_/S vssd1 vssd1 vccd1 vccd1 _5932_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_0_72_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5737_ _4639_/B _5359_/A _3770_/A _5736_/X _6392_/Q vssd1 vssd1 vccd1 vccd1 _5737_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_0_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5668_ _6384_/Q _5600_/X _5665_/X _5594_/Y vssd1 vssd1 vccd1 vccd1 _5668_/X sky130_fd_sc_hd__a22o_1
X_4619_ input8/X _4631_/B vssd1 vssd1 vccd1 vccd1 _4619_/X sky130_fd_sc_hd__and2_1
X_5599_ _5599_/A _5603_/D vssd1 vssd1 vccd1 vccd1 _5610_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_4_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold440 _5645_/X vssd1 vssd1 vccd1 vccd1 _6339_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold462 _5695_/X vssd1 vssd1 vccd1 vccd1 _6343_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold451 _6227_/Q vssd1 vssd1 vccd1 vccd1 hold451/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold473 _5763_/X vssd1 vssd1 vccd1 vccd1 _6372_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold484 _6363_/Q vssd1 vssd1 vccd1 vccd1 hold484/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6438__SET_B fanout171/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold495 _5802_/X vssd1 vssd1 vccd1 vccd1 _6375_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout76_A _3718_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold375_A _6337_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold542_A _6386_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3489__C _5739_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4381__S _4428_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5942__B2 _5096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4053__S0 _5676_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_1_wb_clk_i clkbuf_leaf_6_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6413_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_clkbuf_leaf_43_wb_clk_i_A clkbuf_leaf_6_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__4715__A1_N _6272_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4970_ _6418_/Q _4969_/X _5930_/S vssd1 vssd1 vccd1 vccd1 _4970_/X sky130_fd_sc_hd__mux2_1
X_3921_ hold13/X _4425_/A2 _5597_/B vssd1 vssd1 vccd1 vccd1 _3921_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_86_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3852_ _4111_/A _3852_/B _3852_/C _3852_/D vssd1 vssd1 vccd1 vccd1 _3855_/A sky130_fd_sc_hd__nand4_1
XANTENNA__3539__A3 _3528_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5522_ _5501_/B _5510_/B _5554_/A vssd1 vssd1 vccd1 vccd1 _5522_/X sky130_fd_sc_hd__o21a_1
X_3783_ hold138/X _4483_/A _4438_/A hold97/X vssd1 vssd1 vccd1 vccd1 _3783_/X sky130_fd_sc_hd__o22a_1
X_5453_ _5438_/B _5440_/B _5436_/X vssd1 vssd1 vccd1 vccd1 _5454_/B sky130_fd_sc_hd__a21o_1
X_5384_ _5450_/A _5383_/B _5383_/C vssd1 vssd1 vccd1 vccd1 _5385_/B sky130_fd_sc_hd__a21o_1
X_4404_ hold257/X hold61/X hold266/X hold93/X _5676_/C1 _5676_/B1 vssd1 vssd1 vccd1
+ vccd1 _4404_/X sky130_fd_sc_hd__mux4_2
X_4335_ hold147/X _4148_/X _4336_/S vssd1 vssd1 vccd1 vccd1 _4335_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_10_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4266_ _3132_/B _5315_/A _4265_/X _3289_/A _4230_/X vssd1 vssd1 vccd1 vccd1 _4273_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_5_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3217_ _3549_/A _3502_/A _3232_/C _3216_/X vssd1 vssd1 vccd1 vccd1 _3228_/A sky130_fd_sc_hd__a31o_1
XANTENNA__4672__A1 _5715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3475__A2 _6425_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4466__S _4473_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4197_ _6314_/Q _4197_/B vssd1 vssd1 vccd1 vccd1 _5690_/S sky130_fd_sc_hd__nand2_8
X_6005_ _5560_/D _6004_/X _6026_/B vssd1 vssd1 vccd1 vccd1 _6005_/X sky130_fd_sc_hd__o21a_1
X_3148_ _3525_/A _3278_/A _3116_/A vssd1 vssd1 vccd1 vccd1 _3148_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_69_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3079_ _3079_/A vssd1 vssd1 vccd1 vccd1 _3079_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_92_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold270 _5986_/X vssd1 vssd1 vccd1 vccd1 _6429_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold281 _6195_/Q vssd1 vssd1 vccd1 vccd1 hold281/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold292 _6192_/Q vssd1 vssd1 vccd1 vccd1 hold292/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5000__S _5058_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3926__B1 _3781_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6020__A2_N _6054_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4120_ _4075_/A _4058_/B _4060_/X vssd1 vssd1 vccd1 vccd1 _4121_/B sky130_fd_sc_hd__o21ai_1
X_4051_ _4424_/A _4022_/Y _4050_/X vssd1 vssd1 vccd1 vccd1 _4051_/Y sky130_fd_sc_hd__o21ai_1
Xinput5 io_in[25] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__4654__A1 _6339_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4953_ _6361_/Q _4952_/X _5557_/S vssd1 vssd1 vccd1 vccd1 _4953_/X sky130_fd_sc_hd__mux2_1
X_3904_ _5119_/B vssd1 vssd1 vccd1 vccd1 _5210_/B sky130_fd_sc_hd__inv_2
XFILLER_0_52_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4315__A _4316_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4884_ _6377_/Q _6325_/Q _4901_/S vssd1 vssd1 vccd1 vccd1 _4884_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_74_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3835_ hold45/A hold73/A _3838_/S vssd1 vssd1 vccd1 vccd1 _3835_/X sky130_fd_sc_hd__mux2_1
X_3766_ hold623/X hold637/X _4142_/S _3765_/X vssd1 vssd1 vccd1 vccd1 _3766_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_42_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5505_ hold558/X _5377_/X _5504_/Y _5441_/A vssd1 vssd1 vccd1 vccd1 _5505_/X sky130_fd_sc_hd__a22o_1
X_6485_ _6487_/A vssd1 vssd1 vccd1 vccd1 _6485_/X sky130_fd_sc_hd__buf_1
XFILLER_0_72_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3697_ _5096_/B _3675_/X _3679_/X _5518_/S _3611_/A vssd1 vssd1 vccd1 vccd1 _3697_/X
+ sky130_fd_sc_hd__o2111a_4
X_5436_ _5450_/A _5436_/B _5436_/C vssd1 vssd1 vccd1 vccd1 _5436_/X sky130_fd_sc_hd__and3_1
XFILLER_0_100_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5367_ _5386_/A vssd1 vssd1 vccd1 vccd1 _5367_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3696__A2 _4197_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5298_ _3482_/A _5317_/B _5297_/X _3404_/Y vssd1 vssd1 vccd1 vccd1 _5298_/X sky130_fd_sc_hd__o22a_1
X_4318_ _4767_/A _4318_/B vssd1 vssd1 vccd1 vccd1 _4321_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_10_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4249_ _4255_/B _5328_/B _4734_/B _3297_/X _3109_/B vssd1 vssd1 vccd1 vccd1 _4249_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__6127__D _6127_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4740__S1 _5358_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4924__S _5058_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4884__A1 _6325_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5061__B2 _4867_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5061__A1 _5061_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6087__RESET_B fanout174/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3620_ _5935_/A _3620_/B vssd1 vssd1 vccd1 vccd1 _3621_/A sky130_fd_sc_hd__or2_2
X_3551_ _5096_/A _5578_/A _5325_/A _3654_/B vssd1 vssd1 vccd1 vccd1 _3551_/X sky130_fd_sc_hd__or4_1
X_3482_ _3482_/A _5560_/D _3639_/B vssd1 vssd1 vccd1 vccd1 _3482_/X sky130_fd_sc_hd__and3_1
X_6270_ _6270_/CLK _6270_/D fanout176/X vssd1 vssd1 vccd1 vccd1 _6270_/Q sky130_fd_sc_hd__dfstp_4
X_5221_ _5220_/X _5208_/X _5150_/Y _6297_/Q vssd1 vssd1 vccd1 vccd1 _5221_/X sky130_fd_sc_hd__o2bb2a_2
XANTENNA__3678__A2 _3770_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5152_ _3758_/Y _5128_/Y _5149_/X _6293_/Q _5241_/S vssd1 vssd1 vccd1 vccd1 _5152_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_47_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4103_ _4102_/X hold296/X _4206_/S vssd1 vssd1 vccd1 vccd1 _6073_/D sky130_fd_sc_hd__mux2_1
X_5083_ _5239_/S _5746_/A vssd1 vssd1 vccd1 vccd1 _5083_/Y sky130_fd_sc_hd__nand2_1
X_4034_ _4035_/A _5182_/A vssd1 vssd1 vccd1 vccd1 _4034_/X sky130_fd_sc_hd__or2_1
XFILLER_0_63_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5985_ hold269/X _5982_/S _5979_/Y _5518_/S vssd1 vssd1 vccd1 vccd1 _5985_/X sky130_fd_sc_hd__a22o_1
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4936_ _6216_/Q _6153_/Q _6193_/Q _6069_/Q _5051_/S0 _5052_/S1 vssd1 vssd1 vccd1
+ vccd1 _4936_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_10 _6298_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4867_ _4866_/X _4867_/B _4867_/C vssd1 vssd1 vccd1 vccd1 _4867_/X sky130_fd_sc_hd__and3b_1
XFILLER_0_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3818_ _4594_/A vssd1 vssd1 vccd1 vccd1 _3818_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3366__A1 _5061_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4798_ _4797_/X _6320_/Q _5825_/S vssd1 vssd1 vccd1 vccd1 _4799_/B sky130_fd_sc_hd__mux2_1
X_3749_ _3952_/A _3755_/C _5715_/C _3747_/B _6336_/Q vssd1 vssd1 vccd1 vccd1 _3749_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_15_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6399_ _6399_/CLK _6399_/D fanout174/X vssd1 vssd1 vccd1 vccd1 _6399_/Q sky130_fd_sc_hd__dfrtp_1
X_5419_ hold608/X _5418_/X _5447_/S vssd1 vssd1 vccd1 vccd1 _5419_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4919__S _5053_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4654__S _4674_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5043__B2 _4867_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5043__A1 _5061_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4251__C1 _4222_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5594__A2 _5603_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4554__B1 _3725_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5217__C _6247_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4829__S _4901_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4857__A1 _6323_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5806__A0 _6324_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5282__A1 _5077_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5770_ _5782_/B _5770_/B vssd1 vssd1 vccd1 vccd1 _5770_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_90_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4721_ hold405/X _4314_/S _4727_/S vssd1 vssd1 vccd1 vccd1 _4721_/X sky130_fd_sc_hd__mux2_1
X_4652_ _5715_/B _4650_/Y _4651_/X hold328/X _4635_/Y vssd1 vssd1 vccd1 vccd1 _4652_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_0_4_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3603_ _4347_/C _5327_/A _4348_/A _3603_/D vssd1 vssd1 vccd1 vccd1 _3603_/X sky130_fd_sc_hd__or4_1
XFILLER_0_71_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3899__A2 _6244_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3209__A _3594_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4583_ _5695_/A1 hold441/X _4546_/Y _4582_/X vssd1 vssd1 vccd1 vccd1 _4583_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_12_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3534_ _3534_/A _3534_/B vssd1 vssd1 vccd1 vccd1 _3535_/D sky130_fd_sc_hd__or2_1
X_6322_ _6421_/CLK _6322_/D fanout175/X vssd1 vssd1 vccd1 vccd1 _6322_/Q sky130_fd_sc_hd__dfrtp_4
X_6253_ _6403_/CLK _6253_/D fanout174/X vssd1 vssd1 vccd1 vccd1 _6253_/Q sky130_fd_sc_hd__dfrtp_1
X_3465_ _3465_/A _3465_/B vssd1 vssd1 vccd1 vccd1 _3471_/B sky130_fd_sc_hd__or2_1
X_5204_ _3333_/S _6300_/Q _5111_/A _5111_/B vssd1 vssd1 vccd1 vccd1 _5205_/A sky130_fd_sc_hd__a211o_1
XANTENNA__4848__A1 _6323_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3396_ _3394_/X _3395_/Y _3686_/A vssd1 vssd1 vccd1 vccd1 _3396_/Y sky130_fd_sc_hd__o21ai_1
X_6184_ _6344_/CLK _6184_/D vssd1 vssd1 vccd1 vccd1 _6184_/Q sky130_fd_sc_hd__dfxtp_1
X_5135_ _5135_/A _5135_/B vssd1 vssd1 vccd1 vccd1 _5135_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5066_ _6423_/Q _5065_/X _5930_/S vssd1 vssd1 vccd1 vccd1 _5066_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_79_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4017_ _4017_/A _4017_/B vssd1 vssd1 vccd1 vccd1 _4019_/B sky130_fd_sc_hd__nor2_1
XANTENNA__3823__A2 _3715_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5968_ input9/X hold637/X _5975_/S vssd1 vssd1 vccd1 vccd1 _6416_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_47_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3587__A1 _3278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4919_ _4918_/X _4917_/X _5053_/S vssd1 vssd1 vccd1 vccd1 _4920_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_74_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5899_ _5887_/A _5898_/X _5933_/S vssd1 vssd1 vccd1 vccd1 _5899_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_7_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3119__A _4679_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4222__B _4222_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3780__C _3838_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3814__A2 _3779_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3578__A1 _4541_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4542__A3 _3770_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3250_ _5313_/A _3686_/A vssd1 vssd1 vccd1 vccd1 _4637_/A sky130_fd_sc_hd__or2_4
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3181_ _3091_/X _3144_/X _3277_/A _3100_/B vssd1 vssd1 vccd1 vccd1 _3189_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3266__B1 _4637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3211__B _5715_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5822_ _5821_/A _5821_/B _5820_/X vssd1 vssd1 vccd1 vccd1 _5836_/B sky130_fd_sc_hd__o21ba_1
XANTENNA__3569__A1 _3482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5753_ _5236_/S _6417_/Q _3580_/A _5735_/X vssd1 vssd1 vccd1 vccd1 _5755_/B sky130_fd_sc_hd__o31a_1
XFILLER_0_60_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4704_ _6270_/Q _4681_/X _4703_/X _5371_/A vssd1 vssd1 vccd1 vccd1 _4704_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_44_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4861__S0 _5051_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4323__A _4323_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5684_ _5695_/A1 _3063_/A _5571_/Y _5683_/X vssd1 vssd1 vccd1 vccd1 _5684_/X sky130_fd_sc_hd__a22o_1
X_4635_ _3691_/B _4673_/B _5715_/B vssd1 vssd1 vccd1 vccd1 _4635_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_0_44_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5853__S _5931_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold611 _5169_/X vssd1 vssd1 vccd1 vccd1 _6293_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_25_wb_clk_i _6404_/CLK vssd1 vssd1 vccd1 vccd1 _6295_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold600 _6296_/Q vssd1 vssd1 vccd1 vccd1 hold600/X sky130_fd_sc_hd__dlygate4sd3_1
X_4566_ _4566_/A _4566_/B vssd1 vssd1 vccd1 vccd1 _4566_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_8_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold633 _6302_/Q vssd1 vssd1 vccd1 vccd1 hold633/X sky130_fd_sc_hd__dlygate4sd3_1
X_6305_ _6305_/CLK _6305_/D fanout180/X vssd1 vssd1 vccd1 vccd1 _6305_/Q sky130_fd_sc_hd__dfrtp_4
X_3517_ _4070_/A _3952_/B _3330_/X _4214_/A vssd1 vssd1 vccd1 vccd1 _3517_/X sky130_fd_sc_hd__o211a_1
Xhold622 _5954_/X vssd1 vssd1 vccd1 vccd1 _6393_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold644 _6423_/Q vssd1 vssd1 vccd1 vccd1 hold644/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4469__S _4473_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5730__A2 _5729_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold655 _6291_/Q vssd1 vssd1 vccd1 vccd1 hold655/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold666 _6387_/Q vssd1 vssd1 vccd1 vccd1 hold666/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold677 _6430_/Q vssd1 vssd1 vccd1 vccd1 hold677/X sky130_fd_sc_hd__dlygate4sd3_1
X_4497_ _4054_/X hold284/X _4500_/S vssd1 vssd1 vccd1 vccd1 _6196_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_12_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3448_ _3469_/A _3448_/B vssd1 vssd1 vccd1 vccd1 _3465_/A sky130_fd_sc_hd__nor2_1
X_6236_ _6295_/CLK _6236_/D fanout176/X vssd1 vssd1 vccd1 vccd1 _6236_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA__5494__A1 _6057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3379_ _5303_/A _3379_/B vssd1 vssd1 vccd1 vccd1 _3581_/B sky130_fd_sc_hd__or2_2
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6167_ _6414_/CLK _6167_/D vssd1 vssd1 vccd1 vccd1 _6167_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5118_ _6293_/Q _5117_/X _5347_/B vssd1 vssd1 vccd1 vccd1 _5118_/X sky130_fd_sc_hd__mux2_1
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6119__RESET_B fanout173/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5601__B _5691_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6098_ _6355_/CLK _6098_/D vssd1 vssd1 vccd1 vccd1 _6098_/Q sky130_fd_sc_hd__dfxtp_1
X_5049_ hold405/X _5048_/X _5557_/S vssd1 vssd1 vccd1 vccd1 _5049_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_94_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_2_3__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6404_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_94_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_33_wb_clk_i_A clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__3791__B _3862_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5485__A1 _4313_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5230__C _6423_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4143__A _6022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4420_ _4417_/X _4418_/X _4419_/X _4427_/S vssd1 vssd1 vccd1 vccd1 _4420_/X sky130_fd_sc_hd__a22o_2
XFILLER_0_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3723__A1 _3611_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4351_ hold304/X _4350_/Y _5347_/A vssd1 vssd1 vccd1 vccd1 _6107_/D sky130_fd_sc_hd__mux2_1
XANTENNA__4289__S _6064_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3302_ _3337_/A _3549_/B _5360_/C _3299_/X _3195_/B vssd1 vssd1 vccd1 vccd1 _3302_/X
+ sky130_fd_sc_hd__o2111a_1
X_4282_ hold321/X _4281_/X _5727_/S vssd1 vssd1 vccd1 vccd1 _4282_/X sky130_fd_sc_hd__mux2_1
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3233_ _4522_/B _5258_/B _3233_/C _3233_/D vssd1 vssd1 vccd1 vccd1 _3233_/X sky130_fd_sc_hd__or4_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6021_ _6057_/A _6020_/X _6026_/B vssd1 vssd1 vccd1 vccd1 _6021_/X sky130_fd_sc_hd__o21a_1
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3164_ _5303_/B _5256_/A vssd1 vssd1 vccd1 vccd1 _3164_/Y sky130_fd_sc_hd__nor2_2
XANTENNA__3222__A _3254_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3095_ _3573_/A _3278_/A vssd1 vssd1 vccd1 vccd1 _3683_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_49_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xci2406_z80_194 vssd1 vssd1 vccd1 vccd1 ci2406_z80_194/HI io_oeb[13] sky130_fd_sc_hd__conb_1
Xci2406_z80_183 vssd1 vssd1 vccd1 vccd1 ci2406_z80_183/HI io_oeb[1] sky130_fd_sc_hd__conb_1
XANTENNA__5149__A _6304_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3997_ _6218_/Q _3784_/X _3786_/X _6155_/Q _3996_/X vssd1 vssd1 vccd1 vccd1 _4000_/A
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4203__A2 _5597_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5805_ _5773_/A _5804_/X _4863_/Y vssd1 vssd1 vccd1 vccd1 _5805_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_91_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5736_ _5313_/A _3451_/C _5935_/A vssd1 vssd1 vccd1 vccd1 _5736_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_29_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5667_ _6438_/Q _5588_/X _5603_/X _6376_/Q _5666_/X vssd1 vssd1 vccd1 vccd1 _5670_/A
+ sky130_fd_sc_hd__a221o_1
X_4618_ hold247/X _4615_/X _4617_/Y _4613_/X vssd1 vssd1 vccd1 vccd1 _4618_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_13_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5598_ _3722_/X _5690_/S _5590_/X _5597_/X _5691_/S vssd1 vssd1 vccd1 vccd1 _5598_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4911__A0 _6326_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4549_ _5574_/A _5578_/B _4210_/A vssd1 vssd1 vccd1 vccd1 _4550_/C sky130_fd_sc_hd__o21a_1
Xhold463 _6117_/Q vssd1 vssd1 vccd1 vccd1 _3491_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold430 _4573_/X vssd1 vssd1 vccd1 vccd1 _6242_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold441 _6244_/Q vssd1 vssd1 vccd1 vccd1 hold441/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold452 _4526_/X vssd1 vssd1 vccd1 vccd1 _6227_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold474 _6340_/Q vssd1 vssd1 vccd1 vccd1 _3062_/A sky130_fd_sc_hd__buf_1
Xhold496 _6336_/Q vssd1 vssd1 vccd1 vccd1 hold496/X sky130_fd_sc_hd__clkbuf_2
Xhold485 _5719_/X vssd1 vssd1 vccd1 vccd1 _6363_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6219_ _6331_/CLK _6219_/D vssd1 vssd1 vccd1 vccd1 _6219_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4228__A _4228_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3786__B _3850_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4902__A0 _4900_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3307__A _5578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5458__A1 _5560_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3139__A_N _3656_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3042__A _6389_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3920_ _3724_/A _5251_/A _3910_/Y vssd1 vssd1 vccd1 vccd1 _3920_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_86_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3851_ _3852_/B _3852_/C _3852_/D vssd1 vssd1 vccd1 vccd1 _4574_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_39_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6444__SET_B fanout171/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3782_ _3863_/A _3862_/S _3861_/S vssd1 vssd1 vccd1 vccd1 _4438_/A sky130_fd_sc_hd__or3_4
XFILLER_0_6_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5521_ _5519_/X _5521_/B vssd1 vssd1 vccd1 vccd1 _5524_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_14_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5452_ _5450_/X _5452_/B vssd1 vssd1 vccd1 vccd1 _5454_/A sky130_fd_sc_hd__and2b_1
X_5383_ _5450_/A _5383_/B _5383_/C vssd1 vssd1 vccd1 vccd1 _5383_/X sky130_fd_sc_hd__and3_1
X_4403_ hold11/X _4425_/A2 _5597_/B vssd1 vssd1 vccd1 vccd1 _4403_/X sky130_fd_sc_hd__o21a_1
X_4334_ hold145/X _4102_/X _4336_/S vssd1 vssd1 vccd1 vccd1 _4334_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_10_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5449__A1 _4882_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4265_ _3534_/A _4222_/B _4255_/Y _5315_/B vssd1 vssd1 vccd1 vccd1 _4265_/X sky130_fd_sc_hd__a31o_1
X_6004_ _4321_/A _4807_/X _5400_/Y _5992_/Y vssd1 vssd1 vccd1 vccd1 _6004_/X sky130_fd_sc_hd__o22a_1
X_3216_ _3216_/A _3233_/C _3373_/A vssd1 vssd1 vccd1 vccd1 _3216_/X sky130_fd_sc_hd__and3_1
X_4196_ hold25/X _4425_/A2 _5597_/B vssd1 vssd1 vccd1 vccd1 _4196_/X sky130_fd_sc_hd__o21a_1
X_3147_ _3206_/B vssd1 vssd1 vccd1 vccd1 _3633_/B sky130_fd_sc_hd__inv_2
XANTENNA__3475__A3 _3473_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3880__B1 _4382_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4482__S _4482_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5621__A1 _5695_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3078_ _3078_/A vssd1 vssd1 vccd1 vccd1 _3078_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_9_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4214__C _5258_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_40_wb_clk_i clkbuf_leaf_6_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6447_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_5719_ _6270_/Q hold484/X _5723_/S vssd1 vssd1 vccd1 vccd1 _5719_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3699__B1 _3365_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3127__A _4228_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold271 _6155_/Q vssd1 vssd1 vccd1 vccd1 hold271/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold260 _4428_/X vssd1 vssd1 vccd1 vccd1 _6135_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 _6141_/Q vssd1 vssd1 vccd1 vccd1 hold282/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold293 _4493_/X vssd1 vssd1 vccd1 vccd1 _6192_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_hold652_A _6297_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5488__S _5518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4820__C1 _4313_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5679__B2 _6422_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5679__A1 _6385_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3037__A _3656_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4050_ _3724_/A _6048_/A _4425_/A2 vssd1 vssd1 vccd1 vccd1 _4050_/X sky130_fd_sc_hd__o21a_1
Xinput6 io_in[26] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__clkbuf_2
X_4952_ _6417_/Q _4951_/X _5930_/S vssd1 vssd1 vccd1 vccd1 _4952_/X sky130_fd_sc_hd__mux2_1
X_3903_ _4073_/B _3981_/A _6243_/Q vssd1 vssd1 vccd1 vccd1 _5119_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_19_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4883_ _6325_/Q _4752_/X _4751_/B vssd1 vssd1 vccd1 vccd1 _4883_/X sky130_fd_sc_hd__a21o_1
X_3834_ _3862_/S _3834_/B vssd1 vssd1 vccd1 vccd1 _3834_/Y sky130_fd_sc_hd__nor2_1
X_3765_ _4040_/A _5111_/A _3749_/X _3764_/X _5247_/A vssd1 vssd1 vccd1 vccd1 _3765_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_42_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5427__A _5441_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3696_ _3682_/X _4197_/B _4391_/A2 _3695_/X _5339_/A vssd1 vssd1 vccd1 vccd1 _4510_/A
+ sky130_fd_sc_hd__a41o_4
XFILLER_0_6_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6484_ _6487_/A vssd1 vssd1 vccd1 vccd1 _6484_/X sky130_fd_sc_hd__buf_1
X_5504_ _5504_/A vssd1 vssd1 vccd1 vccd1 _5504_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4590__A1 _6420_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4590__B2 _6271_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5435_ _6438_/Q _4863_/B _5518_/S vssd1 vssd1 vccd1 vccd1 _5436_/C sky130_fd_sc_hd__mux2_1
X_5366_ _5715_/A _6433_/Q _5365_/X vssd1 vssd1 vccd1 vccd1 _5386_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_10_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5297_ _4224_/A _3572_/A _3581_/A _5266_/B vssd1 vssd1 vccd1 vccd1 _5297_/X sky130_fd_sc_hd__a31o_1
XANTENNA__5162__A _6419_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4477__S _4482_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4317_ _6064_/S _4314_/S _5724_/S _6273_/Q _4315_/X vssd1 vssd1 vccd1 vccd1 _4317_/X
+ sky130_fd_sc_hd__o221a_1
X_4248_ _4255_/B _5328_/B vssd1 vssd1 vccd1 vccd1 _4248_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_93_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4179_ _4179_/A _4179_/B vssd1 vssd1 vccd1 vccd1 _4179_/X sky130_fd_sc_hd__or2_1
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3410__A _4541_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5358__A0 _5358_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4030__B1 _6246_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6315__RESET_B fanout173/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5996__A2_N _6054_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5072__A _6032_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5011__S _5557_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3550_ _4685_/A _5096_/A _5324_/C _4734_/B _5291_/A vssd1 vssd1 vccd1 vccd1 _3559_/A
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_24_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5220_ _5120_/A _5219_/X _5218_/X _5215_/X vssd1 vssd1 vccd1 vccd1 _5220_/X sky130_fd_sc_hd__o211a_1
X_3481_ _3505_/A _3486_/B vssd1 vssd1 vccd1 vccd1 _3639_/B sky130_fd_sc_hd__or2_2
X_5151_ _3985_/A _5137_/X _5143_/Y _3761_/A vssd1 vssd1 vccd1 vccd1 _5154_/A sky130_fd_sc_hd__a22o_1
X_5082_ _5239_/S _5746_/A vssd1 vssd1 vccd1 vccd1 _5082_/X sky130_fd_sc_hd__and2_1
XFILLER_0_44_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4102_ _4099_/X _4100_/X _4101_/X _4427_/S vssd1 vssd1 vccd1 vccd1 _4102_/X sky130_fd_sc_hd__a22o_2
X_4033_ _3973_/A _3973_/B _3969_/B vssd1 vssd1 vccd1 vccd1 _5182_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5984_ _5518_/S _5982_/S _5979_/Y _3473_/A vssd1 vssd1 vccd1 vccd1 _6427_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_19_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4935_ _6109_/Q hold51/A _6092_/Q _6137_/Q _5051_/S0 _5052_/S1 vssd1 vssd1 vccd1
+ vccd1 _4935_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_74_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4866_ _6324_/Q _4866_/B vssd1 vssd1 vccd1 vccd1 _4866_/X sky130_fd_sc_hd__and2_1
XFILLER_0_34_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6001__A1 _5560_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_11 _6298_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4797_ _5849_/S _4795_/X _4796_/X _4783_/X vssd1 vssd1 vccd1 vccd1 _4797_/X sky130_fd_sc_hd__a31o_1
X_3817_ _3817_/A _3817_/B vssd1 vssd1 vccd1 vccd1 _4594_/A sky130_fd_sc_hd__nor2_2
X_3748_ _4134_/B vssd1 vssd1 vccd1 vccd1 _3748_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_42_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3679_ _3164_/Y _3553_/Y _3668_/C _3678_/X vssd1 vssd1 vccd1 vccd1 _3679_/X sky130_fd_sc_hd__a211o_1
XANTENNA__4996__A _5054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6398_ _6401_/CLK _6398_/D fanout178/X vssd1 vssd1 vccd1 vccd1 _6398_/Q sky130_fd_sc_hd__dfrtp_1
X_5418_ _6419_/Q _5417_/X _5471_/S vssd1 vssd1 vccd1 vccd1 _5418_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_30_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5349_ _5603_/A _5349_/B vssd1 vssd1 vccd1 vccd1 _5349_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__3405__A _4284_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4618__A2 _4615_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6034__A2_N _6054_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3794__B _3862_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5751__B1 _5747_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5217__D _6248_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4306__B2 _6064_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5514__B _6057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5267__C1 _4224_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output32_A _6287_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5665__S0 _5691_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5990__B1 _5739_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4720_ hold658/X _4719_/X _5447_/S vssd1 vssd1 vccd1 vccd1 _6272_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_44_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4651_ _3691_/B _4649_/X _4673_/B vssd1 vssd1 vccd1 vccd1 _4651_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_44_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3602_ _5560_/A _5270_/A _5324_/A _5480_/D vssd1 vssd1 vccd1 vccd1 _3603_/D sky130_fd_sc_hd__or4_1
X_4582_ _4564_/A _4579_/X _4581_/X vssd1 vssd1 vccd1 vccd1 _4582_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_101_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3533_ hold37/X _3449_/X _3457_/C _6390_/Q vssd1 vssd1 vccd1 vccd1 hold38/A sky130_fd_sc_hd__a22o_1
X_6321_ _6326_/CLK _6321_/D fanout181/X vssd1 vssd1 vccd1 vccd1 _6321_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_3_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6252_ _6403_/CLK _6252_/D fanout179/X vssd1 vssd1 vccd1 vccd1 _6252_/Q sky130_fd_sc_hd__dfrtp_1
X_3464_ _3464_/A _3471_/A _3464_/C vssd1 vssd1 vccd1 vccd1 _6395_/D sky130_fd_sc_hd__or3_1
XFILLER_0_58_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5203_ hold600/X _5202_/X _5347_/A vssd1 vssd1 vccd1 vccd1 _6296_/D sky130_fd_sc_hd__mux2_1
X_6183_ _6414_/CLK _6183_/D vssd1 vssd1 vccd1 vccd1 _6183_/Q sky130_fd_sc_hd__dfxtp_1
X_5134_ _5134_/A _5134_/B vssd1 vssd1 vccd1 vccd1 _5135_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__3225__A _3566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3395_ _5265_/A _3377_/Y _3389_/Y vssd1 vssd1 vccd1 vccd1 _3395_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5065_ _5929_/A1 _5064_/X _5054_/Y vssd1 vssd1 vccd1 vccd1 _5065_/X sky130_fd_sc_hd__a21bo_1
XANTENNA__3808__B1 _3791_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4016_ hold224/X _3715_/X _3794_/X _6140_/Q _4015_/X vssd1 vssd1 vccd1 vccd1 _4017_/B
+ sky130_fd_sc_hd__a221o_1
Xclkbuf_2_2__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_2__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
X_5967_ _4427_/X hold305/X _5967_/S vssd1 vssd1 vccd1 vccd1 _6414_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_90_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3587__A2 _3566_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4918_ _6215_/Q _6192_/Q _6152_/Q _6068_/Q _5052_/S1 _5358_/A0 vssd1 vssd1 vccd1
+ vccd1 _4918_/X sky130_fd_sc_hd__mux4_1
XANTENNA__4490__S _4491_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5898_ _5892_/Y _5897_/X _5932_/S vssd1 vssd1 vccd1 vccd1 _5898_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4536__A1 _6295_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4849_ _4843_/X _4848_/X _5058_/S vssd1 vssd1 vccd1 vccd1 _4849_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_99_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_23_wb_clk_i_A _6404_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4222__C _4541_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout99_A _4639_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4839__A2 _4313_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4147__S0 _5676_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3789__B _3862_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5496__S _6060_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5972__A0 input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6330__RESET_B fanout171/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5724__A0 _6274_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4527__A1 _6270_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3045__A _6425_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3180_ _3220_/A _3243_/B vssd1 vssd1 vccd1 vccd1 _3496_/A sky130_fd_sc_hd__or2_1
XANTENNA__5660__C1 _5676_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4215__B1 _4679_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5821_ _5821_/A _5821_/B vssd1 vssd1 vccd1 vccd1 _5821_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5752_ _5745_/A _5742_/A _5751_/X _5731_/X vssd1 vssd1 vccd1 vccd1 _5752_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_60_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4703_ _6270_/Q _4680_/X _5075_/B hold488/X vssd1 vssd1 vccd1 vccd1 _4703_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_44_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4861__S1 _5052_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5683_ _5683_/A _5683_/B vssd1 vssd1 vccd1 vccd1 _5683_/X sky130_fd_sc_hd__or2_1
XANTENNA__6241__D _6241_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4634_ _5069_/A _4678_/B vssd1 vssd1 vccd1 vccd1 _4636_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold612 _6402_/Q vssd1 vssd1 vccd1 vccd1 hold612/X sky130_fd_sc_hd__buf_1
Xhold601 _6325_/Q vssd1 vssd1 vccd1 vccd1 hold601/X sky130_fd_sc_hd__dlygate4sd3_1
X_4565_ _3798_/B _5249_/B _4604_/S vssd1 vssd1 vccd1 vccd1 _4566_/B sky130_fd_sc_hd__mux2_1
Xhold634 _5306_/X vssd1 vssd1 vccd1 vccd1 _6302_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6304_ _6403_/CLK _6304_/D fanout180/X vssd1 vssd1 vccd1 vccd1 _6304_/Q sky130_fd_sc_hd__dfrtp_4
Xhold623 _6305_/Q vssd1 vssd1 vccd1 vccd1 hold623/X sky130_fd_sc_hd__clkbuf_2
X_3516_ _3344_/A _4747_/D _4223_/B vssd1 vssd1 vccd1 vccd1 _3519_/C sky130_fd_sc_hd__a21oi_1
XFILLER_0_69_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold645 _6420_/Q vssd1 vssd1 vccd1 vccd1 hold645/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold678 _6305_/Q vssd1 vssd1 vccd1 vccd1 _4085_/S sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold656 _6090_/Q vssd1 vssd1 vccd1 vccd1 hold656/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold667 _6313_/Q vssd1 vssd1 vccd1 vccd1 hold667/X sky130_fd_sc_hd__dlygate4sd3_1
X_4496_ _4007_/X hold281/X _4500_/S vssd1 vssd1 vccd1 vccd1 _6195_/D sky130_fd_sc_hd__mux2_1
X_3447_ _5935_/A _3451_/C _5978_/A _6392_/Q vssd1 vssd1 vccd1 vccd1 _3448_/B sky130_fd_sc_hd__or4b_1
X_6235_ _6297_/CLK _6235_/D fanout176/X vssd1 vssd1 vccd1 vccd1 _6235_/Q sky130_fd_sc_hd__dfstp_1
X_3378_ _5303_/A _3379_/B vssd1 vssd1 vccd1 vccd1 _4347_/C sky130_fd_sc_hd__nor2_4
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5494__A2 _5377_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6166_ _6408_/CLK hold90/X vssd1 vssd1 vccd1 vccd1 hold89/A sky130_fd_sc_hd__dfxtp_1
X_5117_ _3760_/B _5108_/Y _5115_/Y _5116_/X vssd1 vssd1 vccd1 vccd1 _5117_/X sky130_fd_sc_hd__o22a_1
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4485__S _4491_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6097_ _6194_/CLK _6097_/D vssd1 vssd1 vccd1 vccd1 _6097_/Q sky130_fd_sc_hd__dfxtp_1
X_5048_ _6422_/Q _5047_/X _5930_/S vssd1 vssd1 vccd1 vccd1 _5048_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_79_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3402__B _3594_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5485__A2 _5377_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3248__A1 _6392_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3248__B2 _5313_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6116__SET_B fanout173/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5230__D _6422_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3420__A1 _3654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5173__A1 _6294_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5173__B2 _5371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3708__C1 _3365_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4350_ _4639_/B _5317_/B _4349_/X _3597_/Y vssd1 vssd1 vccd1 vccd1 _4350_/Y sky130_fd_sc_hd__o2bb2ai_1
X_3301_ _3594_/A _5328_/B vssd1 vssd1 vccd1 vccd1 _3549_/B sky130_fd_sc_hd__nand2_2
XANTENNA__3723__A2 _3473_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4281_ _6335_/Q _6317_/Q _4281_/S vssd1 vssd1 vccd1 vccd1 _4281_/X sky130_fd_sc_hd__mux2_1
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3232_ _3232_/A _3233_/C _3232_/C vssd1 vssd1 vccd1 vccd1 _3232_/Y sky130_fd_sc_hd__nand3_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6020_ _5454_/Y _6054_/B _6057_/B _4882_/B vssd1 vssd1 vccd1 vccd1 _6020_/X sky130_fd_sc_hd__o2bb2a_1
X_3163_ _3573_/A _3572_/A vssd1 vssd1 vccd1 vccd1 _5266_/A sky130_fd_sc_hd__and2_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3094_ _3289_/A _3183_/B _3254_/A vssd1 vssd1 vccd1 vccd1 _3278_/A sky130_fd_sc_hd__nand3b_4
XANTENNA__5633__C1 _5675_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6252__RESET_B fanout179/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3222__B _3566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3649__S input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xci2406_z80_184 vssd1 vssd1 vccd1 vccd1 ci2406_z80_184/HI io_oeb[2] sky130_fd_sc_hd__conb_1
Xci2406_z80_195 vssd1 vssd1 vccd1 vccd1 ci2406_z80_195/HI io_oeb[14] sky130_fd_sc_hd__conb_1
X_5804_ _5803_/X _6324_/Q _5825_/S vssd1 vssd1 vccd1 vccd1 _5804_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout149_A _4284_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3996_ _6111_/Q _3779_/X _3781_/X _6102_/Q vssd1 vssd1 vccd1 vccd1 _3996_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3411__A1 _5158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5735_ _5077_/A _4734_/B _3579_/B hold128/X vssd1 vssd1 vccd1 vccd1 _5735_/X sky130_fd_sc_hd__a31o_4
XFILLER_0_95_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5666_ _6296_/Q _5587_/X _5602_/X _6421_/Q vssd1 vssd1 vccd1 vccd1 _5666_/X sky130_fd_sc_hd__a22o_1
X_4617_ _5371_/A _5372_/C _4615_/X vssd1 vssd1 vccd1 vccd1 _4617_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_0_44_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold420 _6246_/Q vssd1 vssd1 vccd1 vccd1 hold420/X sky130_fd_sc_hd__dlygate4sd3_1
X_5597_ _6314_/Q _5597_/B _5597_/C vssd1 vssd1 vccd1 vccd1 _5597_/X sky130_fd_sc_hd__and3_1
X_4548_ _3343_/Y _4547_/Y _4541_/A vssd1 vssd1 vccd1 vccd1 _4548_/X sky130_fd_sc_hd__o21a_1
Xhold431 _6400_/Q vssd1 vssd1 vccd1 vccd1 _4616_/A sky130_fd_sc_hd__clkbuf_2
Xhold442 _4583_/X vssd1 vssd1 vccd1 vccd1 _6244_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold453 _6226_/Q vssd1 vssd1 vccd1 vccd1 hold453/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4372__C1 _5673_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold464 _6235_/Q vssd1 vssd1 vccd1 vccd1 hold464/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold475 _5658_/X vssd1 vssd1 vccd1 vccd1 _6340_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold486 _6225_/Q vssd1 vssd1 vccd1 vccd1 hold486/X sky130_fd_sc_hd__dlygate4sd3_1
X_4479_ _4405_/X hold218/X _4482_/S vssd1 vssd1 vccd1 vccd1 _4479_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3478__A1 _4323_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold497 _5609_/X vssd1 vssd1 vccd1 vccd1 _6336_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6218_ _6218_/CLK _6218_/D vssd1 vssd1 vccd1 vccd1 _6218_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6149_ _6221_/CLK hold50/X vssd1 vssd1 vccd1 vccd1 hold49/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__5624__C1 _5675_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3786__C _3838_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5155__A1 _6293_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5075__A _5931_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3307__B _5158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4418__B1 _5597_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3850_ _3850_/A _3850_/B _3850_/C vssd1 vssd1 vccd1 vccd1 _3852_/D sky130_fd_sc_hd__or3_1
XFILLER_0_73_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3781_ _3850_/A _3850_/B _3838_/S vssd1 vssd1 vccd1 vccd1 _3781_/X sky130_fd_sc_hd__and3_4
XANTENNA__5394__A1 _4807_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5520_ _5554_/A _5520_/B vssd1 vssd1 vccd1 vccd1 _5521_/B sky130_fd_sc_hd__or2_1
XANTENNA__5146__A1 _6342_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5146__B2 _6339_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5451_ _5450_/A _5450_/B _5450_/C vssd1 vssd1 vccd1 vccd1 _5452_/B sky130_fd_sc_hd__a21o_1
X_5382_ _6434_/Q _4788_/B _6427_/Q vssd1 vssd1 vccd1 vccd1 _5383_/C sky130_fd_sc_hd__mux2_1
XFILLER_0_22_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4402_ _3724_/A _5250_/B _4050_/X vssd1 vssd1 vccd1 vccd1 _4402_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_10_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4333_ hold297/X _4054_/X _4336_/S vssd1 vssd1 vccd1 vccd1 _6095_/D sky130_fd_sc_hd__mux2_1
X_4264_ _5603_/A vssd1 vssd1 vccd1 vccd1 _5599_/A sky130_fd_sc_hd__inv_2
X_3215_ _3293_/B _4224_/A _3215_/C _3566_/B vssd1 vssd1 vccd1 vccd1 _3215_/X sky130_fd_sc_hd__or4_1
XFILLER_0_66_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6003_ _5339_/A _6001_/X _6002_/Y hold437/X _5995_/Y vssd1 vssd1 vccd1 vccd1 _6003_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_0_66_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4195_ _3723_/X _4157_/Y _4194_/Y vssd1 vssd1 vccd1 vccd1 _4195_/X sky130_fd_sc_hd__a21o_1
X_3146_ _4224_/A _3278_/A vssd1 vssd1 vccd1 vccd1 _3206_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_77_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3077_ _6321_/Q vssd1 vssd1 vccd1 vccd1 _4809_/A sky130_fd_sc_hd__inv_2
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3979_ _6243_/Q _6244_/Q _6245_/Q vssd1 vssd1 vccd1 vccd1 _3979_/X sky130_fd_sc_hd__or3_1
XFILLER_0_45_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5718_ _6269_/Q hold416/X _5723_/S vssd1 vssd1 vccd1 vccd1 _5718_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5137__A1 _5560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5649_ _6196_/Q _4382_/B _4200_/S _6072_/Q _5675_/C1 vssd1 vssd1 vccd1 vccd1 _5651_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_32_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3699__A1 _3473_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5688__A2 _6313_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold250 _3504_/X vssd1 vssd1 vccd1 vccd1 _6087_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3127__B _3594_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold261 _6131_/Q vssd1 vssd1 vccd1 vccd1 hold261/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold294 _6308_/Q vssd1 vssd1 vccd1 vccd1 _5988_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold272 _6179_/Q vssd1 vssd1 vccd1 vccd1 hold272/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold283 _6167_/Q vssd1 vssd1 vccd1 vccd1 hold283/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4648__A0 _6244_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold645_A _6420_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3926__A2 _3779_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4848__S _6315_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5300__B2 _3573_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput7 io_in[27] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_36_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3988__A _6339_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4951_ _5929_/A1 _4950_/X _4938_/Y vssd1 vssd1 vccd1 vccd1 _4951_/X sky130_fd_sc_hd__a21bo_1
XANTENNA__4811__A0 _4807_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3902_ _6245_/Q _6295_/Q vssd1 vssd1 vccd1 vccd1 _3981_/A sky130_fd_sc_hd__or2_1
XFILLER_0_59_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4882_ _5054_/A _4882_/B vssd1 vssd1 vccd1 vccd1 _4882_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_86_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3833_ hold39/A hold55/A _3838_/S vssd1 vssd1 vccd1 vccd1 _3834_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_27_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3764_ _3985_/A _5130_/A _3756_/X _3332_/Y _3763_/X vssd1 vssd1 vccd1 vccd1 _3764_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_82_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4612__A _5740_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3695_ _3695_/A _4361_/B _4633_/C vssd1 vssd1 vccd1 vccd1 _3695_/X sky130_fd_sc_hd__or3b_1
X_6483_ _6487_/A vssd1 vssd1 vccd1 vccd1 _6483_/X sky130_fd_sc_hd__buf_1
X_5503_ _5503_/A _5503_/B vssd1 vssd1 vccd1 vccd1 _5504_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_42_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5434_ _5715_/A _6421_/Q vssd1 vssd1 vccd1 vccd1 _5436_/B sky130_fd_sc_hd__or2_1
XFILLER_0_100_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3550__B1 _4734_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5365_ _5553_/S _6416_/Q _5365_/C vssd1 vssd1 vccd1 vccd1 _5365_/X sky130_fd_sc_hd__and3_1
XFILLER_0_10_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4973__S0 _5051_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5296_ _3313_/X _5294_/X _5295_/X vssd1 vssd1 vccd1 vccd1 _5296_/X sky130_fd_sc_hd__a21o_1
X_4316_ _6064_/S _4316_/B vssd1 vssd1 vccd1 vccd1 _5724_/S sky130_fd_sc_hd__nand2_1
X_4247_ _5935_/A _5313_/A vssd1 vssd1 vccd1 vccd1 _4247_/X sky130_fd_sc_hd__or2_2
XANTENNA__5162__B _6418_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4178_ _4178_/A _4179_/B vssd1 vssd1 vccd1 vccd1 _4178_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_97_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4493__S _4500_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3129_ _4228_/A _3656_/A vssd1 vssd1 vccd1 vccd1 _3132_/B sky130_fd_sc_hd__and2b_2
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3410__B _4637_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3837__S _3838_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4522__A _5560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3129__A_N _4228_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3138__A _3254_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold595_A _6379_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4869__A0 _4863_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5072__B _5243_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5499__S _5518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5247__B _5247_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3480_ _3483_/A _3591_/B _3374_/A _4767_/A vssd1 vssd1 vccd1 vccd1 _3486_/B sky130_fd_sc_hd__o211a_1
XANTENNA__4955__S0 _5051_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5150_ _6304_/Q _5150_/B vssd1 vssd1 vccd1 vccd1 _5150_/Y sky130_fd_sc_hd__nand2_1
X_5081_ _5977_/S _5740_/A vssd1 vssd1 vccd1 vccd1 _5746_/A sky130_fd_sc_hd__or2_2
X_4101_ hold85/X hold143/X hold103/X hold246/X _5676_/C1 _4200_/S vssd1 vssd1 vccd1
+ vccd1 _4101_/X sky130_fd_sc_hd__mux4_1
X_4032_ _4059_/A _4032_/B vssd1 vssd1 vccd1 vccd1 _4035_/A sky130_fd_sc_hd__and2_1
Xclkbuf_2_1__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_9_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__5202__S _5243_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5037__A0 _6385_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5983_ _3473_/A _5982_/S _5979_/Y _3577_/A vssd1 vssd1 vccd1 vccd1 _6426_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_59_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4326__B _4326_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4934_ hold427/X _4933_/X _5068_/S vssd1 vssd1 vccd1 vccd1 _4934_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_19_wb_clk_i _6404_/CLK vssd1 vssd1 vccd1 vccd1 _6305_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_86_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_12 _3577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4865_ _6324_/Q _4866_/B vssd1 vssd1 vccd1 vccd1 _4867_/C sky130_fd_sc_hd__or2_1
X_4796_ _6372_/Q _4796_/B vssd1 vssd1 vccd1 vccd1 _4796_/X sky130_fd_sc_hd__or2_1
X_3816_ _6181_/Q _3715_/X _3794_/X _6212_/Q _3815_/X vssd1 vssd1 vccd1 vccd1 _3817_/B
+ sky130_fd_sc_hd__a221o_1
X_3747_ _6301_/Q _3747_/B vssd1 vssd1 vccd1 vccd1 _4134_/B sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_leaf_13_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_70_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3678_ _5265_/A _3770_/A _3677_/Y vssd1 vssd1 vccd1 vccd1 _3678_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_42_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6397_ _6397_/CLK _6397_/D fanout174/X vssd1 vssd1 vccd1 vccd1 _6397_/Q sky130_fd_sc_hd__dfrtp_1
X_5417_ _5413_/Y _5415_/X _5416_/X _5560_/D vssd1 vssd1 vccd1 vccd1 _5417_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_2_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4488__S _4491_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5348_ _5077_/A _5347_/A _5315_/A _5347_/Y vssd1 vssd1 vccd1 vccd1 _5348_/X sky130_fd_sc_hd__a31o_1
X_5279_ _3573_/A _4685_/A _5322_/A _5276_/X _3334_/C vssd1 vssd1 vccd1 vccd1 _5279_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__5028__A0 _6421_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5579__A1 _3654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xmax_cap58 _4756_/Y vssd1 vssd1 vccd1 vccd1 _5056_/A2 sky130_fd_sc_hd__buf_4
XANTENNA_clkbuf_leaf_52_wb_clk_i_A clkbuf_leaf_6_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__4251__A1 _3254_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_hold510_A _6384_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold608_A _6322_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3794__C _3838_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5751__A1 _5932_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3762__A0 _6336_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5267__B1 _5317_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5022__S _5060_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5019__A0 _6384_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5665__S1 _5690_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5990__A1 _3611_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5258__A _5578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4650_ _6040_/A _4673_/B vssd1 vssd1 vccd1 vccd1 _4650_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_56_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput10 io_in[30] vssd1 vssd1 vccd1 vccd1 _6403_/D sky130_fd_sc_hd__buf_1
X_3601_ _4765_/A _5324_/B vssd1 vssd1 vccd1 vccd1 _4348_/A sky130_fd_sc_hd__or2_1
X_6320_ _6421_/CLK _6320_/D fanout175/X vssd1 vssd1 vccd1 vccd1 _6320_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4581_ hold435/X _4567_/Y _4568_/X _6443_/Q _4580_/X vssd1 vssd1 vccd1 vccd1 _4581_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__6206__RESET_B fanout174/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3532_ hold33/X _3449_/X _3471_/C vssd1 vssd1 vccd1 vccd1 hold34/A sky130_fd_sc_hd__a21o_1
XFILLER_0_12_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6251_ _6403_/CLK _6251_/D fanout179/X vssd1 vssd1 vccd1 vccd1 _6251_/Q sky130_fd_sc_hd__dfrtp_1
X_3463_ _3466_/B _3453_/B _3462_/X _3449_/X _3465_/B vssd1 vssd1 vccd1 vccd1 _3464_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_58_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5202_ _4087_/Y _5201_/X _5243_/S vssd1 vssd1 vccd1 vccd1 _5202_/X sky130_fd_sc_hd__mux2_1
X_6182_ _6408_/CLK _6182_/D vssd1 vssd1 vccd1 vccd1 _6182_/Q sky130_fd_sc_hd__dfxtp_1
X_5133_ _5133_/A _5133_/B vssd1 vssd1 vccd1 vccd1 _5134_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__3225__B _3566_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3394_ _4318_/B _5322_/D _3394_/C _3394_/D vssd1 vssd1 vccd1 vccd1 _3394_/X sky130_fd_sc_hd__or4_1
XFILLER_0_74_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5064_ _6334_/Q _5928_/A2 _5928_/B1 _5063_/X vssd1 vssd1 vccd1 vccd1 _5064_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_79_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4015_ _6095_/Q _3789_/X _3791_/X _6196_/Q vssd1 vssd1 vccd1 vccd1 _4015_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4337__A _4510_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3241__A _4679_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout179_A fanout180/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4728__A1_N _6274_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5966_ _4420_/X hold236/X _5967_/S vssd1 vssd1 vccd1 vccd1 _5966_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_74_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5897_ _5896_/X _5887_/A _5931_/S vssd1 vssd1 vccd1 vccd1 _5897_/X sky130_fd_sc_hd__mux2_1
X_4917_ _6108_/Q _6091_/Q hold97/A _6136_/Q _5052_/S1 _5051_/S0 vssd1 vssd1 vccd1
+ vccd1 _4917_/X sky130_fd_sc_hd__mux4_1
X_4848_ _6375_/Q _6323_/Q _6315_/Q vssd1 vssd1 vccd1 vccd1 _4848_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_43_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4779_ _6319_/Q _5825_/S _5850_/B1 _4778_/X _5054_/A vssd1 vssd1 vccd1 vccd1 _4779_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_99_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3135__B _3573_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4946__S _5060_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4147__S1 _5676_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4247__A _5935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3983__A0 _6339_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3061__A _3061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5660__B1 _5676_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5820_ _5836_/A _5820_/B vssd1 vssd1 vccd1 vccd1 _5820_/X sky130_fd_sc_hd__or2_1
XFILLER_0_84_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5751_ _5932_/S _5745_/Y _5747_/A _5750_/X vssd1 vssd1 vccd1 vccd1 _5751_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_71_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4702_ hold648/X _4701_/X _4732_/S vssd1 vssd1 vccd1 vccd1 _6269_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_71_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5682_ _6273_/Q _5589_/X _5603_/X _6377_/Q _5681_/X vssd1 vssd1 vccd1 vccd1 _5683_/B
+ sky130_fd_sc_hd__a221o_1
X_4633_ _5988_/C _4633_/B _4633_/C _4633_/D vssd1 vssd1 vccd1 vccd1 _4678_/B sky130_fd_sc_hd__and4_1
Xhold602 _5460_/X vssd1 vssd1 vccd1 vccd1 _6325_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4564_ _4564_/A vssd1 vssd1 vccd1 vccd1 _4566_/A sky130_fd_sc_hd__inv_2
Xhold624 _6258_/Q vssd1 vssd1 vccd1 vccd1 hold624/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_6303_ _6403_/CLK _6303_/D fanout179/X vssd1 vssd1 vccd1 vccd1 _6303_/Q sky130_fd_sc_hd__dfrtp_4
Xhold635 _6301_/Q vssd1 vssd1 vccd1 vccd1 hold635/X sky130_fd_sc_hd__dlygate4sd3_1
X_3515_ _3657_/A _3337_/B _4734_/B _3337_/Y _3600_/B vssd1 vssd1 vccd1 vccd1 _3515_/X
+ sky130_fd_sc_hd__a32o_1
Xhold613 _6295_/Q vssd1 vssd1 vccd1 vccd1 hold613/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold679 _6305_/Q vssd1 vssd1 vccd1 vccd1 _3906_/S sky130_fd_sc_hd__buf_1
X_6234_ _6270_/CLK _6234_/D fanout176/X vssd1 vssd1 vccd1 vccd1 _6234_/Q sky130_fd_sc_hd__dfstp_1
Xhold657 _4327_/X vssd1 vssd1 vccd1 vccd1 _6090_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold668 _5350_/X vssd1 vssd1 vccd1 vccd1 _6313_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold646 _6271_/Q vssd1 vssd1 vccd1 vccd1 hold646/X sky130_fd_sc_hd__dlygate4sd3_1
X_4495_ _3965_/X hold244/X _4500_/S vssd1 vssd1 vccd1 vccd1 _4495_/X sky130_fd_sc_hd__mux2_1
X_3446_ _5560_/B _3443_/A _5956_/B vssd1 vssd1 vccd1 vccd1 _5978_/A sky130_fd_sc_hd__a21o_2
XFILLER_0_85_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3377_ _3426_/B _3377_/B vssd1 vssd1 vccd1 vccd1 _3377_/Y sky130_fd_sc_hd__nor2_1
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4297__A4 _4287_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4151__B1 _3786_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6165_ _6181_/CLK _6165_/D vssd1 vssd1 vccd1 vccd1 _6165_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5116_ _5115_/A _5115_/B _3740_/Y vssd1 vssd1 vccd1 vccd1 _5116_/X sky130_fd_sc_hd__a21o_1
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6096_ _6354_/CLK _6096_/D vssd1 vssd1 vccd1 vccd1 _6096_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4067__A _6247_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5047_ _5929_/A1 _5046_/X _5034_/Y vssd1 vssd1 vccd1 vccd1 _5047_/X sky130_fd_sc_hd__a21bo_1
Xclkbuf_leaf_34_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6368_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__3402__C _4222_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5949_ _6396_/Q _5949_/B _5949_/C vssd1 vssd1 vccd1 vccd1 _5949_/X sky130_fd_sc_hd__and3b_1
XFILLER_0_47_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3146__A _4224_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3056__A _6242_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3300_ _3656_/A _5328_/B vssd1 vssd1 vccd1 vccd1 _5360_/C sky130_fd_sc_hd__nand2_2
XANTENNA__5970__S _5975_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4280_ _5599_/A _5349_/B vssd1 vssd1 vccd1 vccd1 _4281_/S sky130_fd_sc_hd__nor2_1
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3231_ _3183_/B _4744_/B _3573_/A _3143_/X vssd1 vssd1 vccd1 vccd1 _3231_/Y sky130_fd_sc_hd__a31oi_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3162_ _5256_/A _3369_/B vssd1 vssd1 vccd1 vccd1 _3572_/A sky130_fd_sc_hd__nor2_4
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3093_ _4744_/B _3232_/A vssd1 vssd1 vccd1 vccd1 _3194_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_89_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3222__C _3566_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xci2406_z80_185 vssd1 vssd1 vccd1 vccd1 ci2406_z80_185/HI io_oeb[3] sky130_fd_sc_hd__conb_1
Xci2406_z80_196 vssd1 vssd1 vccd1 vccd1 ci2406_z80_196/HI io_oeb[15] sky130_fd_sc_hd__conb_1
X_5803_ _6376_/Q _5849_/S _4864_/X vssd1 vssd1 vccd1 vccd1 _5803_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_76_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3995_ _3724_/A _6044_/A _4425_/A2 vssd1 vssd1 vccd1 vccd1 _3995_/Y sky130_fd_sc_hd__o21ai_1
X_5734_ _3039_/Y _4767_/B _3511_/D _5733_/X _3770_/A vssd1 vssd1 vccd1 vccd1 _5734_/X
+ sky130_fd_sc_hd__a32o_1
X_5665_ _5664_/X _5661_/X _4101_/X _4411_/X _5691_/S _5690_/S vssd1 vssd1 vccd1 vccd1
+ _5665_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_88_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4616_ _4616_/A _4616_/B vssd1 vssd1 vccd1 vccd1 _5372_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_4_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5596_ _5690_/S _4364_/X _5592_/X _5595_/X _5603_/D vssd1 vssd1 vccd1 vccd1 _5596_/X
+ sky130_fd_sc_hd__a221o_1
Xhold410 _5050_/X vssd1 vssd1 vccd1 vccd1 _6289_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6122__SET_B fanout180/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4547_ _3379_/B _3535_/D _5303_/A vssd1 vssd1 vccd1 vccd1 _4547_/Y sky130_fd_sc_hd__a21oi_1
Xhold432 _5955_/X vssd1 vssd1 vccd1 vccd1 _6400_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold421 _4593_/X vssd1 vssd1 vccd1 vccd1 _6246_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold454 _4525_/X vssd1 vssd1 vccd1 vccd1 _6226_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold443 _6231_/Q vssd1 vssd1 vccd1 vccd1 hold443/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold465 _4534_/X vssd1 vssd1 vccd1 vccd1 _6235_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold476 _6229_/Q vssd1 vssd1 vccd1 vccd1 hold476/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold487 _4524_/X vssd1 vssd1 vccd1 vccd1 _6225_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4478_ _4399_/X hold272/X _4482_/S vssd1 vssd1 vccd1 vccd1 _4478_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_96_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3429_ _3386_/B _3377_/B _4541_/B vssd1 vssd1 vccd1 vccd1 _3429_/X sky130_fd_sc_hd__o21a_1
Xhold498 _6433_/Q vssd1 vssd1 vccd1 vccd1 hold498/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4496__S _4500_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6217_ _6217_/CLK _6217_/D vssd1 vssd1 vccd1 vccd1 _6217_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4675__A1 _6245_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3478__A2 _5560_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6148_ _6413_/CLK hold62/X vssd1 vssd1 vccd1 vccd1 hold61/A sky130_fd_sc_hd__dfxtp_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6079_ _6368_/CLK _6079_/D fanout169/X vssd1 vssd1 vccd1 vccd1 _6079_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold423_A _6389_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6309__RESET_B fanout173/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4244__B _5725_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5927__A1 _6386_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5075__B _5075_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3323__B _4070_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3626__C1 _3047_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5091__A1 _3573_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5918__A1 _6385_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3780_ _3863_/A _3862_/S _3838_/S vssd1 vssd1 vccd1 vccd1 _4483_/A sky130_fd_sc_hd__or3_4
XFILLER_0_39_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4170__A _5217_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5450_ _5450_/A _5450_/B _5450_/C vssd1 vssd1 vccd1 vccd1 _5450_/X sky130_fd_sc_hd__and3_1
XANTENNA__5146__A2 _4255_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4401_ _4401_/A _4401_/B vssd1 vssd1 vccd1 vccd1 _5250_/B sky130_fd_sc_hd__xnor2_1
X_5381_ _5715_/A _6417_/Q vssd1 vssd1 vccd1 vccd1 _5383_/B sky130_fd_sc_hd__or2_1
X_4332_ hold252/X _4007_/X _4336_/S vssd1 vssd1 vccd1 vccd1 _4332_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_1_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4263_ _3254_/A _4247_/X _4262_/X _5952_/A vssd1 vssd1 vccd1 vccd1 _5603_/A sky130_fd_sc_hd__a22oi_4
XANTENNA__4106__B1 _3791_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3214_ _6257_/Q _6258_/Q _3334_/C vssd1 vssd1 vccd1 vccd1 _3566_/B sky130_fd_sc_hd__nand3b_4
XANTENNA__4657__A1 _5715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6002_ _6036_/A _6026_/B vssd1 vssd1 vccd1 vccd1 _6002_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_10_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3233__B _5258_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4194_ _3724_/A _6026_/A _4391_/A2 vssd1 vssd1 vccd1 vccd1 _4194_/Y sky130_fd_sc_hd__o21ai_1
X_3145_ _3116_/A _3144_/X _3193_/B vssd1 vssd1 vccd1 vccd1 _3177_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_82_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3076_ _6320_/Q vssd1 vssd1 vccd1 vccd1 _3076_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_89_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6402__RESET_B fanout178/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout161_A _5077_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6031__B1 _6063_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3978_ _6243_/Q _6244_/Q _6245_/Q _4073_/B vssd1 vssd1 vccd1 vccd1 _3978_/Y sky130_fd_sc_hd__a31oi_1
XFILLER_0_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5717_ _6268_/Q hold377/X _5723_/S vssd1 vssd1 vccd1 vccd1 _5717_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_72_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5137__A2 _6293_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5648_ _5648_/A _5648_/B vssd1 vssd1 vccd1 vccd1 _5648_/X sky130_fd_sc_hd__or2_1
X_5579_ _3654_/A _5323_/C _5578_/Y _4551_/Y _4347_/C vssd1 vssd1 vccd1 vccd1 _5579_/X
+ sky130_fd_sc_hd__a32o_1
Xhold240 _5961_/X vssd1 vssd1 vccd1 vccd1 _6408_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold251 _6133_/Q vssd1 vssd1 vccd1 vccd1 hold251/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold262 _4400_/X vssd1 vssd1 vccd1 vccd1 _6131_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold295 _5336_/X vssd1 vssd1 vccd1 vccd1 _6308_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold284 _6196_/Q vssd1 vssd1 vccd1 vccd1 hold284/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold273 _4478_/X vssd1 vssd1 vccd1 vccd1 _6179_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4648__A1 _6338_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3424__A _4309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4255__A _4541_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4887__A1 _6325_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3334__A _4284_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput8 io_in[28] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__clkbuf_2
Xclkbuf_2_0__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_6_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_59_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4165__A _5217_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4950_ _6328_/Q _5928_/A2 _5928_/B1 _4949_/X vssd1 vssd1 vccd1 vccd1 _4950_/X sky130_fd_sc_hd__a22o_1
X_3901_ _6295_/Q _4071_/C vssd1 vssd1 vccd1 vccd1 _4073_/B sky130_fd_sc_hd__nor2_1
X_4881_ _4880_/X _4879_/X _5053_/S vssd1 vssd1 vccd1 vccd1 _4882_/B sky130_fd_sc_hd__mux2_2
X_3832_ _4111_/A _4394_/B vssd1 vssd1 vccd1 vccd1 _3870_/A sky130_fd_sc_hd__nand2_1
X_3763_ _6242_/Q _3758_/Y _3761_/A _5216_/A vssd1 vssd1 vccd1 vccd1 _3763_/X sky130_fd_sc_hd__a22o_1
X_5502_ _5502_/A _5502_/B vssd1 vssd1 vccd1 vccd1 _5503_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_27_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3694_ _6310_/Q _5989_/B _4633_/D vssd1 vssd1 vccd1 vccd1 _4361_/B sky130_fd_sc_hd__or3_1
X_6482_ _6487_/A vssd1 vssd1 vccd1 vccd1 _6482_/X sky130_fd_sc_hd__buf_1
XFILLER_0_14_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5433_ hold606/X _5432_/X _5472_/S vssd1 vssd1 vccd1 vccd1 _5433_/X sky130_fd_sc_hd__mux2_1
X_5364_ _5553_/S _5364_/B vssd1 vssd1 vccd1 vccd1 _5471_/S sky130_fd_sc_hd__nand2_4
XANTENNA__3550__A1 _4685_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4973__S1 _5052_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4315_ _4316_/B _4315_/B vssd1 vssd1 vccd1 vccd1 _4315_/X sky130_fd_sc_hd__or2_1
X_5295_ hold624/X _3400_/B _5277_/Y _4228_/A vssd1 vssd1 vccd1 vccd1 _5295_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5827__A0 _6325_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4246_ hold1/X _4245_/X _5727_/S vssd1 vssd1 vccd1 vccd1 hold2/A sky130_fd_sc_hd__mux2_1
XFILLER_0_93_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3302__A1 _3337_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4177_ _4177_/A _4177_/B vssd1 vssd1 vccd1 vccd1 _4179_/B sky130_fd_sc_hd__nor2_1
X_3128_ _4685_/A _3334_/C _3290_/B vssd1 vssd1 vccd1 vccd1 _3193_/B sky130_fd_sc_hd__or3_2
XANTENNA__5055__A1 _6274_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3059_ _6247_/Q vssd1 vssd1 vccd1 vccd1 _4075_/A sky130_fd_sc_hd__inv_2
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_42_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_37_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4404__S0 _5676_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4955__S1 _5052_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3064__A _6292_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5080_ hold490/X _4520_/Y _5079_/X vssd1 vssd1 vccd1 vccd1 _5080_/Y sky130_fd_sc_hd__o21ai_1
X_4100_ hold27/X _4425_/A2 _5597_/B vssd1 vssd1 vccd1 vccd1 _4100_/X sky130_fd_sc_hd__o21a_1
XANTENNA__5285__B2 _5560_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4031_ _6246_/Q _4031_/B _4031_/C vssd1 vssd1 vccd1 vccd1 _4032_/B sky130_fd_sc_hd__or3_1
XFILLER_0_47_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4088__A2 _6052_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5982_ _5981_/X _3577_/A _5982_/S vssd1 vssd1 vccd1 vccd1 _6425_/D sky130_fd_sc_hd__mux2_1
X_4933_ hold397/X _4932_/X _5557_/S vssd1 vssd1 vccd1 vccd1 _4933_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_19_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4623__A input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_13 _4347_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4864_ _6324_/Q _4752_/X _4751_/B vssd1 vssd1 vccd1 vccd1 _4864_/X sky130_fd_sc_hd__a21o_1
X_4795_ _6417_/Q _4758_/X _4789_/X _4793_/X _4794_/X vssd1 vssd1 vccd1 vccd1 _4795_/X
+ sky130_fd_sc_hd__a2111o_1
X_3815_ _6133_/Q _3789_/X _3791_/X _6412_/Q vssd1 vssd1 vccd1 vccd1 _3815_/X sky130_fd_sc_hd__a22o_1
X_3746_ _3755_/C _3747_/B vssd1 vssd1 vccd1 vccd1 _3746_/X sky130_fd_sc_hd__and2_4
XANTENNA_fanout124_A _4214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3677_ _4270_/B _3676_/X _5097_/B vssd1 vssd1 vccd1 vccd1 _3677_/Y sky130_fd_sc_hd__o21ai_1
X_5416_ hold608/X input3/X _5469_/S vssd1 vssd1 vccd1 vccd1 _5416_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_2_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6396_ _6397_/CLK _6396_/D fanout173/X vssd1 vssd1 vccd1 vccd1 _6396_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_9_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_100_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5347_ _5347_/A _5347_/B vssd1 vssd1 vccd1 vccd1 _5347_/Y sky130_fd_sc_hd__nor2_1
X_5278_ _3572_/A _3581_/A _5266_/C _5266_/D vssd1 vssd1 vccd1 vccd1 _5278_/X sky130_fd_sc_hd__a211o_1
X_4229_ _4541_/D _3553_/Y _4228_/Y _4209_/Y vssd1 vssd1 vccd1 vccd1 _4229_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_84_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3762__A1 _6340_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5364__A _5553_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5258__B _5258_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput11 io_in[31] vssd1 vssd1 vccd1 vccd1 _3082_/A sky130_fd_sc_hd__buf_1
XANTENNA__3059__A _6247_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3600_ _3600_/A _3600_/B _3600_/C _5272_/B vssd1 vssd1 vccd1 vccd1 _5327_/A sky130_fd_sc_hd__or4_1
XFILLER_0_71_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5973__S _5975_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4580_ _6418_/Q _4569_/X _4570_/X _6269_/Q vssd1 vssd1 vccd1 vccd1 _4580_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3753__A1 _4679_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3531_ _5560_/B hold289/X _3403_/B _3528_/Y _3530_/X vssd1 vssd1 vccd1 vccd1 _3531_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_12_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4589__S _4604_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6250_ _6401_/CLK _6250_/D fanout179/X vssd1 vssd1 vccd1 vccd1 _6250_/Q sky130_fd_sc_hd__dfrtp_1
X_3462_ hold31/X _3507_/B hold47/X _3507_/C vssd1 vssd1 vccd1 vccd1 _3462_/X sky130_fd_sc_hd__or4_1
X_3393_ _3384_/Y _3387_/X _3391_/A _5270_/A _3392_/Y vssd1 vssd1 vccd1 vccd1 _3394_/D
+ sky130_fd_sc_hd__a221o_1
X_5201_ _3905_/X _5178_/A _5195_/X _5200_/Y vssd1 vssd1 vccd1 vccd1 _5201_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_58_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6181_ _6181_/CLK _6181_/D vssd1 vssd1 vccd1 vccd1 _6181_/Q sky130_fd_sc_hd__dfxtp_1
X_5132_ _5211_/C _5211_/D vssd1 vssd1 vccd1 vccd1 _5133_/B sky130_fd_sc_hd__xor2_1
XANTENNA__3269__B1 _5560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5063_ _6367_/Q _5062_/X _5927_/S vssd1 vssd1 vccd1 vccd1 _5063_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3808__A2 _3789_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4014_ hold212/X _3784_/X _3786_/X hold235/X _4013_/X vssd1 vssd1 vccd1 vccd1 _4017_/A
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4233__A2 _5733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5430__A1 input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5965_ _4412_/X hold291/X _5967_/S vssd1 vssd1 vccd1 vccd1 _6412_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_90_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5896_ _6420_/Q _5895_/X _5930_/S vssd1 vssd1 vccd1 vccd1 _5896_/X sky130_fd_sc_hd__mux2_1
X_4916_ hold346/X _4915_/X _4916_/S vssd1 vssd1 vccd1 vccd1 _4916_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_90_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4847_ _4866_/B _4867_/B _4847_/C vssd1 vssd1 vccd1 vccd1 _4852_/A sky130_fd_sc_hd__and3b_1
XFILLER_0_74_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5883__S _5931_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4941__A0 _6380_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4778_ _6319_/Q _4777_/X _5849_/S vssd1 vssd1 vccd1 vccd1 _4778_/X sky130_fd_sc_hd__mux2_1
X_3729_ _6303_/Q _3755_/C vssd1 vssd1 vccd1 vccd1 _5087_/B sky130_fd_sc_hd__and2_2
XANTENNA__4499__S _4500_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6448_ _6448_/CLK _6448_/D fanout181/X vssd1 vssd1 vccd1 vccd1 _6448_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_0_100_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6379_ _6383_/CLK _6379_/D fanout168/X vssd1 vssd1 vccd1 vccd1 _6379_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_100_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4247__B _5313_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4962__S _5058_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5421__A1 _4843_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3983__A1 _6343_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4932__A0 _6416_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_4_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6407_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_0_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5032__S0 _5051_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5488__A1 _4938_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5033__S _5053_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5968__S _5975_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4215__A2 _5715_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5750_ _6319_/Q _5728_/D _4742_/X _5749_/X vssd1 vssd1 vccd1 vccd1 _5750_/X sky130_fd_sc_hd__a22o_1
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5681_ hold414/X _5588_/X _5594_/Y _5678_/X vssd1 vssd1 vccd1 vccd1 _5681_/X sky130_fd_sc_hd__a22o_1
X_4701_ _3960_/Y _4700_/X _4731_/S vssd1 vssd1 vccd1 vccd1 _4701_/X sky130_fd_sc_hd__mux2_1
X_4632_ hold624/X _4615_/X _4617_/Y _4631_/X vssd1 vssd1 vccd1 vccd1 _4632_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_60_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4923__A0 _6379_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4563_ _4568_/C _4570_/B vssd1 vssd1 vccd1 vccd1 _4564_/A sky130_fd_sc_hd__nor2_4
Xhold603 _6380_/Q vssd1 vssd1 vccd1 vccd1 _5856_/A sky130_fd_sc_hd__buf_1
XFILLER_0_4_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6302_ _6403_/CLK _6302_/D fanout179/X vssd1 vssd1 vccd1 vccd1 _6302_/Q sky130_fd_sc_hd__dfrtp_1
Xhold625 _4632_/X vssd1 vssd1 vccd1 vccd1 _6258_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold636 _5287_/X vssd1 vssd1 vccd1 vccd1 _6301_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3514_ hold118/X _3513_/X _5472_/S vssd1 vssd1 vccd1 vccd1 _3514_/X sky130_fd_sc_hd__mux2_1
Xhold614 _6116_/Q vssd1 vssd1 vccd1 vccd1 hold614/X sky130_fd_sc_hd__buf_1
X_4494_ _3923_/X hold238/X _4500_/S vssd1 vssd1 vccd1 vccd1 _6193_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_100_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3445_ _3473_/B _3473_/A vssd1 vssd1 vccd1 vccd1 _5956_/B sky130_fd_sc_hd__and2b_2
X_6233_ _6270_/CLK _6233_/D fanout176/X vssd1 vssd1 vccd1 vccd1 _6233_/Q sky130_fd_sc_hd__dfstp_1
Xhold669 _6292_/Q vssd1 vssd1 vccd1 vccd1 hold669/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold658 _6272_/Q vssd1 vssd1 vccd1 vccd1 hold658/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold647 _6273_/Q vssd1 vssd1 vccd1 vccd1 hold647/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5479__A1 _4313_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6080__RESET_B fanout169/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3376_ _5322_/C _3376_/B _5326_/B _5272_/A vssd1 vssd1 vccd1 vccd1 _3377_/B sky130_fd_sc_hd__or4_1
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6164_ _6412_/CLK _6164_/D vssd1 vssd1 vccd1 vccd1 _6164_/Q sky130_fd_sc_hd__dfxtp_1
X_5115_ _5115_/A _5115_/B vssd1 vssd1 vccd1 vccd1 _5115_/Y sky130_fd_sc_hd__nor2_1
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6095_ _6218_/CLK _6095_/D vssd1 vssd1 vccd1 vccd1 _6095_/Q sky130_fd_sc_hd__dfxtp_1
X_5046_ _6333_/Q _5928_/A2 _5928_/B1 _5045_/X vssd1 vssd1 vccd1 vccd1 _5046_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5948_ _3621_/A _3625_/B hold545/X _3623_/A _3466_/B vssd1 vssd1 vccd1 vccd1 _5948_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_90_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5879_ _6363_/Q _6382_/Q _5927_/S vssd1 vssd1 vccd1 vccd1 _5879_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_35_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5167__B1 _5243_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4914__A0 _6326_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3146__B _3278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4957__S _5053_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5014__S0 _5358_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5890__A1 _6379_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6433__SET_B fanout171/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3708__A1 _3473_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3337__A _3337_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3230_ _3549_/A _3152_/Y _4679_/D _3566_/B _3525_/B vssd1 vssd1 vccd1 vccd1 _3230_/X
+ sky130_fd_sc_hd__o32a_1
XANTENNA__4133__A1 _6292_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5330__A0 _4214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3161_ _3289_/A _3534_/A vssd1 vssd1 vccd1 vccd1 _3369_/B sky130_fd_sc_hd__or2_4
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3092_ _4744_/A _3183_/B vssd1 vssd1 vccd1 vccd1 _3232_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_55_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xci2406_z80_186 vssd1 vssd1 vccd1 vccd1 ci2406_z80_186/HI io_oeb[5] sky130_fd_sc_hd__conb_1
Xci2406_z80_197 vssd1 vssd1 vccd1 vccd1 ci2406_z80_197/HI io_oeb[16] sky130_fd_sc_hd__conb_1
X_5802_ _5791_/A _5742_/A _5801_/X _5731_/X vssd1 vssd1 vccd1 vccd1 _5802_/X sky130_fd_sc_hd__o22a_1
X_3994_ _6044_/A vssd1 vssd1 vccd1 vccd1 _3994_/Y sky130_fd_sc_hd__inv_2
X_5733_ _5733_/A _5733_/B _5360_/X vssd1 vssd1 vccd1 vccd1 _5733_/X sky130_fd_sc_hd__or3b_1
XFILLER_0_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4631__A input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5664_ _5664_/A _5664_/B vssd1 vssd1 vccd1 vccd1 _5664_/X sky130_fd_sc_hd__or2_1
X_4615_ _4615_/A _4615_/B vssd1 vssd1 vccd1 vccd1 _4615_/X sky130_fd_sc_hd__and2_4
X_5595_ _6314_/Q _5597_/B _5595_/C vssd1 vssd1 vccd1 vccd1 _5595_/X sky130_fd_sc_hd__and3_1
XFILLER_0_32_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6261__RESET_B fanout177/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4546_ _4568_/C _4567_/B _5339_/A vssd1 vssd1 vccd1 vccd1 _4546_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_0_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold411 _6444_/Q vssd1 vssd1 vccd1 vccd1 hold411/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold400 _6049_/X vssd1 vssd1 vccd1 vccd1 _6445_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold422 _6426_/Q vssd1 vssd1 vccd1 vccd1 hold422/X sky130_fd_sc_hd__clkbuf_2
Xhold444 _4530_/X vssd1 vssd1 vccd1 vccd1 _6231_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold433 _6314_/Q vssd1 vssd1 vccd1 vccd1 hold433/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold466 _6230_/Q vssd1 vssd1 vccd1 vccd1 hold466/X sky130_fd_sc_hd__dlygate4sd3_1
X_4477_ _4392_/X hold155/X _4482_/S vssd1 vssd1 vccd1 vccd1 _4477_/X sky130_fd_sc_hd__mux2_1
Xhold477 _4528_/X vssd1 vssd1 vccd1 vccd1 _6229_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold455 _6436_/Q vssd1 vssd1 vccd1 vccd1 hold455/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3428_ _3386_/B _4734_/B _3384_/Y _5292_/C _3426_/X vssd1 vssd1 vccd1 vccd1 _3428_/X
+ sky130_fd_sc_hd__a221o_1
Xhold488 _6228_/Q vssd1 vssd1 vccd1 vccd1 hold488/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold499 _5999_/X vssd1 vssd1 vccd1 vccd1 _6433_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6216_ _6217_/CLK _6216_/D vssd1 vssd1 vccd1 vccd1 _6216_/Q sky130_fd_sc_hd__dfxtp_1
X_3359_ _5313_/A _3359_/B _3359_/C vssd1 vssd1 vccd1 vccd1 _4757_/B sky130_fd_sc_hd__or3_4
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6147_ _6413_/CLK hold60/X vssd1 vssd1 vccd1 vccd1 hold59/A sky130_fd_sc_hd__dfxtp_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6078_ _6368_/CLK _6078_/D fanout169/X vssd1 vssd1 vccd1 vccd1 _6078_/Q sky130_fd_sc_hd__dfrtp_2
X_5029_ _6365_/Q _5028_/X _5029_/S vssd1 vssd1 vccd1 vccd1 _5029_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_82_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5372__A _5739_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3626__B1 _3639_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3620__A _5935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5091__A2 _5217_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4170__B _6248_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3067__A _6416_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4400_ hold261/X _4399_/X _4428_/S vssd1 vssd1 vccd1 vccd1 _4400_/X sky130_fd_sc_hd__mux2_1
X_5380_ _5518_/S _5380_/B _5380_/C vssd1 vssd1 vccd1 vccd1 _5450_/A sky130_fd_sc_hd__or3_4
XFILLER_0_22_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4331_ hold216/X _3965_/X _4336_/S vssd1 vssd1 vccd1 vccd1 _4331_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_22_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4262_ _3530_/D _4254_/X _4256_/X _4261_/X _5584_/A1 vssd1 vssd1 vccd1 vccd1 _4262_/X
+ sky130_fd_sc_hd__a32o_1
X_3213_ _4228_/A _3534_/A vssd1 vssd1 vccd1 vccd1 _3215_/C sky130_fd_sc_hd__nand2_1
X_6001_ _5560_/D _6000_/X _6026_/B vssd1 vssd1 vccd1 vccd1 _6001_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_5_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4193_ _6026_/A vssd1 vssd1 vccd1 vccd1 _4193_/Y sky130_fd_sc_hd__inv_2
X_3144_ _3534_/A _3121_/Y _3143_/X vssd1 vssd1 vccd1 vccd1 _3144_/X sky130_fd_sc_hd__o21ba_1
XANTENNA__5606__A1 _4070_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3075_ _6272_/Q vssd1 vssd1 vccd1 vccd1 _3075_/Y sky130_fd_sc_hd__inv_2
XANTENNA__5606__B2 _6267_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_32_wb_clk_i_A clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_82_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6031__A1 _4313_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3977_ _6243_/Q _6244_/Q _6245_/Q vssd1 vssd1 vccd1 vccd1 _4073_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_64_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5457__A _5560_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5790__B1 _5735_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5716_ _6267_/Q hold397/X _5723_/S vssd1 vssd1 vccd1 vccd1 _5716_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4593__A1 _5695_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3148__A2 _3278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5647_ _6132_/Q _4198_/B _5676_/B1 _6211_/Q _5676_/C1 vssd1 vssd1 vccd1 vccd1 _5648_/B
+ sky130_fd_sc_hd__o221a_1
XANTENNA__3408__C _6390_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5578_ _5578_/A _5578_/B vssd1 vssd1 vccd1 vccd1 _5578_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_13_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4529_ hold466/X _6272_/Q _4539_/S vssd1 vssd1 vccd1 vccd1 _4529_/X sky130_fd_sc_hd__mux2_1
Xhold241 _6175_/Q vssd1 vssd1 vccd1 vccd1 hold241/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold230 _4433_/X vssd1 vssd1 vccd1 vccd1 _6139_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold252 _6094_/Q vssd1 vssd1 vccd1 vccd1 hold252/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold274 _6185_/Q vssd1 vssd1 vccd1 vccd1 hold274/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold296 _6073_/Q vssd1 vssd1 vccd1 vccd1 hold296/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold263 _6197_/Q vssd1 vssd1 vccd1 vccd1 hold263/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold285 _6163_/Q vssd1 vssd1 vccd1 vccd1 hold285/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5073__A2 _5247_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4255__B _4255_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4820__A2 _5728_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3615__A _4541_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3334__B _5226_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3311__A2 _3309_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput9 io_in[29] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__4165__B _6343_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3900_ _6243_/Q _6244_/Q _6245_/Q vssd1 vssd1 vccd1 vccd1 _4066_/B sky130_fd_sc_hd__o21ai_2
XFILLER_0_59_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6013__A1 _4313_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4880_ hold89/A hold81/A _6413_/Q _6182_/Q _5358_/A0 _4326_/B vssd1 vssd1 vccd1 vccd1
+ _4880_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_52_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3831_ _3831_/A _3831_/B _3831_/C vssd1 vssd1 vccd1 vccd1 _4394_/B sky130_fd_sc_hd__or3_4
X_3762_ _6336_/Q _6340_/Q _6301_/Q vssd1 vssd1 vccd1 vccd1 _5216_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_6_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5501_ _5554_/A _5501_/B vssd1 vssd1 vccd1 vccd1 _5502_/B sky130_fd_sc_hd__nor2_1
X_3693_ _6308_/Q _6309_/Q vssd1 vssd1 vccd1 vccd1 _4633_/D sky130_fd_sc_hd__and2_1
X_6481_ _6487_/A vssd1 vssd1 vccd1 vccd1 _6481_/X sky130_fd_sc_hd__buf_1
X_5432_ _6420_/Q _5431_/X _5471_/S vssd1 vssd1 vccd1 vccd1 _5432_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4327__A1 _5339_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5363_ _4214_/A _4639_/B _5359_/X _5362_/X _4767_/A vssd1 vssd1 vccd1 vccd1 _5364_/B
+ sky130_fd_sc_hd__a32o_1
XANTENNA__3550__A2 _5096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4314_ _4310_/C _4313_/Y _4314_/S vssd1 vssd1 vccd1 vccd1 _4315_/B sky130_fd_sc_hd__mux2_1
X_5294_ _5294_/A _5294_/B _5294_/C _5294_/D vssd1 vssd1 vccd1 vccd1 _5294_/X sky130_fd_sc_hd__or4_1
XFILLER_0_10_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5740__A _5740_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4245_ _6317_/Q _6335_/Q _4245_/S vssd1 vssd1 vccd1 vccd1 _4245_/X sky130_fd_sc_hd__mux2_1
X_4176_ _4176_/A _4176_/B vssd1 vssd1 vccd1 vccd1 _4178_/A sky130_fd_sc_hd__nand2_1
X_3127_ _4228_/A _3594_/A _4214_/B vssd1 vssd1 vccd1 vccd1 _3194_/B sky130_fd_sc_hd__and3_1
XFILLER_0_89_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3058_ _6246_/Q vssd1 vssd1 vccd1 vccd1 _4066_/A sky130_fd_sc_hd__inv_2
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4802__A2 _4313_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4015__B1 _3791_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3526__C1 _5560_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3829__B1 _3791_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6481__A _6487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4101__S0 _5676_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3517__C1 _4214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4404__S1 _5676_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3345__A _5560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3296__A1 _5578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4030_ _4031_/B _4031_/C _6246_/Q vssd1 vssd1 vccd1 vccd1 _4059_/A sky130_fd_sc_hd__o21ai_2
XANTENNA__5560__A _5560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5981_ _5981_/A _5981_/B vssd1 vssd1 vccd1 vccd1 _5981_/X sky130_fd_sc_hd__or2_1
XFILLER_0_47_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4932_ _6416_/Q _4931_/X _5930_/S vssd1 vssd1 vccd1 vccd1 _4932_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5993__B1 _4313_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4904__A _6323_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4623__B _4631_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4863_ _5054_/A _4863_/B vssd1 vssd1 vccd1 vccd1 _4863_/Y sky130_fd_sc_hd__nand2_1
X_3814_ _6189_/Q _3779_/X _3781_/X hold49/A _3813_/X vssd1 vssd1 vccd1 vccd1 _3817_/A
+ sky130_fd_sc_hd__a221o_1
X_4794_ _6434_/Q _4756_/Y _4757_/Y _4788_/B _4754_/X vssd1 vssd1 vccd1 vccd1 _4794_/X
+ sky130_fd_sc_hd__a221o_1
X_3745_ _6303_/Q _3938_/A _6304_/Q vssd1 vssd1 vccd1 vccd1 _3747_/B sky130_fd_sc_hd__and3b_1
XFILLER_0_42_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3676_ _3254_/A _5578_/A _3566_/B _3136_/B _3289_/A vssd1 vssd1 vccd1 vccd1 _3676_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_88_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5415_ _5441_/A _5414_/X _5371_/A vssd1 vssd1 vccd1 vccd1 _5415_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_88_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3255__A _3278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6395_ _6397_/CLK _6395_/D fanout172/X vssd1 vssd1 vccd1 vccd1 _6395_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_28_wb_clk_i _6404_/CLK vssd1 vssd1 vccd1 vccd1 _6421_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_23_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3523__A2 _3164_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5346_ _4633_/B _5345_/X _5727_/S vssd1 vssd1 vccd1 vccd1 _6311_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_2_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5277_ _3337_/A _3502_/A _3400_/B vssd1 vssd1 vccd1 vccd1 _5277_/Y sky130_fd_sc_hd__a21oi_1
X_4228_ _4228_/A _4541_/A vssd1 vssd1 vccd1 vccd1 _4228_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_97_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4159_ _4121_/A _4121_/B _4122_/B vssd1 vssd1 vccd1 vccd1 _4160_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_92_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5736__B1 _5935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4539__A1 _6298_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4398__S0 _5673_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4695__S _4731_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5267__A2 _3770_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5380__A _5518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5672__C1 _3721_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5975__A0 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput12 io_in[35] vssd1 vssd1 vccd1 vccd1 _3083_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__3753__A2 _6243_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3530_ _5560_/B _5360_/C _4228_/A _3530_/D vssd1 vssd1 vccd1 vccd1 _3530_/X sky130_fd_sc_hd__and4bb_1
XFILLER_0_3_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3461_ _3507_/C _3449_/X _3465_/B vssd1 vssd1 vccd1 vccd1 _3461_/X sky130_fd_sc_hd__a21o_1
XANTENNA__3075__A _6272_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3392_ _3337_/A _4747_/D _3297_/X _3581_/B _3654_/A vssd1 vssd1 vccd1 vccd1 _3392_/Y
+ sky130_fd_sc_hd__o32ai_4
X_5200_ _5102_/B _5199_/Y _5178_/A vssd1 vssd1 vccd1 vccd1 _5200_/Y sky130_fd_sc_hd__a21oi_1
X_6180_ _6410_/CLK _6180_/D vssd1 vssd1 vccd1 vccd1 _6180_/Q sky130_fd_sc_hd__dfxtp_1
X_5131_ _5211_/A _5211_/B vssd1 vssd1 vccd1 vccd1 _5133_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_58_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5062_ _6386_/Q _4754_/X _5056_/X _5061_/X vssd1 vssd1 vccd1 vccd1 _5062_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_42_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3269__A1 _4309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5663__C1 _5673_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4013_ _6112_/Q _3779_/X _3781_/X hold77/A vssd1 vssd1 vccd1 vccd1 _4013_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_79_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4233__A3 _3770_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5964_ _4405_/X hold300/X _5967_/S vssd1 vssd1 vccd1 vccd1 _6411_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_90_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3441__A1 _3047_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5895_ _5929_/A1 _5894_/X _4996_/Y vssd1 vssd1 vccd1 vccd1 _5895_/X sky130_fd_sc_hd__a21bo_1
X_4915_ hold157/X _4914_/X _5029_/S vssd1 vssd1 vccd1 vccd1 _4915_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5718__A0 _6269_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4846_ _6323_/Q _4846_/B vssd1 vssd1 vccd1 vccd1 _4866_/B sky130_fd_sc_hd__and2_1
XFILLER_0_62_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3744__A2 _6242_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4777_ _6371_/Q _4754_/X _4760_/X _4776_/X vssd1 vssd1 vccd1 vccd1 _4777_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_7_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6060__S _6060_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3728_ _6304_/Q _5196_/S vssd1 vssd1 vccd1 vccd1 _4040_/A sky130_fd_sc_hd__nand2_4
XFILLER_0_70_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3659_ _3657_/A _3657_/B _3658_/Y vssd1 vssd1 vccd1 vccd1 _3659_/X sky130_fd_sc_hd__a21o_1
X_6447_ _6447_/CLK _6447_/D fanout168/X vssd1 vssd1 vccd1 vccd1 _6447_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_0_30_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6378_ _6383_/CLK _6378_/D fanout168/X vssd1 vssd1 vccd1 vccd1 _6378_/Q sky130_fd_sc_hd__dfrtp_4
X_5329_ _4224_/A _5270_/B _4734_/B _5328_/X vssd1 vssd1 vccd1 vccd1 _5329_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_11_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3680__A1 _5096_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5957__B1 _3443_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4544__A _5339_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_hold613_A _6295_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_2_3__f_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5032__S1 _5052_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5660__A2 _4198_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3671__B2 _3164_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4620__B1 _4617_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4700_ _4697_/X _4699_/X _5240_/S vssd1 vssd1 vccd1 vccd1 _4700_/X sky130_fd_sc_hd__mux2_1
X_5680_ _6297_/Q _5587_/X _5610_/X _6447_/Q _5679_/X vssd1 vssd1 vccd1 vccd1 _5683_/A
+ sky130_fd_sc_hd__a221o_1
X_4631_ input7/X _4631_/B vssd1 vssd1 vccd1 vccd1 _4631_/X sky130_fd_sc_hd__and2_1
XANTENNA__5176__A1 _6294_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4562_ _5725_/A _4568_/B vssd1 vssd1 vccd1 vccd1 _4570_/B sky130_fd_sc_hd__nor2_2
Xhold626 _6303_/Q vssd1 vssd1 vccd1 vccd1 hold626/X sky130_fd_sc_hd__dlygate4sd3_1
X_6301_ _6305_/CLK _6301_/D fanout179/X vssd1 vssd1 vccd1 vccd1 _6301_/Q sky130_fd_sc_hd__dfrtp_4
X_3513_ _4767_/A _3511_/X _3512_/Y vssd1 vssd1 vccd1 vccd1 _3513_/X sky130_fd_sc_hd__a21bo_1
Xhold615 _3493_/X vssd1 vssd1 vccd1 vccd1 _6116_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold604 _5864_/X vssd1 vssd1 vccd1 vccd1 _6380_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4493_ _3881_/X hold292/X _4500_/S vssd1 vssd1 vccd1 vccd1 _4493_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_40_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold659 _6252_/Q vssd1 vssd1 vccd1 vccd1 hold659/X sky130_fd_sc_hd__buf_1
X_3444_ _4901_/S _3622_/A vssd1 vssd1 vccd1 vccd1 _3469_/A sky130_fd_sc_hd__or2_1
Xhold637 _6416_/Q vssd1 vssd1 vccd1 vccd1 hold637/X sky130_fd_sc_hd__dlygate4sd3_1
X_6232_ _6343_/CLK _6232_/D fanout170/X vssd1 vssd1 vccd1 vccd1 _6232_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA__5479__A2 _5377_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold648 _6269_/Q vssd1 vssd1 vccd1 vccd1 hold648/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4687__B1 _4731_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4629__A input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3375_ _5733_/A _5481_/A _5324_/B _5481_/B vssd1 vssd1 vccd1 vccd1 _5272_/A sky130_fd_sc_hd__or4_1
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4151__A2 _3784_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6163_ _6410_/CLK _6163_/D vssd1 vssd1 vccd1 vccd1 _6163_/Q sky130_fd_sc_hd__dfxtp_1
X_5114_ _5114_/A _5114_/B vssd1 vssd1 vccd1 vccd1 _5115_/B sky130_fd_sc_hd__xnor2_1
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6094_ _6218_/CLK _6094_/D vssd1 vssd1 vccd1 vccd1 _6094_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3252__B _3725_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5636__C1 _5675_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5045_ _6366_/Q _5044_/X _5927_/S vssd1 vssd1 vccd1 vccd1 _5045_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_79_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5547__A2_N _5377_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5947_ _5952_/A _3043_/A _5949_/B _5936_/Y vssd1 vssd1 vccd1 vccd1 _5947_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_47_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5878_ _5889_/B _5878_/B vssd1 vssd1 vccd1 vccd1 _5878_/Y sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_43_wb_clk_i clkbuf_leaf_6_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6445_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_4829_ _6374_/Q _6322_/Q _4901_/S vssd1 vssd1 vccd1 vccd1 _4829_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_62_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5989__D_N _4633_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5014__S1 _4326_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3443__A _3443_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5890__A2 _6380_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3162__B _3369_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5833__A _6378_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4669__A0 _6338_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3160_ _3289_/A _3289_/C _4222_/B vssd1 vssd1 vccd1 vccd1 _5317_/A sky130_fd_sc_hd__and3_2
XANTENNA__5271__C _5322_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3091_ _3525_/B _3334_/C _6258_/Q _6257_/Q vssd1 vssd1 vccd1 vccd1 _3091_/X sky130_fd_sc_hd__or4bb_2
Xhold1 hold1/A vssd1 vssd1 vccd1 vccd1 hold1/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_22_wb_clk_i_A _6404_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5633__A2 _4382_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3644__A1 _3048_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xci2406_z80_187 vssd1 vssd1 vccd1 vccd1 ci2406_z80_187/HI io_oeb[6] sky130_fd_sc_hd__conb_1
X_5801_ _5815_/S _5796_/X _5800_/X _5747_/A vssd1 vssd1 vccd1 vccd1 _5801_/X sky130_fd_sc_hd__o22a_1
X_5732_ _3109_/B _5270_/B _3373_/B _3579_/B _4214_/A vssd1 vssd1 vccd1 vccd1 _5733_/B
+ sky130_fd_sc_hd__o41a_1
X_3993_ _4142_/S _3991_/X _3992_/X vssd1 vssd1 vccd1 vccd1 _6044_/A sky130_fd_sc_hd__a21oi_4
Xci2406_z80_198 vssd1 vssd1 vccd1 vccd1 ci2406_z80_198/HI io_oeb[17] sky130_fd_sc_hd__conb_1
XFILLER_0_29_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4631__B _4631_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3528__A _5560_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5663_ _6096_/Q _4382_/B _4200_/S _6141_/Q _5673_/C1 vssd1 vssd1 vccd1 vccd1 _5664_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_29_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4614_ hold587/X _5313_/A _5740_/A vssd1 vssd1 vccd1 vccd1 _4615_/B sky130_fd_sc_hd__a21o_1
X_5594_ _5599_/A _5603_/B _5603_/C vssd1 vssd1 vccd1 vccd1 _5594_/Y sky130_fd_sc_hd__a21oi_4
X_4545_ _5725_/A _4568_/B vssd1 vssd1 vccd1 vccd1 _4567_/B sky130_fd_sc_hd__nand2_2
XANTENNA__4372__A2 _4382_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold401 _6287_/Q vssd1 vssd1 vccd1 vccd1 hold401/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold423 _6389_/Q vssd1 vssd1 vccd1 vccd1 _3457_/A sky130_fd_sc_hd__buf_1
Xhold434 _5351_/X vssd1 vssd1 vccd1 vccd1 _6314_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold445 _6232_/Q vssd1 vssd1 vccd1 vccd1 hold445/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold412 _6045_/X vssd1 vssd1 vccd1 vccd1 _6444_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold478 _6238_/Q vssd1 vssd1 vccd1 vccd1 hold478/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold467 _4529_/X vssd1 vssd1 vccd1 vccd1 _6230_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold456 _6011_/X vssd1 vssd1 vccd1 vccd1 _6436_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4476_ _4380_/X hold115/X _4482_/S vssd1 vssd1 vccd1 vccd1 _4476_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_96_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3427_ _5325_/A _3427_/B vssd1 vssd1 vccd1 vccd1 _5292_/C sky130_fd_sc_hd__nand2_1
Xhold489 _4527_/X vssd1 vssd1 vccd1 vccd1 _6228_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6215_ _6354_/CLK _6215_/D vssd1 vssd1 vccd1 vccd1 _6215_/Q sky130_fd_sc_hd__dfxtp_1
X_3358_ _3257_/X _3356_/Y _3357_/X _3349_/X vssd1 vssd1 vccd1 vccd1 _3359_/C sky130_fd_sc_hd__o31a_1
X_6146_ _6209_/CLK hold56/X vssd1 vssd1 vccd1 vccd1 hold55/A sky130_fd_sc_hd__dfxtp_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3289_ _3289_/A _4214_/B _3289_/C vssd1 vssd1 vccd1 vccd1 _3657_/A sky130_fd_sc_hd__and3_2
X_6077_ _6351_/CLK _6077_/D vssd1 vssd1 vccd1 vccd1 _6077_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5624__A2 _4198_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5028_ _6421_/Q _5027_/X _5930_/S vssd1 vssd1 vccd1 vccd1 _5028_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_67_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5388__B2 _5441_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4541__B _4541_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold409_A _6289_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4994__S0 _5051_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5312__B2 _5578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3901__A _6295_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6484__A _6487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3626__A1 _6415_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5379__A1 _5472_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3562__B1 _5096_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4330_ hold199/X _3923_/X _4336_/S vssd1 vssd1 vccd1 vccd1 _4330_/X sky130_fd_sc_hd__mux2_1
X_4261_ _3226_/Y _3654_/A _4259_/X _4228_/A _4260_/X vssd1 vssd1 vccd1 vccd1 _4261_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4106__A2 _3789_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3212_ _3122_/X _3148_/X _3211_/X _3241_/B _3208_/X vssd1 vssd1 vccd1 vccd1 _3212_/X
+ sky130_fd_sc_hd__a32o_1
X_6000_ _6057_/B _4788_/B _5387_/Y _5992_/Y vssd1 vssd1 vccd1 vccd1 _6000_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_5_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4192_ _4142_/S _4191_/X _4158_/X vssd1 vssd1 vccd1 vccd1 _6026_/A sky130_fd_sc_hd__a21oi_4
XFILLER_0_66_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3143_ _3289_/A _6254_/Q _3289_/C vssd1 vssd1 vccd1 vccd1 _3143_/X sky130_fd_sc_hd__and3_1
X_3074_ _6270_/Q vssd1 vssd1 vccd1 vccd1 _3074_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_82_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3976_ _5087_/A _6245_/Q _6339_/Q _3740_/Y _3975_/X vssd1 vssd1 vccd1 vccd1 _5205_/B
+ sky130_fd_sc_hd__o41a_2
XFILLER_0_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5715_ _5715_/A _5715_/B _5715_/C _5226_/C vssd1 vssd1 vccd1 vccd1 _5723_/S sky130_fd_sc_hd__or4b_4
XANTENNA__5790__A1 _5236_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3258__A _5096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5646_ _6411_/Q _4198_/B _5676_/B1 _6180_/Q _5675_/C1 vssd1 vssd1 vccd1 vccd1 _5648_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_33_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5577_ _3418_/A _3337_/B _4248_/Y _4268_/B vssd1 vssd1 vccd1 vccd1 _5577_/X sky130_fd_sc_hd__o211a_1
Xhold220 _6138_/Q vssd1 vssd1 vccd1 vccd1 hold220/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold242 _4473_/X vssd1 vssd1 vccd1 vccd1 _6175_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4528_ hold476/X _6271_/Q _4539_/S vssd1 vssd1 vccd1 vccd1 _4528_/X sky130_fd_sc_hd__mux2_1
Xhold231 _6218_/Q vssd1 vssd1 vccd1 vccd1 hold231/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold253 _4332_/X vssd1 vssd1 vccd1 vccd1 _6094_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold264 _6429_/Q vssd1 vssd1 vccd1 vccd1 hold264/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold275 _4485_/X vssd1 vssd1 vccd1 vccd1 _6185_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4459_ _4392_/X hold111/X _4464_/S vssd1 vssd1 vccd1 vccd1 _4459_/X sky130_fd_sc_hd__mux2_1
Xhold286 _6199_/Q vssd1 vssd1 vccd1 vccd1 hold286/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold297 _6095_/Q vssd1 vssd1 vccd1 vccd1 hold297/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6129_ _6344_/CLK hold76/X vssd1 vssd1 vccd1 vccd1 hold75/A sky130_fd_sc_hd__dfxtp_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3608__A1 _3577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5069__C_N _4633_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3631__A _3632_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3350__B _5578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4024__A1 _6292_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3830_ _6179_/Q _3715_/X _3794_/X _6210_/Q _3829_/X vssd1 vssd1 vccd1 vccd1 _3831_/C
+ sky130_fd_sc_hd__a221o_1
X_3761_ _3761_/A vssd1 vssd1 vccd1 vccd1 _3761_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_27_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4575__A2 _4604_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5500_ _5554_/A _5501_/B vssd1 vssd1 vccd1 vccd1 _5502_/A sky130_fd_sc_hd__and2_1
X_3692_ _5247_/A _6304_/Q _5196_/S _3691_/Y vssd1 vssd1 vccd1 vccd1 _4633_/C sky130_fd_sc_hd__o31a_2
XFILLER_0_54_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5431_ _5427_/Y _5429_/X _5430_/X _5740_/A vssd1 vssd1 vccd1 vccd1 _5431_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_2_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5362_ _3410_/Y _3511_/D _5361_/Y _4214_/A vssd1 vssd1 vccd1 vccd1 _5362_/X sky130_fd_sc_hd__a22o_1
X_4313_ _6064_/S _4313_/B _4313_/C _4313_/D vssd1 vssd1 vccd1 vccd1 _4313_/Y sky130_fd_sc_hd__nand4_1
X_5293_ _5293_/A _5293_/B _5293_/C vssd1 vssd1 vccd1 vccd1 _5294_/D sky130_fd_sc_hd__or3_1
X_4244_ _5725_/B _5725_/A vssd1 vssd1 vccd1 vccd1 _4245_/S sky130_fd_sc_hd__nand2b_1
X_4175_ _6248_/Q _4174_/C _5217_/A vssd1 vssd1 vccd1 vccd1 _4176_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__4637__A _4637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3126_ _3183_/B _3116_/A _3285_/B _3116_/C vssd1 vssd1 vccd1 vccd1 _3126_/X sky130_fd_sc_hd__o211a_1
X_3057_ _6245_/Q vssd1 vssd1 vccd1 vccd1 _3970_/A sky130_fd_sc_hd__inv_2
XFILLER_0_89_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4263__A1 _3254_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6004__A2 _4807_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6063__S _6063_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3959_ _3061_/Y _3958_/X _4142_/S vssd1 vssd1 vccd1 vccd1 _6040_/A sky130_fd_sc_hd__mux2_8
XFILLER_0_18_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5763__B2 _5933_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5515__A1 _6057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5629_ _6269_/Q _5589_/X _5594_/Y _5628_/X vssd1 vssd1 vccd1 vccd1 _5629_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5407__S _5553_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3451__A _5935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold643_A _6422_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6046__A2_N _6054_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5097__B _5097_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6333__RESET_B fanout171/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6002__A _6036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5560__B _5560_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3296__A2 _5258_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5980_ _6424_/Q _5982_/S _5979_/Y hold306/X vssd1 vssd1 vccd1 vccd1 _5980_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5442__A0 _3952_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4931_ _5773_/A _4930_/X _4920_/Y vssd1 vssd1 vccd1 vccd1 _4931_/X sky130_fd_sc_hd__a21bo_1
XANTENNA__5993__A1 _6057_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4904__B _6324_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4862_ _4861_/X _4860_/X _5053_/S vssd1 vssd1 vccd1 vccd1 _4863_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_74_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3813_ _6165_/Q _3784_/X _3786_/X hold87/A vssd1 vssd1 vccd1 vccd1 _3813_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_74_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4793_ _4827_/C _4867_/B _4793_/C vssd1 vssd1 vccd1 vccd1 _4793_/X sky130_fd_sc_hd__and3b_1
X_3744_ _5087_/A _6242_/Q _6336_/Q _3740_/Y _3743_/X vssd1 vssd1 vccd1 vccd1 _5111_/A
+ sky130_fd_sc_hd__o41a_2
XFILLER_0_12_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4920__A _5054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3675_ _5322_/D _3661_/X _3662_/X _3655_/Y vssd1 vssd1 vccd1 vccd1 _3675_/X sky130_fd_sc_hd__o31a_1
XFILLER_0_15_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5414_ _4284_/A _6322_/Q _5442_/S vssd1 vssd1 vccd1 vccd1 _5414_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_88_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6394_ _6401_/CLK _6394_/D fanout179/X vssd1 vssd1 vccd1 vccd1 _6394_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5345_ _5339_/D _5344_/X _5979_/A vssd1 vssd1 vccd1 vccd1 _5345_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_56_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5276_ _3100_/B _4346_/B _4347_/C _3581_/A _5273_/X vssd1 vssd1 vccd1 vccd1 _5276_/X
+ sky130_fd_sc_hd__a221o_1
X_4227_ _5096_/B _4219_/X _4226_/X vssd1 vssd1 vccd1 vccd1 _5725_/A sky130_fd_sc_hd__o21ai_4
X_4158_ _4158_/A _4158_/B vssd1 vssd1 vccd1 vccd1 _4158_/X sky130_fd_sc_hd__and2_1
XFILLER_0_69_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5897__S _5931_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4236__A1 _4222_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3109_ _4255_/B _3109_/B vssd1 vssd1 vccd1 vccd1 _3459_/B sky130_fd_sc_hd__nand2_1
X_4089_ _6113_/Q _3779_/X _3781_/X _6104_/Q vssd1 vssd1 vccd1 vccd1 _4089_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5984__A1 _5518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5984__B2 _3473_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5736__A1 _5313_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4830__A _5058_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4227__A1 _5096_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput13 io_in[4] vssd1 vssd1 vccd1 vccd1 _3473_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_0_71_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3460_ _5560_/B _3443_/A _3449_/X _3459_/Y vssd1 vssd1 vccd1 vccd1 _3465_/B sky130_fd_sc_hd__a211oi_2
X_3391_ _3391_/A vssd1 vssd1 vccd1 vccd1 _3391_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_20_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5130_ _5130_/A _5130_/B vssd1 vssd1 vccd1 vccd1 _5134_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_58_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5061_ _5061_/A1 _5058_/X _5060_/X _4867_/B vssd1 vssd1 vccd1 vccd1 _5061_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3269__A2 _4222_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4012_ _3876_/X _3919_/A _4009_/X _4011_/X vssd1 vssd1 vccd1 vccd1 _4022_/A sky130_fd_sc_hd__o31ai_4
XANTENNA__5415__B1 _5371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5963_ _4399_/X hold301/X _5967_/S vssd1 vssd1 vccd1 vccd1 _6410_/D sky130_fd_sc_hd__mux2_1
XANTENNA__6255__RESET_B fanout179/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3977__B1 _6245_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4914_ _6326_/Q _4913_/X _5852_/S vssd1 vssd1 vccd1 vccd1 _4914_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_90_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5894_ _6331_/Q _5928_/A2 _5928_/B1 _5893_/X vssd1 vssd1 vccd1 vccd1 _5894_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_47_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3965__S _4427_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4845_ _6323_/Q _4846_/B vssd1 vssd1 vccd1 vccd1 _4847_/C sky130_fd_sc_hd__or2_1
XANTENNA__4650__A _6040_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5194__A2 _5075_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4776_ _5061_/A1 _4762_/X _4867_/B _4775_/X vssd1 vssd1 vccd1 vccd1 _4776_/X sky130_fd_sc_hd__a22o_1
X_3727_ _6304_/Q _5196_/S vssd1 vssd1 vccd1 vccd1 _3727_/X sky130_fd_sc_hd__and2_1
XFILLER_0_15_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3744__A3 _6336_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3658_ _4270_/B _3658_/B vssd1 vssd1 vccd1 vccd1 _3658_/Y sky130_fd_sc_hd__nor2_1
X_6446_ _6447_/CLK _6446_/D fanout171/X vssd1 vssd1 vccd1 vccd1 _6446_/Q sky130_fd_sc_hd__dfstp_1
X_3589_ _3334_/C _5733_/A _5480_/C _5481_/B _3588_/Y vssd1 vssd1 vccd1 vccd1 _4772_/A
+ sky130_fd_sc_hd__a2111o_1
XANTENNA__4154__B1 _3794_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6377_ _6386_/CLK _6377_/D fanout168/X vssd1 vssd1 vccd1 vccd1 _6377_/Q sky130_fd_sc_hd__dfrtp_4
X_5328_ _6390_/Q _5328_/B _5328_/C vssd1 vssd1 vccd1 vccd1 _5328_/X sky130_fd_sc_hd__and3_1
XANTENNA__4809__B _4809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5259_ _3116_/C _3148_/X _3152_/Y vssd1 vssd1 vccd1 vccd1 _5294_/C sky130_fd_sc_hd__a21oi_1
XFILLER_0_97_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5957__A1 _5715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold439_A _6339_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold606_A _6323_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5590__C1 _5676_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6487__A _6487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3499__A2 _5258_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_12_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_69_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output23_A _4732_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4630_ hold597/X _4615_/X _4617_/Y _4629_/X vssd1 vssd1 vccd1 vccd1 _4630_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_71_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6300_ _6403_/CLK _6300_/D fanout179/X vssd1 vssd1 vccd1 vccd1 _6300_/Q sky130_fd_sc_hd__dfrtp_1
X_4561_ _3183_/B _5313_/A _3686_/A _4555_/X _4560_/X vssd1 vssd1 vccd1 vccd1 _4604_/S
+ sky130_fd_sc_hd__a221o_4
XFILLER_0_71_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold627 _5307_/X vssd1 vssd1 vccd1 vccd1 _6303_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold616 _6304_/Q vssd1 vssd1 vccd1 vccd1 hold616/X sky130_fd_sc_hd__dlygate4sd3_1
X_3512_ _4639_/B _5359_/A vssd1 vssd1 vccd1 vccd1 _3512_/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_69_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold605 _6447_/Q vssd1 vssd1 vccd1 vccd1 _6054_/A sky130_fd_sc_hd__dlygate4sd3_1
X_4492_ _4510_/A _5959_/A vssd1 vssd1 vccd1 vccd1 _4500_/S sky130_fd_sc_hd__or2_4
XFILLER_0_40_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold638 _6396_/Q vssd1 vssd1 vccd1 vccd1 _5936_/B sky130_fd_sc_hd__buf_1
X_3443_ _3443_/A _5931_/S vssd1 vssd1 vccd1 vccd1 _3622_/A sky130_fd_sc_hd__or2_1
X_6231_ _6343_/CLK _6231_/D fanout170/X vssd1 vssd1 vccd1 vccd1 _6231_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_0_0_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold649 _6267_/Q vssd1 vssd1 vccd1 vccd1 _3072_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6162_ _6414_/CLK _6162_/D vssd1 vssd1 vccd1 vccd1 _6162_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_51_wb_clk_i_A clkbuf_leaf_6_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__4687__A1 _5240_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4629__B _4631_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5113_ _5113_/A _5113_/B vssd1 vssd1 vccd1 vccd1 _5114_/B sky130_fd_sc_hd__xnor2_1
X_3374_ _3374_/A _5328_/B vssd1 vssd1 vccd1 vccd1 _5481_/B sky130_fd_sc_hd__and2_1
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6093_ _6217_/CLK _6093_/D vssd1 vssd1 vccd1 vccd1 _6093_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5100__A2 _5192_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3252__C _4679_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5044_ _6385_/Q _4754_/X _5036_/X _5043_/X vssd1 vssd1 vccd1 vccd1 _5044_/X sky130_fd_sc_hd__a211o_1
XANTENNA__4645__A _6036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5240__S _5240_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout177_A fanout178/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5946_ _3621_/A _3625_/B hold566/X _3623_/A _3043_/A vssd1 vssd1 vccd1 vccd1 _5946_/X
+ sky130_fd_sc_hd__a32o_1
X_5877_ _6381_/Q _5926_/A _5868_/X vssd1 vssd1 vccd1 vccd1 _5878_/B sky130_fd_sc_hd__a21o_1
X_4828_ _6322_/Q _4828_/B vssd1 vssd1 vccd1 vccd1 _4828_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_90_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5167__A2 _5158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4759_ _5365_/C _4757_/Y _4758_/X _6416_/Q vssd1 vssd1 vccd1 vccd1 _4759_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_31_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6429_ _6430_/CLK _6429_/D fanout172/X vssd1 vssd1 vccd1 vccd1 _6429_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_12_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6209_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_101_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3443__B _5931_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5890__A3 _6381_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4850__B2 _4843_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4366__B1 _4382_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4669__A1 _6342_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3341__A1 _3654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6010__A _6044_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3892__A2 _6243_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3090_ _3290_/B _4522_/B vssd1 vssd1 vccd1 vccd1 _3206_/A sky130_fd_sc_hd__nor2_1
Xhold2 hold2/A vssd1 vssd1 vccd1 vccd1 hold2/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5094__A1 _5243_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5060__S _5060_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6043__B1 _6063_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3992_ _3992_/A _4158_/B vssd1 vssd1 vccd1 vccd1 _3992_/X sky130_fd_sc_hd__and2_1
Xci2406_z80_188 vssd1 vssd1 vccd1 vccd1 ci2406_z80_188/HI io_oeb[7] sky130_fd_sc_hd__conb_1
X_5800_ _6323_/Q _5852_/S _5799_/X vssd1 vssd1 vccd1 vccd1 _5800_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_71_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5731_ _5740_/A _5729_/X _3477_/X vssd1 vssd1 vccd1 vccd1 _5731_/X sky130_fd_sc_hd__a21o_2
Xci2406_z80_199 vssd1 vssd1 vccd1 vccd1 ci2406_z80_199/HI io_oeb[18] sky130_fd_sc_hd__conb_1
XFILLER_0_84_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5662_ _6197_/Q _4382_/B _4200_/S _6073_/Q _5675_/C1 vssd1 vssd1 vccd1 vccd1 _5664_/A
+ sky130_fd_sc_hd__o221a_1
X_4613_ input9/X _4631_/B vssd1 vssd1 vccd1 vccd1 _4613_/X sky130_fd_sc_hd__and2_1
XANTENNA__3528__B _4637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5593_ _6207_/Q _6313_/Q _3718_/Y _6128_/Q _3721_/Y vssd1 vssd1 vccd1 vccd1 _5595_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_44_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4544_ _5339_/C vssd1 vssd1 vccd1 vccd1 _4568_/C sky130_fd_sc_hd__inv_2
Xhold402 _5012_/X vssd1 vssd1 vccd1 vccd1 _6287_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold424 _3457_/X vssd1 vssd1 vccd1 vccd1 _3471_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold413 hold681/X vssd1 vssd1 vccd1 vccd1 _5989_/A sky130_fd_sc_hd__clkbuf_2
Xhold435 _6435_/Q vssd1 vssd1 vccd1 vccd1 hold435/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold468 _6240_/Q vssd1 vssd1 vccd1 vccd1 hold468/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold457 _6341_/Q vssd1 vssd1 vccd1 vccd1 _4056_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold446 _4531_/X vssd1 vssd1 vccd1 vccd1 _6232_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4475_ _4367_/X hold214/X _4482_/S vssd1 vssd1 vccd1 vccd1 _4475_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_13_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6214_ _6410_/CLK _6214_/D vssd1 vssd1 vccd1 vccd1 _6214_/Q sky130_fd_sc_hd__dfxtp_1
X_3426_ _3426_/A _3426_/B _3426_/C vssd1 vssd1 vccd1 vccd1 _3426_/X sky130_fd_sc_hd__or3_1
Xhold479 _4537_/X vssd1 vssd1 vccd1 vccd1 _6238_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3263__B _3654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3357_ _3686_/A _5359_/A _3357_/C _3357_/D vssd1 vssd1 vccd1 vccd1 _3357_/X sky130_fd_sc_hd__or4_1
X_6145_ _6344_/CLK _6145_/D vssd1 vssd1 vccd1 vccd1 _6145_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6076_ _6428_/CLK hold2/X vssd1 vssd1 vccd1 vccd1 hold1/A sky130_fd_sc_hd__dfxtp_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3288_ _3658_/B _4550_/B _3367_/B vssd1 vssd1 vccd1 vccd1 _3339_/A sky130_fd_sc_hd__and3_1
X_5027_ _5929_/A1 _5026_/X _5016_/Y vssd1 vssd1 vccd1 vccd1 _5027_/X sky130_fd_sc_hd__a21bo_1
XANTENNA__4832__B2 _4830_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5388__A2 _5377_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6034__B1 _6057_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5929_ _5929_/A1 _5928_/X _5054_/Y vssd1 vssd1 vccd1 vccd1 _5929_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_63_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4994__S1 _4326_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4984__S _5060_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3626__A2 _4287_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4285__A _4685_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4260_ _4260_/A _4260_/B vssd1 vssd1 vccd1 vccd1 _4260_/X sky130_fd_sc_hd__or2_1
XFILLER_0_10_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3211_ _3496_/A _5715_/C vssd1 vssd1 vccd1 vccd1 _3211_/X sky130_fd_sc_hd__or2_1
X_4191_ _6423_/Q _4190_/X _4191_/S vssd1 vssd1 vccd1 vccd1 _4191_/X sky130_fd_sc_hd__mux2_1
X_3142_ _3091_/X _3379_/B _3426_/A vssd1 vssd1 vccd1 vccd1 _3600_/A sky130_fd_sc_hd__o21bai_2
X_3073_ _3073_/A vssd1 vssd1 vccd1 vccd1 _3073_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4814__A1 _4867_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3530__C _4228_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4290__A2 _4287_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6016__B1 _6057_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3975_ _3740_/Y _3973_/X _3974_/X vssd1 vssd1 vccd1 vccd1 _3975_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_92_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5790__A2 _6420_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5714_ hold25/X _4156_/B _6064_/S vssd1 vssd1 vccd1 vccd1 hold26/A sky130_fd_sc_hd__mux2_1
XANTENNA__3258__B _6389_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5645_ _5695_/A1 _3992_/A _5571_/Y _5644_/X vssd1 vssd1 vccd1 vccd1 _5645_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5576_ _3572_/A _4551_/Y _5575_/X _5317_/A vssd1 vssd1 vccd1 vccd1 _5576_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_5_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold210 _6181_/Q vssd1 vssd1 vccd1 vccd1 hold210/X sky130_fd_sc_hd__dlygate4sd3_1
X_4527_ hold488/X _6270_/Q _4539_/S vssd1 vssd1 vccd1 vccd1 _4527_/X sky130_fd_sc_hd__mux2_1
Xhold221 _4432_/X vssd1 vssd1 vccd1 vccd1 _6138_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold232 _4514_/X vssd1 vssd1 vccd1 vccd1 _6218_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold243 _6198_/Q vssd1 vssd1 vccd1 vccd1 hold243/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold265 _5987_/X vssd1 vssd1 vccd1 vccd1 _6430_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold254 _6145_/Q vssd1 vssd1 vccd1 vccd1 hold254/X sky130_fd_sc_hd__dlygate4sd3_1
X_4458_ _4380_/X hold167/X _4464_/S vssd1 vssd1 vccd1 vccd1 _4458_/X sky130_fd_sc_hd__mux2_1
Xhold287 _4500_/X vssd1 vssd1 vccd1 vccd1 _6199_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold276 _6183_/Q vssd1 vssd1 vccd1 vccd1 hold276/X sky130_fd_sc_hd__dlygate4sd3_1
X_3409_ _4210_/A _3409_/B vssd1 vssd1 vccd1 vccd1 _4637_/B sky130_fd_sc_hd__nand2_4
Xhold298 _6068_/Q vssd1 vssd1 vccd1 vccd1 hold298/X sky130_fd_sc_hd__dlygate4sd3_1
X_6128_ _6209_/CLK _6128_/D vssd1 vssd1 vccd1 vccd1 _6128_/Q sky130_fd_sc_hd__dfxtp_1
X_4389_ _4389_/A _5249_/C vssd1 vssd1 vccd1 vccd1 _4389_/X sky130_fd_sc_hd__xor2_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3608__A2 _5956_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6059_ _6022_/A _6063_/S _6056_/Y _6058_/X vssd1 vssd1 vccd1 vccd1 _6059_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_95_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4979__S _6315_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3544__A1 _5097_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5297__A1 _4224_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4272__A2 _3654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3760_ _3757_/B _3760_/B _6304_/Q vssd1 vssd1 vccd1 vccd1 _3761_/A sky130_fd_sc_hd__and3b_4
XANTENNA__5221__B2 _6297_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3359__A _5313_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3691_ _5247_/A _3691_/B vssd1 vssd1 vccd1 vccd1 _3691_/Y sky130_fd_sc_hd__nand2_1
X_5430_ hold606/X input2/X _5469_/S vssd1 vssd1 vccd1 vccd1 _5430_/X sky130_fd_sc_hd__mux2_1
X_5361_ _3611_/A _3367_/B _5360_/X vssd1 vssd1 vccd1 vccd1 _5361_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_2_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3525__C _5077_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5292_ _5292_/A _5292_/B _5292_/C _5292_/D vssd1 vssd1 vccd1 vccd1 _5293_/C sky130_fd_sc_hd__or4_1
XFILLER_0_77_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4312_ _4313_/B _4311_/Y _5447_/S vssd1 vssd1 vccd1 vccd1 _4312_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_2_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5288__A1 _6256_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4243_ _4279_/A _4243_/B vssd1 vssd1 vccd1 vccd1 _5725_/B sky130_fd_sc_hd__nand2_1
X_4174_ _5217_/A _6248_/Q _4174_/C vssd1 vssd1 vccd1 vccd1 _4176_/A sky130_fd_sc_hd__or3_1
XANTENNA__4637__B _4637_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3125_ _3116_/A _4522_/D _3122_/X _4679_/C vssd1 vssd1 vccd1 vccd1 _3125_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_96_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3056_ _6242_/Q vssd1 vssd1 vccd1 vccd1 _4183_/B sky130_fd_sc_hd__inv_2
XFILLER_0_89_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4653__A _6044_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4015__A2 _3789_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3958_ _5393_/B _3957_/X _6305_/Q vssd1 vssd1 vccd1 vccd1 _3958_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_9_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3889_ _3889_/A _3889_/B vssd1 vssd1 vccd1 vccd1 _3889_/X sky130_fd_sc_hd__xor2_1
XANTENNA__5484__A _5553_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5628_ _5627_/X _4388_/X _5691_/S vssd1 vssd1 vccd1 vccd1 _5628_/X sky130_fd_sc_hd__mux2_1
X_5559_ hold526/X _5558_/X _6060_/S vssd1 vssd1 vccd1 vccd1 _5559_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3716__B _3850_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5279__A1 _3573_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3732__A _6242_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3829__A2 _3789_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4828__A _6322_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout72_A _5673_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3451__B _6392_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4254__A2 _5315_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4962__A0 _4958_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4502__S _4509_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3517__A1 _4070_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6373__RESET_B fanout169/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6302__RESET_B fanout179/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6439__SET_B fanout181/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3642__A _5077_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4738__A _5728_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5442__A1 _6324_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4930_ _6327_/Q _5825_/S _5928_/B1 _4929_/X vssd1 vssd1 vccd1 vccd1 _4930_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_74_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4861_ _6165_/Q hold87/A _6412_/Q _6181_/Q _5051_/S0 _5052_/S1 vssd1 vssd1 vccd1
+ vccd1 _4861_/X sky130_fd_sc_hd__mux4_1
XANTENNA__4904__C _6325_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3812_ _4394_/A _4599_/A vssd1 vssd1 vccd1 vccd1 _4416_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__3756__A1 _6336_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4792_ _5060_/S _4905_/C vssd1 vssd1 vccd1 vccd1 _4827_/C sky130_fd_sc_hd__and2_1
X_3743_ _3737_/X _3738_/Y _3740_/Y _3742_/X vssd1 vssd1 vccd1 vccd1 _3743_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_70_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5508__S _6060_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4920__B _4920_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3674_ _3674_/A _3674_/B vssd1 vssd1 vccd1 vccd1 _5991_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_70_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6393_ _6430_/CLK _6393_/D fanout172/X vssd1 vssd1 vccd1 vccd1 _6393_/Q sky130_fd_sc_hd__dfrtp_1
X_5413_ _5441_/A _5413_/B vssd1 vssd1 vccd1 vccd1 _5413_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_30_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4181__A1 _6292_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5344_ _5584_/A1 _5341_/X _5343_/X _3530_/D _5313_/X vssd1 vssd1 vccd1 vccd1 _5344_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_23_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5275_ _5096_/B _5268_/X _5274_/X _3530_/D _5263_/X vssd1 vssd1 vccd1 vccd1 _5275_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5243__S _5243_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4226_ _4228_/A _4225_/X _4221_/X _4260_/B vssd1 vssd1 vccd1 vccd1 _4226_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_49_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3271__B _3502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4157_ _4157_/A _4157_/B vssd1 vssd1 vccd1 vccd1 _4157_/Y sky130_fd_sc_hd__xnor2_1
X_3108_ _4223_/B _3344_/A vssd1 vssd1 vccd1 vccd1 _3451_/C sky130_fd_sc_hd__nor2_2
X_4088_ _3724_/A _6052_/A _4425_/A2 vssd1 vssd1 vccd1 vccd1 _4088_/Y sky130_fd_sc_hd__o21ai_1
X_3039_ _5265_/A vssd1 vssd1 vccd1 vccd1 _3039_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_37_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6384_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5736__A2 _3451_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4830__B _4830_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3727__A _6304_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput14 rst_n vssd1 vssd1 vccd1 vccd1 input14/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_52_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_41_wb_clk_i_A clkbuf_leaf_6_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_3390_ _3770_/A _5728_/B _3611_/A vssd1 vssd1 vccd1 vccd1 _3391_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_20_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3372__A _4520_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5060_ _6423_/Q _5059_/X _5060_/S vssd1 vssd1 vccd1 vccd1 _5060_/X sky130_fd_sc_hd__mux2_1
X_4011_ _3934_/B _4009_/X _4010_/Y vssd1 vssd1 vccd1 vccd1 _4011_/X sky130_fd_sc_hd__o21a_1
XANTENNA__4218__A2 _5733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5415__A1 _5441_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5962_ _4392_/X hold130/X _5967_/S vssd1 vssd1 vccd1 vccd1 _5962_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3977__A1 _6243_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4913_ _5773_/A _4912_/X _4900_/Y vssd1 vssd1 vccd1 vccd1 _4913_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_90_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5893_ _6364_/Q _6383_/Q _5927_/S vssd1 vssd1 vccd1 vccd1 _5893_/X sky130_fd_sc_hd__mux2_1
X_4844_ _5054_/A _4843_/X _5728_/D vssd1 vssd1 vccd1 vccd1 _4844_/X sky130_fd_sc_hd__a21o_1
X_4775_ _6319_/Q _5060_/S vssd1 vssd1 vccd1 vccd1 _4775_/X sky130_fd_sc_hd__xor2_1
XANTENNA__4926__A0 _6416_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6030__A2_N _6054_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6224__RESET_B fanout179/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3726_ _4158_/B vssd1 vssd1 vccd1 vccd1 _4142_/S sky130_fd_sc_hd__inv_4
XFILLER_0_43_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3657_ _3657_/A _3657_/B vssd1 vssd1 vccd1 vccd1 _4274_/A sky130_fd_sc_hd__and2_1
XFILLER_0_15_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6445_ _6445_/CLK _6445_/D fanout171/X vssd1 vssd1 vccd1 vccd1 _6445_/Q sky130_fd_sc_hd__dfstp_1
X_3588_ _4679_/C _4679_/D vssd1 vssd1 vccd1 vccd1 _3588_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_2_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6376_ _6376_/CLK _6376_/D fanout166/X vssd1 vssd1 vccd1 vccd1 _6376_/Q sky130_fd_sc_hd__dfrtp_4
X_5327_ _5327_/A _5482_/A _5327_/C _5327_/D vssd1 vssd1 vccd1 vccd1 _5330_/S sky130_fd_sc_hd__or4_1
X_5258_ _5578_/A _5258_/B vssd1 vssd1 vccd1 vccd1 _5258_/Y sky130_fd_sc_hd__nor2_1
X_4209_ _4747_/D _4349_/C vssd1 vssd1 vccd1 vccd1 _4209_/Y sky130_fd_sc_hd__nor2_1
X_5189_ _5186_/X _5188_/X _5102_/B _5185_/Y vssd1 vssd1 vccd1 vccd1 _5189_/X sky130_fd_sc_hd__a2bb2o_1
XANTENNA__5701__S _6060_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3417__B1 _4541_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3432__A3 _4734_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4090__B1 _3786_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4393__A1 _4392_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5590__B1 _5676_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5645__A1 _5695_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout180 fanout181/X vssd1 vssd1 vccd1 vccd1 fanout180/X sky130_fd_sc_hd__buf_4
XFILLER_0_88_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_8_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__4620__A2 _4615_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4560_ _4260_/A _4559_/X _5096_/B vssd1 vssd1 vccd1 vccd1 _4560_/X sky130_fd_sc_hd__o21a_1
XANTENNA__5058__S _5058_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3511_ _3511_/A _5292_/C _3511_/C _3511_/D vssd1 vssd1 vccd1 vccd1 _3511_/X sky130_fd_sc_hd__or4_1
Xhold606 _6323_/Q vssd1 vssd1 vccd1 vccd1 hold606/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold617 _6298_/Q vssd1 vssd1 vccd1 vccd1 hold617/X sky130_fd_sc_hd__dlygate4sd3_1
X_4491_ hold71/X _4427_/X _4491_/S vssd1 vssd1 vccd1 vccd1 hold72/A sky130_fd_sc_hd__mux2_1
XFILLER_0_100_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4136__A1 _6248_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold639 _5943_/X vssd1 vssd1 vccd1 vccd1 hold639/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold628 _6392_/Q vssd1 vssd1 vccd1 vccd1 _4323_/A sky130_fd_sc_hd__clkbuf_2
X_3442_ _5931_/S vssd1 vssd1 vccd1 vccd1 _5979_/A sky130_fd_sc_hd__inv_2
X_6230_ _6271_/CLK _6230_/D fanout170/X vssd1 vssd1 vccd1 vccd1 _6230_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_0_100_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3373_ _3373_/A _3373_/B vssd1 vssd1 vccd1 vccd1 _5324_/B sky130_fd_sc_hd__or2_1
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6161_ _6407_/CLK _6161_/D vssd1 vssd1 vccd1 vccd1 _6161_/Q sky130_fd_sc_hd__dfxtp_1
X_5112_ _5112_/A _5205_/B vssd1 vssd1 vccd1 vccd1 _5113_/B sky130_fd_sc_hd__xnor2_1
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6092_ _6217_/CLK _6092_/D vssd1 vssd1 vccd1 vccd1 _6092_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5043_ _5061_/A1 _5038_/X _5042_/X _4867_/B vssd1 vssd1 vccd1 vccd1 _5043_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_79_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6061__A1 _6057_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5945_ _5952_/A _3457_/A hold565/X _5937_/Y vssd1 vssd1 vccd1 vccd1 _5945_/X sky130_fd_sc_hd__a22o_1
XANTENNA__6405__RESET_B fanout178/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5876_ _5876_/A _5926_/A vssd1 vssd1 vccd1 vccd1 _5889_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_7_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4827_ _6321_/Q _6322_/Q _4827_/C vssd1 vssd1 vccd1 vccd1 _4846_/B sky130_fd_sc_hd__and3_1
XFILLER_0_90_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4375__A1 _5690_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4758_ _4757_/B _4758_/B _4758_/C vssd1 vssd1 vccd1 vccd1 _4758_/X sky130_fd_sc_hd__and3b_4
XFILLER_0_7_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3709_ _3700_/C _3702_/X _3707_/X _3708_/Y vssd1 vssd1 vccd1 vccd1 _3850_/B sky130_fd_sc_hd__o31ai_4
X_4689_ _6032_/A _4731_/S _4688_/X vssd1 vssd1 vccd1 vccd1 _4689_/Y sky130_fd_sc_hd__o21ai_1
X_6428_ _6428_/CLK _6428_/D fanout172/X vssd1 vssd1 vccd1 vccd1 _6428_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6359_ _6444_/CLK hold26/X vssd1 vssd1 vccd1 vccd1 hold25/A sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_52_wb_clk_i clkbuf_leaf_6_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6412_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_98_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold549_A _6243_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5866__A1 _6379_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5618__A1 _6292_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3892__A3 _6337_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold3 hold3/A vssd1 vssd1 vccd1 vccd1 hold3/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6043__A1 _6057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3991_ _6419_/Q _3990_/X _4085_/S vssd1 vssd1 vccd1 vccd1 _3991_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_71_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5730_ _5740_/A _5729_/X _3477_/X vssd1 vssd1 vccd1 vccd1 _5933_/S sky130_fd_sc_hd__a21oi_4
Xci2406_z80_189 vssd1 vssd1 vccd1 vccd1 ci2406_z80_189/HI io_oeb[8] sky130_fd_sc_hd__conb_1
XFILLER_0_29_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3801__B1 _3786_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5661_ _5661_/A _5661_/B vssd1 vssd1 vccd1 vccd1 _5661_/X sky130_fd_sc_hd__or2_1
XFILLER_0_72_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4612_ _5740_/A _5372_/B vssd1 vssd1 vccd1 vccd1 _4631_/B sky130_fd_sc_hd__nand2_2
X_5592_ _6176_/Q _4382_/B _3718_/Y _6407_/Q _5673_/C1 vssd1 vssd1 vccd1 vccd1 _5592_/X
+ sky130_fd_sc_hd__a221o_1
X_4543_ _5096_/B _4540_/X _4542_/X _3530_/D vssd1 vssd1 vccd1 vccd1 _5339_/C sky130_fd_sc_hd__a22oi_4
XFILLER_0_4_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold425 _6342_/Q vssd1 vssd1 vccd1 vccd1 _3063_/A sky130_fd_sc_hd__buf_1
Xhold403 _6288_/Q vssd1 vssd1 vccd1 vccd1 hold403/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold414 _6439_/Q vssd1 vssd1 vccd1 vccd1 hold414/X sky130_fd_sc_hd__buf_1
Xhold436 _6007_/X vssd1 vssd1 vccd1 vccd1 _6435_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold469 _4539_/X vssd1 vssd1 vccd1 vccd1 _6240_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold458 _5671_/X vssd1 vssd1 vccd1 vccd1 _6341_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold447 _6290_/Q vssd1 vssd1 vccd1 vccd1 hold447/X sky130_fd_sc_hd__dlygate4sd3_1
X_4474_ _4474_/A _5959_/B vssd1 vssd1 vccd1 vccd1 _4482_/S sky130_fd_sc_hd__or2_4
X_6213_ _6413_/CLK _6213_/D vssd1 vssd1 vccd1 vccd1 _6213_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3425_ _3391_/A _3424_/X _5270_/A vssd1 vssd1 vccd1 vccd1 _3426_/C sky130_fd_sc_hd__o21a_1
X_3356_ _3224_/X _3501_/B _3611_/A vssd1 vssd1 vccd1 vccd1 _3356_/Y sky130_fd_sc_hd__a21oi_1
X_6144_ _6344_/CLK hold92/X vssd1 vssd1 vccd1 vccd1 hold91/A sky130_fd_sc_hd__dfxtp_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5609__A1 _5695_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3287_ _4550_/B _3367_/B vssd1 vssd1 vccd1 vccd1 _3287_/Y sky130_fd_sc_hd__nand2_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6075_ _6355_/CLK _6075_/D vssd1 vssd1 vccd1 vccd1 _6075_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5026_ _6332_/Q _5928_/A2 _5928_/B1 _5025_/X vssd1 vssd1 vccd1 vccd1 _5026_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_95_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6034__B2 _4938_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5928_ _6334_/Q _5928_/A2 _5928_/B1 _5927_/X vssd1 vssd1 vccd1 vccd1 _5928_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4596__A1 _6421_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4596__B2 _6272_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3719__B _5597_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5859_ _6361_/Q _6380_/Q _5927_/S vssd1 vssd1 vccd1 vccd1 _5859_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_8_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4330__S _4336_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6398__RESET_B fanout178/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4285__B _5553_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6327__RESET_B fanout168/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6025__A1 _6057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4505__S _4509_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5784__A0 _6322_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3562__A2 _4734_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5839__A1 _6326_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4190_ _4040_/A _5109_/B _4182_/X _4189_/X vssd1 vssd1 vccd1 vccd1 _4190_/X sky130_fd_sc_hd__a211o_1
X_3210_ _4284_/A _5226_/A vssd1 vssd1 vccd1 vccd1 _5715_/C sky130_fd_sc_hd__or2_4
X_3141_ _3549_/A _3220_/A _3186_/B vssd1 vssd1 vccd1 vccd1 _3426_/A sky130_fd_sc_hd__nor3_4
XANTENNA__3380__A _4214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3072_ _3072_/A vssd1 vssd1 vccd1 vccd1 _3072_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4027__A0 _6245_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6016__B2 _4863_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4578__A1 _5695_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3974_ _5087_/B _3969_/X _3973_/A _3741_/X vssd1 vssd1 vccd1 vccd1 _3974_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_57_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5713_ hold29/X _4111_/B _6064_/S vssd1 vssd1 vccd1 vccd1 hold30/A sky130_fd_sc_hd__mux2_1
XFILLER_0_60_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5790__A3 _3580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5644_ _5644_/A _5644_/B vssd1 vssd1 vccd1 vccd1 _5644_/X sky130_fd_sc_hd__or2_1
XFILLER_0_32_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5575_ _3546_/Y _4550_/C _5574_/Y _4257_/Y _4224_/A vssd1 vssd1 vccd1 vccd1 _5575_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_79_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold200 _4330_/X vssd1 vssd1 vccd1 vccd1 _6092_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold211 _4480_/X vssd1 vssd1 vccd1 vccd1 _6181_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3274__B _4520_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4526_ hold451/X _6269_/Q _4539_/S vssd1 vssd1 vccd1 vccd1 _4526_/X sky130_fd_sc_hd__mux2_1
Xhold244 _6194_/Q vssd1 vssd1 vccd1 vccd1 hold244/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold233 _6152_/Q vssd1 vssd1 vccd1 vccd1 hold233/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold222 _6132_/Q vssd1 vssd1 vccd1 vccd1 hold222/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold255 _4440_/X vssd1 vssd1 vccd1 vccd1 _6145_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4457_ _4367_/X hold95/X _4464_/S vssd1 vssd1 vccd1 vccd1 hold96/A sky130_fd_sc_hd__mux2_1
Xhold266 _6164_/Q vssd1 vssd1 vccd1 vccd1 hold266/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold277 _4482_/X vssd1 vssd1 vccd1 vccd1 _6183_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3408_ _4210_/A _5574_/A _6390_/Q vssd1 vssd1 vccd1 vccd1 _4767_/B sky130_fd_sc_hd__and3_2
Xhold288 _6217_/Q vssd1 vssd1 vccd1 vccd1 hold288/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold299 _3882_/X vssd1 vssd1 vccd1 vccd1 _6068_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6127_ _6406_/CLK _6127_/D fanout180/X vssd1 vssd1 vccd1 vccd1 _6127_/Q sky130_fd_sc_hd__dfstp_1
X_4388_ _5690_/S _4385_/X _4386_/X _4387_/X vssd1 vssd1 vccd1 vccd1 _4388_/X sky130_fd_sc_hd__o31a_1
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3339_ _3339_/A _3339_/B vssd1 vssd1 vccd1 vccd1 _3349_/B sky130_fd_sc_hd__nor2_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6058_ _6054_/A _5557_/S _6063_/S _6057_/X vssd1 vssd1 vccd1 vccd1 _6058_/X sky130_fd_sc_hd__o211a_1
X_5009_ _5929_/A1 _5008_/X _4996_/Y vssd1 vssd1 vccd1 vccd1 _5009_/X sky130_fd_sc_hd__a21bo_1
XANTENNA__6007__A1 _5339_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3449__B _5956_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5156__S _5240_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4995__S _5053_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3690_ _5097_/A _3690_/B vssd1 vssd1 vccd1 vccd1 _3691_/B sky130_fd_sc_hd__or2_4
XANTENNA__3375__A _5733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_502 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5360_ _3600_/C _5360_/B _5360_/C vssd1 vssd1 vccd1 vccd1 _5360_/X sky130_fd_sc_hd__and3b_1
XFILLER_0_2_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3094__B _3183_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3525__D _4070_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5291_ _5291_/A _5291_/B _3367_/B vssd1 vssd1 vccd1 vccd1 _5292_/D sky130_fd_sc_hd__or3b_1
XFILLER_0_65_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4311_ _3075_/Y _4305_/S _4310_/X vssd1 vssd1 vccd1 vccd1 _4311_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_10_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4242_ _4568_/B vssd1 vssd1 vccd1 vccd1 _4243_/B sky130_fd_sc_hd__inv_2
XFILLER_0_10_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4173_ _4172_/C _4172_/B _4171_/X vssd1 vssd1 vccd1 vccd1 _4173_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_0_93_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3124_ _3525_/B _3243_/B vssd1 vssd1 vccd1 vccd1 _4679_/C sky130_fd_sc_hd__or2_2
X_3055_ _6244_/Q vssd1 vssd1 vccd1 vccd1 _3939_/A sky130_fd_sc_hd__inv_2
XANTENNA__5996__B1 _6057_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout152_A _3566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3957_ _4040_/A _5112_/A _3956_/X vssd1 vssd1 vccd1 vccd1 _3957_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_73_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3888_ _4183_/B _3732_/B _3738_/Y vssd1 vssd1 vccd1 vccd1 _3889_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__5484__B _5484_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5627_ _5626_/X _3964_/X _5690_/S vssd1 vssd1 vccd1 vccd1 _5627_/X sky130_fd_sc_hd__mux2_1
X_5558_ _6423_/Q _5557_/X _5558_/S vssd1 vssd1 vccd1 vccd1 _5558_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4723__A1 _6273_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4723__B2 _5371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4509_ hold151/X _4427_/X _4509_/S vssd1 vssd1 vccd1 vccd1 _4509_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5279__A2 _4685_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5489_ _5554_/A _5489_/B vssd1 vssd1 vccd1 vccd1 _5492_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__5704__S _6060_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4239__B1 _4221_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3451__C _3451_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3517__A2 _3952_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_31_wb_clk_i_A clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_20_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_7_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6351_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__3642__B _4255_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5675__C1 _5675_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5560__D _5560_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output46_A _3048_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4860_ _6189_/Q hold49/A _6133_/Q _6212_/Q _5051_/S0 _5052_/S1 vssd1 vssd1 vccd1
+ vccd1 _4860_/X sky130_fd_sc_hd__mux4_1
XANTENNA__4904__D _6326_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3811_ _4599_/A vssd1 vssd1 vccd1 vccd1 _3811_/Y sky130_fd_sc_hd__inv_2
X_4791_ _6319_/Q _6320_/Q vssd1 vssd1 vccd1 vccd1 _4905_/C sky130_fd_sc_hd__and2_1
X_3742_ _5087_/B _3731_/X _3738_/A _3741_/X vssd1 vssd1 vccd1 vccd1 _3742_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_12_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3673_ _5096_/B _3671_/X _3672_/X _3655_/Y vssd1 vssd1 vccd1 vccd1 _3674_/B sky130_fd_sc_hd__a22oi_4
XFILLER_0_42_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6392_ _6430_/CLK _6392_/D fanout172/X vssd1 vssd1 vccd1 vccd1 _6392_/Q sky130_fd_sc_hd__dfrtp_4
X_5412_ _5412_/A _5412_/B vssd1 vssd1 vccd1 vccd1 _5413_/B sky130_fd_sc_hd__xor2_1
X_5343_ _5343_/A _5343_/B _5343_/C _5343_/D vssd1 vssd1 vccd1 vccd1 _5343_/X sky130_fd_sc_hd__or4_1
XFILLER_0_88_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5274_ _4210_/A _4347_/C _5273_/X _3549_/A vssd1 vssd1 vccd1 vccd1 _5274_/X sky130_fd_sc_hd__a22o_1
X_4225_ _3594_/A _5341_/B _5341_/A vssd1 vssd1 vccd1 vccd1 _4225_/X sky130_fd_sc_hd__a21o_1
XANTENNA__6083__RESET_B fanout169/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4156_ _4156_/A _4156_/B vssd1 vssd1 vccd1 vccd1 _4157_/B sky130_fd_sc_hd__xnor2_1
X_3107_ _5258_/B _3292_/C vssd1 vssd1 vccd1 vccd1 _3344_/A sky130_fd_sc_hd__nand2_2
XANTENNA__5969__A0 input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4087_ _6052_/A vssd1 vssd1 vccd1 vccd1 _4087_/Y sky130_fd_sc_hd__inv_2
X_3038_ _4541_/A vssd1 vssd1 vccd1 vccd1 _4210_/A sky130_fd_sc_hd__clkinv_4
XFILLER_0_93_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3995__A2 _6044_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5197__A1 _6341_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4989_ _5929_/A1 _4988_/X _4976_/Y vssd1 vssd1 vccd1 vccd1 _4989_/X sky130_fd_sc_hd__a21bo_1
XANTENNA__6445__SET_B fanout171/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4558__B _5578_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5672__A2 _6313_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4632__B1 _4617_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5188__A1 _5371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4513__S _4518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3910__A2 _6036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5663__A2 _4382_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4010_ _3930_/B _4001_/B _4111_/A vssd1 vssd1 vccd1 vccd1 _4010_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_79_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4218__A3 _3770_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5961_ _4380_/X hold239/X _5967_/S vssd1 vssd1 vccd1 vccd1 _5961_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3977__A2 _6244_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4912_ _6326_/Q _5825_/S _5850_/B1 _4911_/X vssd1 vssd1 vccd1 vccd1 _4912_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_47_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5892_ _5892_/A _5892_/B vssd1 vssd1 vccd1 vccd1 _5892_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_74_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4843_ _4842_/X _4841_/X _5053_/S vssd1 vssd1 vccd1 vccd1 _4843_/X sky130_fd_sc_hd__mux2_4
X_4774_ _4774_/A _4774_/B vssd1 vssd1 vccd1 vccd1 _4809_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_7_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3725_ _5560_/A _3725_/B _3725_/C vssd1 vssd1 vccd1 vccd1 _4158_/B sky130_fd_sc_hd__nor3_4
XFILLER_0_70_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6444_ _6444_/CLK _6444_/D fanout171/X vssd1 vssd1 vccd1 vccd1 _6444_/Q sky130_fd_sc_hd__dfstp_1
X_3656_ _3656_/A _5322_/D vssd1 vssd1 vccd1 vccd1 _3656_/X sky130_fd_sc_hd__and2_1
XANTENNA_fanout115_A _5553_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6264__RESET_B fanout177/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3587_ _3278_/A _3566_/B _4745_/B _3586_/X vssd1 vssd1 vccd1 vccd1 _3587_/X sky130_fd_sc_hd__o31a_1
XFILLER_0_61_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4154__A2 _3715_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6375_ _6376_/CLK _6375_/D fanout169/X vssd1 vssd1 vccd1 vccd1 _6375_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__5351__A1 _5603_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4785__S0 _4326_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5326_ _5481_/A _5326_/B _5326_/C _5326_/D vssd1 vssd1 vccd1 vccd1 _5327_/D sky130_fd_sc_hd__or4_1
XFILLER_0_11_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5257_ _3549_/A _5256_/B _5256_/Y _3373_/A _5258_/B vssd1 vssd1 vccd1 vccd1 _5257_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA__3282__B _3573_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5103__A1 _6292_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5103__B2 _5740_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4208_ _4223_/B _4208_/B vssd1 vssd1 vccd1 vccd1 _4349_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_48_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5188_ _5371_/A _5187_/X _5102_/Y vssd1 vssd1 vccd1 vccd1 _5188_/X sky130_fd_sc_hd__a21bo_1
X_4139_ _3758_/Y _5120_/A _4136_/X _4138_/X vssd1 vssd1 vccd1 vccd1 _4139_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_97_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4614__B1 _5740_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4333__S _4336_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5342__A1 _3770_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3473__A _3473_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout181 input14/X vssd1 vssd1 vccd1 vccd1 fanout181/X sky130_fd_sc_hd__clkbuf_8
Xfanout170 fanout181/X vssd1 vssd1 vccd1 vccd1 fanout170/X sky130_fd_sc_hd__buf_4
XFILLER_0_44_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4508__S _4509_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4908__B2 _4900_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3510_ _6405_/Q _3510_/B _6400_/Q vssd1 vssd1 vccd1 vccd1 _3511_/D sky130_fd_sc_hd__and3b_1
XFILLER_0_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold607 _5433_/X vssd1 vssd1 vccd1 vccd1 _6323_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold618 _5244_/X vssd1 vssd1 vccd1 vccd1 _6298_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4490_ hold159/X _4420_/X _4491_/S vssd1 vssd1 vccd1 vccd1 _4490_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_100_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold629 _5951_/X vssd1 vssd1 vccd1 vccd1 _6392_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3441_ _3047_/Y _3439_/S _3436_/B _3435_/Y _3440_/Y vssd1 vssd1 vccd1 vccd1 _5977_/S
+ sky130_fd_sc_hd__o41a_4
XANTENNA__5333__A1 _4604_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3372_ _4520_/B _5291_/B _4541_/D vssd1 vssd1 vccd1 vccd1 _5326_/B sky130_fd_sc_hd__or3_1
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6160_ _6407_/CLK hold96/X vssd1 vssd1 vccd1 vccd1 hold95/A sky130_fd_sc_hd__dfxtp_1
X_5111_ _5111_/A _5111_/B vssd1 vssd1 vccd1 vccd1 _5113_/A sky130_fd_sc_hd__xor2_1
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4198__B _4198_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5636__A2 _4198_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6091_ _6221_/CLK _6091_/D vssd1 vssd1 vccd1 vccd1 _6091_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5042_ _6422_/Q _5041_/Y _5060_/S vssd1 vssd1 vccd1 vccd1 _5042_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4844__B1 _5728_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5944_ _3621_/A _3625_/B hold639/X _3623_/A _3457_/A vssd1 vssd1 vccd1 vccd1 _5944_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5875_ _5865_/A _5742_/A _5874_/X _5731_/X vssd1 vssd1 vccd1 vccd1 _5875_/X sky130_fd_sc_hd__o22a_1
X_4826_ _5054_/A _4830_/B _5728_/D vssd1 vssd1 vccd1 vccd1 _4826_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_7_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4757_ _4758_/B _4757_/B vssd1 vssd1 vccd1 vccd1 _4757_/Y sky130_fd_sc_hd__nor2_8
XFILLER_0_7_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3708_ _3473_/A _3697_/X _3674_/A _3365_/B vssd1 vssd1 vccd1 vccd1 _3708_/Y sky130_fd_sc_hd__o211ai_4
XANTENNA__4780__C1 _5740_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4688_ _4683_/X _5240_/S _4687_/Y vssd1 vssd1 vccd1 vccd1 _4688_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_70_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3639_ _3639_/A _3639_/B _3639_/C _3630_/X vssd1 vssd1 vccd1 vccd1 _3641_/B sky130_fd_sc_hd__or4b_1
X_6427_ _6428_/CLK _6427_/D fanout172/X vssd1 vssd1 vccd1 vccd1 _6427_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__3335__A0 _4255_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6358_ _6408_/CLK hold30/X vssd1 vssd1 vccd1 vccd1 hold29/A sky130_fd_sc_hd__dfxtp_1
X_5309_ _5077_/A _4216_/B _5308_/X _4639_/B vssd1 vssd1 vccd1 vccd1 _5309_/X sky130_fd_sc_hd__a211o_1
X_6289_ _6290_/CLK _6289_/D fanout167/X vssd1 vssd1 vccd1 vccd1 _6289_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__5712__S _6064_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4835__A0 _6322_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_21_wb_clk_i _6404_/CLK vssd1 vssd1 vccd1 vccd1 _6406_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_93_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5157__B1_N _5242_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5866__A2 _6380_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4 hold4/A vssd1 vssd1 vccd1 vccd1 hold4/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4826__B1 _5728_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3990_ _4040_/A _5205_/B _3986_/X _3989_/X vssd1 vssd1 vccd1 vccd1 _3990_/X sky130_fd_sc_hd__a211o_1
XANTENNA__4054__B2 _4427_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5660_ _6133_/Q _4198_/B _5676_/B1 _6212_/Q _5676_/C1 vssd1 vssd1 vccd1 vccd1 _5661_/B
+ sky130_fd_sc_hd__o221a_1
XANTENNA__3097__B _4685_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4611_ _4616_/A hold359/X _5728_/A hold673/X vssd1 vssd1 vccd1 vccd1 _5372_/B sky130_fd_sc_hd__a211o_1
XANTENNA__5003__B1 _5060_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6059__A2_N _6063_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5591_ _6136_/Q _4198_/B _5676_/B1 _6091_/Q _5675_/C1 vssd1 vssd1 vccd1 vccd1 _5597_/C
+ sky130_fd_sc_hd__a221o_1
X_4542_ _4541_/C _5733_/A _3770_/A _4541_/X vssd1 vssd1 vccd1 vccd1 _4542_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_80_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4701__S _4731_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5306__A1 _5715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold426 _5684_/X vssd1 vssd1 vccd1 vccd1 _6342_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4473_ _4427_/X hold241/X _4473_/S vssd1 vssd1 vccd1 vccd1 _4473_/X sky130_fd_sc_hd__mux2_1
Xhold404 _5030_/X vssd1 vssd1 vccd1 vccd1 _6288_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold415 _6023_/X vssd1 vssd1 vccd1 vccd1 _6439_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3317__B1 _3369_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3424_ _4309_/A _5728_/B vssd1 vssd1 vccd1 vccd1 _3424_/X sky130_fd_sc_hd__and2_1
Xhold459 _6239_/Q vssd1 vssd1 vccd1 vccd1 hold459/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold448 _5068_/X vssd1 vssd1 vccd1 vccd1 _6290_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6212_ _6412_/CLK _6212_/D vssd1 vssd1 vccd1 vccd1 _6212_/Q sky130_fd_sc_hd__dfxtp_1
Xhold437 _6434_/Q vssd1 vssd1 vccd1 vccd1 hold437/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3355_ _3431_/A _5359_/B _4346_/B vssd1 vssd1 vccd1 vccd1 _3357_/D sky130_fd_sc_hd__o21a_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6143_ _6355_/CLK _6143_/D vssd1 vssd1 vccd1 vccd1 _6143_/Q sky130_fd_sc_hd__dfxtp_1
X_3286_ _3290_/B _3220_/A _3379_/B _3091_/X vssd1 vssd1 vccd1 vccd1 _3367_/B sky130_fd_sc_hd__o22a_2
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6074_ _6221_/CLK _6074_/D vssd1 vssd1 vccd1 vccd1 _6074_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5025_ _6365_/Q _5024_/X _5927_/S vssd1 vssd1 vccd1 vccd1 _5025_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5927_ _6367_/Q _6386_/Q _5927_/S vssd1 vssd1 vccd1 vccd1 _5927_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_48_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5858_ _5858_/A _5858_/B vssd1 vssd1 vccd1 vccd1 _5858_/Y sky130_fd_sc_hd__xnor2_1
X_4809_ _4809_/A _4809_/B _4905_/C vssd1 vssd1 vccd1 vccd1 _4828_/B sky130_fd_sc_hd__or3b_1
X_5789_ _5778_/A _5742_/A _5788_/X _5731_/X vssd1 vssd1 vccd1 vccd1 _5789_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_90_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3556__B1 _4637_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3859__A1 _3850_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3751__A _3952_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4285__C _4727_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5617__S _5691_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3547__B1 _5096_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3140_ _3292_/C _3152_/A vssd1 vssd1 vccd1 vccd1 _3186_/B sky130_fd_sc_hd__nand2_2
XANTENNA__4275__B2 _3656_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3071_ _4633_/B vssd1 vssd1 vccd1 vccd1 _5989_/B sky130_fd_sc_hd__inv_2
XFILLER_0_89_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4027__A1 _6247_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5588__A _5603_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4492__A _4510_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5775__A1 _5932_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3973_ _3973_/A _3973_/B vssd1 vssd1 vccd1 vccd1 _3973_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_85_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5712_ hold27/X _4094_/Y _6064_/S vssd1 vssd1 vccd1 vccd1 hold28/A sky130_fd_sc_hd__mux2_1
XANTENNA__5775__B2 _5747_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5527__A1 _6057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5643_ _6270_/Q _5589_/X _5610_/X hold411/X _5642_/X vssd1 vssd1 vccd1 vccd1 _5644_/B
+ sky130_fd_sc_hd__a221o_1
X_5574_ _5574_/A _5574_/B vssd1 vssd1 vccd1 vccd1 _5574_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__4431__S _4437_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4525_ hold453/X _6268_/Q _4539_/S vssd1 vssd1 vccd1 vccd1 _4525_/X sky130_fd_sc_hd__mux2_1
Xhold201 _6075_/Q vssd1 vssd1 vccd1 vccd1 hold201/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold212 _6219_/Q vssd1 vssd1 vccd1 vccd1 hold212/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold234 _4448_/X vssd1 vssd1 vccd1 vccd1 _6152_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold223 _4406_/X vssd1 vssd1 vccd1 vccd1 _6132_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold267 _6250_/Q vssd1 vssd1 vccd1 vccd1 _3639_/A sky130_fd_sc_hd__buf_1
Xhold256 _6119_/Q vssd1 vssd1 vccd1 vccd1 _3541_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold245 _4495_/X vssd1 vssd1 vccd1 vccd1 _6194_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold278 _6136_/Q vssd1 vssd1 vccd1 vccd1 hold278/X sky130_fd_sc_hd__dlygate4sd3_1
X_4456_ _4510_/B _5959_/B vssd1 vssd1 vccd1 vccd1 _4464_/S sky130_fd_sc_hd__or2_4
Xhold289 _6086_/Q vssd1 vssd1 vccd1 vccd1 hold289/X sky130_fd_sc_hd__dlygate4sd3_1
X_3407_ _6389_/Q _4558_/A vssd1 vssd1 vccd1 vccd1 _3409_/B sky130_fd_sc_hd__nor2_1
X_4387_ _6314_/Q _4197_/B _5675_/C1 _4384_/X _4383_/X vssd1 vssd1 vccd1 vccd1 _4387_/X
+ sky130_fd_sc_hd__a221o_1
X_6126_ _6406_/CLK _6126_/D fanout180/X vssd1 vssd1 vccd1 vccd1 _6126_/Q sky130_fd_sc_hd__dfstp_1
X_3338_ _3290_/B _3220_/A _3337_/Y _3654_/A vssd1 vssd1 vccd1 vccd1 _3339_/B sky130_fd_sc_hd__o31a_1
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3269_ _4309_/A _4222_/B _3267_/Y _3725_/C _5560_/A vssd1 vssd1 vccd1 vccd1 _3269_/X
+ sky130_fd_sc_hd__a41o_1
X_6057_ _6057_/A _6057_/B _6057_/C vssd1 vssd1 vccd1 vccd1 _6057_/X sky130_fd_sc_hd__or3_1
X_5008_ _6331_/Q _5928_/A2 _5928_/B1 _5007_/X vssd1 vssd1 vccd1 vccd1 _5008_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_95_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4341__S _4345_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_21_wb_clk_i_A _6404_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4516__S _4518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3656__A _3656_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6032__A _6032_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3094__C _3254_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5290_ _4214_/B _5578_/B _5288_/Y _5289_/Y _3196_/B vssd1 vssd1 vccd1 vccd1 _5293_/B
+ sky130_fd_sc_hd__a311o_1
X_4310_ _4316_/B _4310_/B _4310_/C vssd1 vssd1 vccd1 vccd1 _4310_/X sky130_fd_sc_hd__or3_1
XFILLER_0_2_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4241_ _3572_/Y _3666_/A _4240_/Y _4238_/Y vssd1 vssd1 vccd1 vccd1 _4568_/B sky130_fd_sc_hd__a31o_2
X_4172_ _4171_/X _4172_/B _4172_/C vssd1 vssd1 vccd1 vccd1 _4172_/X sky130_fd_sc_hd__and3b_1
X_3123_ _3334_/C _3292_/C vssd1 vssd1 vccd1 vccd1 _3243_/B sky130_fd_sc_hd__nand2_1
X_3054_ _6243_/Q vssd1 vssd1 vccd1 vccd1 _3886_/A sky130_fd_sc_hd__inv_2
XANTENNA__5996__B2 _5365_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3330__S _6297_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3956_ _3746_/X _3953_/B _3955_/X _3951_/X vssd1 vssd1 vccd1 vccd1 _3956_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_73_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4420__B2 _4427_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3887_ _3885_/B _3887_/B vssd1 vssd1 vccd1 vccd1 _3889_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_91_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3566__A _3566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5626_ _5626_/A _5626_/B vssd1 vssd1 vccd1 vccd1 _5626_/X sky130_fd_sc_hd__or2_1
XFILLER_0_33_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5557_ hold526/X _5556_/X _5557_/S vssd1 vssd1 vccd1 vccd1 _5557_/X sky130_fd_sc_hd__mux2_1
X_5488_ _6442_/Q _4938_/B _5518_/S vssd1 vssd1 vccd1 vccd1 _5489_/B sky130_fd_sc_hd__mux2_1
X_4508_ hold153/X _4420_/X _4509_/S vssd1 vssd1 vccd1 vccd1 _4508_/X sky130_fd_sc_hd__mux2_1
X_4439_ hold91/X _4367_/X _4446_/S vssd1 vssd1 vccd1 vccd1 hold92/A sky130_fd_sc_hd__mux2_1
XANTENNA__4239__A1 _3656_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3451__D _5978_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5720__S _5723_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6109_ _6217_/CLK _6109_/D vssd1 vssd1 vccd1 vccd1 _6109_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3998__B1 _3791_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4336__S _4336_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5956__A _5977_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4175__B1 _5217_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5675__B1 _5676_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3642__C _3642_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6382__RESET_B fanout168/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6311__RESET_B fanout173/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3810_ _3810_/A _3810_/B vssd1 vssd1 vccd1 vccd1 _4599_/A sky130_fd_sc_hd__nor2_2
X_4790_ _6319_/Q _5060_/S _6320_/Q vssd1 vssd1 vccd1 vccd1 _4793_/C sky130_fd_sc_hd__a21o_1
X_3741_ _6303_/Q _6301_/Q _5087_/A vssd1 vssd1 vccd1 vccd1 _3741_/X sky130_fd_sc_hd__and3_2
XFILLER_0_55_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3672_ _3482_/A _5322_/D _3661_/X _3662_/X vssd1 vssd1 vccd1 vccd1 _3672_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6391_ _6397_/CLK _6391_/D fanout172/X vssd1 vssd1 vccd1 vccd1 _6391_/Q sky130_fd_sc_hd__dfrtp_2
X_5411_ _5397_/B _5399_/B _5395_/X vssd1 vssd1 vccd1 vccd1 _5412_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_2_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5342_ _3770_/A _3273_/C _4207_/X _5315_/B vssd1 vssd1 vccd1 vccd1 _5343_/D sky130_fd_sc_hd__a211o_1
XANTENNA__3913__B1 _3791_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5273_ _5292_/B _5273_/B _5273_/C _5273_/D vssd1 vssd1 vccd1 vccd1 _5273_/X sky130_fd_sc_hd__or4_2
X_4224_ _4224_/A _5359_/A _4224_/C vssd1 vssd1 vccd1 vccd1 _5341_/B sky130_fd_sc_hd__and3_1
XANTENNA__5418__A0 _6419_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4155_ _4155_/A _4155_/B vssd1 vssd1 vccd1 vccd1 _4156_/B sky130_fd_sc_hd__or2_1
X_3106_ _3502_/A _5303_/A vssd1 vssd1 vccd1 vccd1 _3109_/B sky130_fd_sc_hd__nor2_2
XANTENNA__3692__A2 _6304_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5540__S _6060_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4086_ _4142_/S _4085_/X _4056_/X vssd1 vssd1 vccd1 vccd1 _6052_/A sky130_fd_sc_hd__a21oi_4
X_3037_ _3656_/A vssd1 vssd1 vccd1 vccd1 _3594_/A sky130_fd_sc_hd__inv_2
XFILLER_0_77_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5197__A2 _3502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4680__A _5931_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4988_ _6330_/Q _5928_/A2 _5928_/B1 _4987_/X vssd1 vssd1 vccd1 vccd1 _4988_/X sky130_fd_sc_hd__a22o_1
X_3939_ _3939_/A _3939_/B vssd1 vssd1 vccd1 vccd1 _3940_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_80_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5609_ _5695_/A1 hold496/X _5571_/Y _5608_/X vssd1 vssd1 vccd1 vccd1 _5609_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_46_wb_clk_i clkbuf_leaf_6_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6331_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_14_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5016__A _5054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold474_A _6340_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold641_A _6419_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4574__B _4604_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5593__C1 _3721_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5896__A0 _6420_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4699__A1 _6269_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4699__B2 _5371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3653__B _5931_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4871__B2 _5061_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4871__A1 _6421_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5960_ _4367_/X hold302/X _5967_/S vssd1 vssd1 vccd1 vccd1 _5960_/X sky130_fd_sc_hd__mux2_1
X_5891_ _5847_/X _5858_/A _5889_/Y _5890_/X vssd1 vssd1 vccd1 vccd1 _5892_/B sky130_fd_sc_hd__a31o_1
XANTENNA_clkbuf_2_0__f_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4911_ _6326_/Q _4910_/X _5849_/S vssd1 vssd1 vccd1 vccd1 _4911_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_7_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4842_ _6164_/Q _6172_/Q _6411_/Q _6180_/Q _5051_/S0 _5052_/S1 vssd1 vssd1 vccd1
+ vccd1 _4842_/X sky130_fd_sc_hd__mux4_1
X_4773_ _4768_/A _4766_/Y _4768_/B _4772_/Y _4639_/B vssd1 vssd1 vccd1 vccd1 _4774_/B
+ sky130_fd_sc_hd__a41o_1
XANTENNA__4387__B1 _5675_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3724_ _3724_/A vssd1 vssd1 vccd1 vccd1 _4424_/A sky130_fd_sc_hd__inv_2
X_3655_ _3661_/A _3654_/X _5560_/A vssd1 vssd1 vccd1 vccd1 _3655_/Y sky130_fd_sc_hd__a21oi_2
X_6443_ _6447_/CLK _6443_/D fanout171/X vssd1 vssd1 vccd1 vccd1 _6443_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_0_70_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3586_ _3224_/X _3501_/B _4346_/B vssd1 vssd1 vccd1 vccd1 _3586_/X sky130_fd_sc_hd__a21o_1
XANTENNA_fanout108_A _5347_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6374_ _6374_/CLK _6374_/D fanout169/X vssd1 vssd1 vccd1 vccd1 _6374_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__4785__S1 _5358_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5325_ _5325_/A _5360_/C vssd1 vssd1 vccd1 vccd1 _5326_/D sky130_fd_sc_hd__nand2_1
XFILLER_0_11_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5256_ _5256_/A _5256_/B vssd1 vssd1 vccd1 vccd1 _5256_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_54_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4207_ _4541_/A _4223_/B _3109_/B _4541_/D _3553_/Y vssd1 vssd1 vccd1 vccd1 _4207_/X
+ sky130_fd_sc_hd__a32o_1
X_5187_ _6237_/Q _4520_/Y _5076_/Y _5078_/Y vssd1 vssd1 vccd1 vccd1 _5187_/X sky130_fd_sc_hd__a2bb2o_1
X_4138_ _4255_/B _3746_/X _4137_/X _6342_/Q vssd1 vssd1 vccd1 vccd1 _4138_/X sky130_fd_sc_hd__a22o_1
X_6065__2 _6406_/CLK vssd1 vssd1 vccd1 vccd1 _6123_/CLK sky130_fd_sc_hd__inv_2
X_4069_ _4070_/A _5126_/B vssd1 vssd1 vccd1 vccd1 _4179_/A sky130_fd_sc_hd__nor2_1
XANTENNA__4090__A2 _3784_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5590__A2 _4198_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3473__B _3473_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout160 hold614/X vssd1 vssd1 vccd1 vccd1 _3530_/D sky130_fd_sc_hd__buf_4
Xfanout171 fanout181/X vssd1 vssd1 vccd1 vccd1 fanout171/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__5180__S _5243_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4605__B2 _6274_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4605__A1 _6423_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold608 _6322_/Q vssd1 vssd1 vccd1 vccd1 hold608/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3440_ _5981_/B vssd1 vssd1 vccd1 vccd1 _3440_/Y sky130_fd_sc_hd__inv_2
XANTENNA__6040__A _6040_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold619 _6274_/Q vssd1 vssd1 vccd1 vccd1 hold619/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3371_ _3483_/A _3600_/C _3511_/A _3371_/D vssd1 vssd1 vccd1 vccd1 _3376_/B sky130_fd_sc_hd__or4_1
X_5110_ _5110_/A _5206_/B vssd1 vssd1 vccd1 vccd1 _5114_/A sky130_fd_sc_hd__xor2_1
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6090_ _6433_/CLK _6090_/D vssd1 vssd1 vccd1 vccd1 _6090_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4198__C _4427_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5041_ _5059_/B _5041_/B vssd1 vssd1 vccd1 vccd1 _5041_/Y sky130_fd_sc_hd__nor2_1
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4844__A1 _5054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
XANTENNA__6046__B1 _6057_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5943_ _3081_/Y _5936_/B _5937_/Y _5096_/A _5952_/A vssd1 vssd1 vccd1 vccd1 _5943_/X
+ sky130_fd_sc_hd__a32o_1
X_5874_ _5932_/S _5869_/Y _5873_/X _5747_/A vssd1 vssd1 vccd1 vccd1 _5874_/X sky130_fd_sc_hd__o22a_1
XANTENNA__4434__S _4437_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4825_ _4824_/X _4823_/X _5053_/S vssd1 vssd1 vccd1 vccd1 _4830_/B sky130_fd_sc_hd__mux2_4
XFILLER_0_90_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5309__C1 _4639_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4756_ _4756_/A _4758_/C _4757_/B vssd1 vssd1 vccd1 vccd1 _4756_/Y sky130_fd_sc_hd__nor3_4
XANTENNA__3574__A _5096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3707_ hold21/A _4391_/A2 _4382_/C vssd1 vssd1 vccd1 vccd1 _3707_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_43_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4687_ _5240_/S _4686_/X _4731_/S vssd1 vssd1 vccd1 vccd1 _4687_/Y sky130_fd_sc_hd__o21ai_1
X_3638_ _3638_/A _3641_/A _3638_/C vssd1 vssd1 vccd1 vccd1 _3638_/X sky130_fd_sc_hd__and3_1
X_6426_ _6428_/CLK _6426_/D fanout172/X vssd1 vssd1 vccd1 vccd1 _6426_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3569_ _3482_/A _3568_/X _5320_/B vssd1 vssd1 vccd1 vccd1 _3569_/Y sky130_fd_sc_hd__a21oi_1
X_6357_ _6444_/CLK hold28/X vssd1 vssd1 vccd1 vccd1 hold27/A sky130_fd_sc_hd__dfxtp_1
X_5308_ _5277_/Y _5313_/A vssd1 vssd1 vccd1 vccd1 _5308_/X sky130_fd_sc_hd__and2b_1
X_6288_ _6290_/CLK _6288_/D fanout167/X vssd1 vssd1 vccd1 vccd1 _6288_/Q sky130_fd_sc_hd__dfrtp_4
X_5239_ _6240_/Q _6298_/Q _5239_/S vssd1 vssd1 vccd1 vccd1 _5239_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_98_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4344__S _4345_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4771__B1 _4637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3484__A _5560_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4299__B _5739_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5079__A1 _4070_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4826__A1 _5054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5 hold5/A vssd1 vssd1 vccd1 vccd1 hold5/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3801__A2 _3784_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4610_ _3639_/A _4609_/X _6405_/Q vssd1 vssd1 vccd1 vccd1 _4610_/X sky130_fd_sc_hd__o21ba_1
X_5590_ _6068_/Q _4198_/B _5676_/B1 _6192_/Q _5676_/C1 vssd1 vssd1 vccd1 vccd1 _5590_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4762__A0 _5365_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4541_ _4541_/A _4541_/B _4541_/C _4541_/D vssd1 vssd1 vccd1 vccd1 _4541_/X sky130_fd_sc_hd__and4_1
XFILLER_0_52_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold427 _6283_/Q vssd1 vssd1 vccd1 vccd1 hold427/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold405 _6366_/Q vssd1 vssd1 vccd1 vccd1 hold405/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold416 _6362_/Q vssd1 vssd1 vccd1 vccd1 hold416/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4472_ _4420_/X hold81/X _4473_/S vssd1 vssd1 vccd1 vccd1 hold82/A sky130_fd_sc_hd__mux2_1
X_3423_ _3686_/A _3389_/Y _3421_/X _3422_/X vssd1 vssd1 vccd1 vccd1 _3436_/B sky130_fd_sc_hd__a31oi_2
Xhold449 _6316_/Q vssd1 vssd1 vccd1 vccd1 _3363_/B sky130_fd_sc_hd__buf_1
X_6211_ _6413_/CLK _6211_/D vssd1 vssd1 vccd1 vccd1 _6211_/Q sky130_fd_sc_hd__dfxtp_1
Xhold438 _6003_/X vssd1 vssd1 vccd1 vccd1 _6434_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6142_ _6181_/CLK _6142_/D vssd1 vssd1 vccd1 vccd1 _6142_/Q sky130_fd_sc_hd__dfxtp_1
X_3354_ _3611_/A _3632_/B vssd1 vssd1 vccd1 vccd1 _5359_/B sky130_fd_sc_hd__nor2_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3285_ _3290_/B _3285_/B vssd1 vssd1 vccd1 vccd1 _4550_/B sky130_fd_sc_hd__or2_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6073_ _6354_/CLK _6073_/D vssd1 vssd1 vccd1 vccd1 _6073_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5024_ _6384_/Q _4754_/X _5018_/X _5023_/X vssd1 vssd1 vccd1 vccd1 _5024_/X sky130_fd_sc_hd__a211o_1
XANTENNA_fanout175_A fanout178/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5242__A1 _6423_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5926_ _5926_/A _5926_/B vssd1 vssd1 vccd1 vccd1 _5926_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_61_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5857_ _5845_/A _5926_/A _5847_/X vssd1 vssd1 vccd1 vccd1 _5858_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_35_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_11_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_8_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4202__C1 _5675_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4808_ _6321_/Q _4827_/C vssd1 vssd1 vccd1 vccd1 _4808_/X sky130_fd_sc_hd__or2_1
X_5788_ _5932_/S _5783_/X _5787_/X _5747_/A vssd1 vssd1 vccd1 vccd1 _5788_/X sky130_fd_sc_hd__o22a_1
X_4739_ _6184_/Q _6128_/Q hold91/A _6207_/Q _4326_/B _5358_/A0 vssd1 vssd1 vccd1 vccd1
+ _4739_/X sky130_fd_sc_hd__mux4_1
X_6409_ _6414_/CLK _6409_/D vssd1 vssd1 vccd1 vccd1 _6409_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5723__S _5723_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout88_A _3642_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4847__B _4867_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3751__B _4070_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4339__S _4345_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4863__A _5054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_50_wb_clk_i_A clkbuf_leaf_6_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__3198__B _4679_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4419__S0 _5673_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3070_ _3070_/A vssd1 vssd1 vccd1 vccd1 _5988_/C sky130_fd_sc_hd__inv_2
XFILLER_0_89_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3972_ _3942_/A _3942_/B _3938_/B vssd1 vssd1 vccd1 vccd1 _3973_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_85_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5711_ hold17/X _4020_/B _6064_/S vssd1 vssd1 vccd1 vccd1 hold18/A sky130_fd_sc_hd__mux2_1
XFILLER_0_45_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5642_ _6382_/Q _5600_/X _5639_/X _5594_/Y vssd1 vssd1 vccd1 vccd1 _5642_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_31_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5573_ _3686_/A _4222_/B _4255_/Y _4247_/X vssd1 vssd1 vccd1 vccd1 _5573_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_72_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4735__B1 _6389_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4524_ hold486/X _6267_/Q _4539_/S vssd1 vssd1 vccd1 vccd1 _4524_/X sky130_fd_sc_hd__mux2_1
Xhold202 _4206_/X vssd1 vssd1 vccd1 vccd1 _6075_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold224 _6072_/Q vssd1 vssd1 vccd1 vccd1 hold224/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold235 _6156_/Q vssd1 vssd1 vccd1 vccd1 hold235/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold213 _4515_/X vssd1 vssd1 vccd1 vccd1 _6219_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold268 _5958_/X vssd1 vssd1 vccd1 vccd1 _6405_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold246 _6113_/Q vssd1 vssd1 vccd1 vccd1 hold246/X sky130_fd_sc_hd__dlygate4sd3_1
X_4455_ _4205_/X hold149/X _4455_/S vssd1 vssd1 vccd1 vccd1 _4455_/X sky130_fd_sc_hd__mux2_1
Xhold257 _6172_/Q vssd1 vssd1 vccd1 vccd1 hold257/X sky130_fd_sc_hd__dlygate4sd3_1
X_3406_ _3572_/A _4270_/B _3384_/Y _4639_/C _3405_/Y vssd1 vssd1 vccd1 vccd1 _3406_/Y
+ sky130_fd_sc_hd__a221oi_1
X_4386_ _6409_/Q _4382_/B _4384_/S _6178_/Q _5675_/C1 vssd1 vssd1 vccd1 vccd1 _4386_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_0_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold279 _4430_/X vssd1 vssd1 vccd1 vccd1 _6136_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3337_ _3337_/A _3337_/B vssd1 vssd1 vccd1 vccd1 _3337_/Y sky130_fd_sc_hd__nand2_1
X_6125_ _6125_/CLK _6125_/D fanout176/X vssd1 vssd1 vccd1 vccd1 _6125_/Q sky130_fd_sc_hd__dfstp_1
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4266__A2 _5315_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3268_ _4255_/B _5258_/B vssd1 vssd1 vccd1 vccd1 _3725_/C sky130_fd_sc_hd__or2_1
X_6056_ _6057_/B _6056_/B vssd1 vssd1 vccd1 vccd1 _6056_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__5463__A1 _4900_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4897__S0 _6318_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3199_ _3379_/B _3628_/B vssd1 vssd1 vccd1 vccd1 _4318_/B sky130_fd_sc_hd__nor2_2
X_5007_ _6364_/Q _5006_/X _5927_/S vssd1 vssd1 vccd1 vccd1 _5007_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_95_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3226__B1 _3566_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5909_ _5909_/A _5909_/B vssd1 vssd1 vccd1 vccd1 _5909_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__5718__S _5723_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold671_A _6256_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3701__A1 _4197_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5628__S _5691_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3656__B _5322_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4717__A0 hold534/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6032__B _6063_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4240_ _3132_/B _5341_/B _4239_/X vssd1 vssd1 vccd1 vccd1 _4240_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_77_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4171_ _5217_/A _5142_/A _4171_/S vssd1 vssd1 vccd1 vccd1 _4171_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5693__B2 _6423_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5693__A1 _6386_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3122_ _3254_/A _3534_/B _3121_/Y _3136_/B vssd1 vssd1 vccd1 vccd1 _3122_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_93_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3053_ _5088_/B vssd1 vssd1 vccd1 vccd1 _5087_/A sky130_fd_sc_hd__inv_2
XANTENNA__5445__B2 _5740_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4879__S0 _5358_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4707__S _4731_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6258__RESET_B fanout179/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3955_ _3758_/Y _5209_/B _3954_/X _6338_/Q vssd1 vssd1 vccd1 vccd1 _3955_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5538__S _5557_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4442__S _4446_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3886_ _3886_/A _3886_/B vssd1 vssd1 vccd1 vccd1 _3887_/B sky130_fd_sc_hd__nand2_1
XANTENNA__3566__B _3566_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5625_ _6093_/Q _4198_/B _5676_/B1 _6138_/Q _5676_/C1 vssd1 vssd1 vccd1 vccd1 _5626_/B
+ sky130_fd_sc_hd__o221a_1
XANTENNA__4184__A1 _4679_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5556_ hold526/X _5377_/X _5555_/Y _5441_/A vssd1 vssd1 vccd1 vccd1 _5556_/X sky130_fd_sc_hd__a22o_1
X_4507_ hold189/X _4412_/X _4509_/S vssd1 vssd1 vccd1 vccd1 _4507_/X sky130_fd_sc_hd__mux2_1
X_5487_ _5485_/X _5486_/X _3046_/A hold522/X vssd1 vssd1 vccd1 vccd1 _5487_/X sky130_fd_sc_hd__a2bb2o_1
X_4438_ _4438_/A _5959_/B vssd1 vssd1 vccd1 vccd1 _4446_/S sky130_fd_sc_hd__nor2_4
XANTENNA__5684__A1 _5695_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4369_ _6185_/Q _4382_/B _4382_/C vssd1 vssd1 vccd1 vccd1 _4369_/X sky130_fd_sc_hd__or3_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6108_ _6194_/CLK _6108_/D vssd1 vssd1 vccd1 vccd1 _6108_/Q sky130_fd_sc_hd__dfxtp_1
X_6039_ _6057_/A _6038_/X _6063_/S vssd1 vssd1 vccd1 vccd1 _6039_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_68_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5956__B _5956_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4175__A1 _6248_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6123__SET_B fanout180/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3642__D _4222_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3740_ _6303_/Q _3740_/B vssd1 vssd1 vccd1 vccd1 _3740_/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_27_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3610__B1 _4309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3671_ _5097_/B _4745_/B _3553_/Y _3164_/Y vssd1 vssd1 vccd1 vccd1 _3671_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_12_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6390_ _6397_/CLK _6390_/D fanout172/X vssd1 vssd1 vccd1 vccd1 _6390_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_23_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5410_ _5410_/A _5410_/B vssd1 vssd1 vccd1 vccd1 _5412_/A sky130_fd_sc_hd__nand2_1
X_5341_ _5341_/A _5341_/B _5316_/X vssd1 vssd1 vccd1 vccd1 _5341_/X sky130_fd_sc_hd__or3b_1
XFILLER_0_2_334 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5272_ _5272_/A _5272_/B _5272_/C _5272_/D vssd1 vssd1 vccd1 vccd1 _5273_/D sky130_fd_sc_hd__or4_1
XANTENNA__5666__B2 _6421_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5666__A1 _6296_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4223_ _4541_/A _4223_/B _5096_/D vssd1 vssd1 vccd1 vccd1 _5341_/A sky130_fd_sc_hd__and3_1
XANTENNA__3677__B1 _5097_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4154_ hold201/X _3715_/X _3794_/X hold165/X _4153_/X vssd1 vssd1 vccd1 vccd1 _4155_/B
+ sky130_fd_sc_hd__a221o_1
X_3105_ _6258_/Q _6257_/Q vssd1 vssd1 vccd1 vccd1 _5303_/A sky130_fd_sc_hd__or2_4
XANTENNA__3429__B1 _4541_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4085_ _6421_/Q _4084_/X _4085_/S vssd1 vssd1 vccd1 vccd1 _4085_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4437__S _4437_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3036_ _5226_/A vssd1 vssd1 vccd1 vccd1 _4685_/A sky130_fd_sc_hd__clkinv_4
XANTENNA__4680__B _5192_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3577__A _3577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4987_ _6363_/Q _4986_/X _5927_/S vssd1 vssd1 vccd1 vccd1 _4987_/X sky130_fd_sc_hd__mux2_1
X_3938_ _3938_/A _3938_/B vssd1 vssd1 vccd1 vccd1 _3938_/X sky130_fd_sc_hd__or2_1
XFILLER_0_61_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3869_ _4111_/A _4394_/B _3868_/B vssd1 vssd1 vccd1 vccd1 _3870_/C sky130_fd_sc_hd__o21bai_1
XFILLER_0_61_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5608_ _6379_/Q _5600_/X _5603_/X _5745_/A _5607_/X vssd1 vssd1 vccd1 vccd1 _5608_/X
+ sky130_fd_sc_hd__a221o_1
X_5539_ _6421_/Q _5538_/X _5558_/S vssd1 vssd1 vccd1 vccd1 _5539_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_14_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_15_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6399_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_fanout70_A _4636_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4632__A2 _4615_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5593__B1 _3718_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4148__B2 _4427_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4810__S _6315_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5890_ _6379_/Q _6380_/Q _6381_/Q _6382_/Q _5926_/A vssd1 vssd1 vccd1 vccd1 _5890_/X
+ sky130_fd_sc_hd__o41a_1
X_4910_ _6378_/Q _4796_/B _4908_/X _4909_/X vssd1 vssd1 vccd1 vccd1 _4910_/X sky130_fd_sc_hd__o22a_1
X_4841_ hold93/A hold61/A _6132_/Q _6211_/Q _5051_/S0 _5052_/S1 vssd1 vssd1 vccd1
+ vccd1 _4841_/X sky130_fd_sc_hd__mux4_1
XANTENNA__3397__A _5096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4387__A1 _6314_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4772_ _4772_/A _4772_/B vssd1 vssd1 vccd1 vccd1 _4772_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_55_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3723_ _3611_/A _3473_/A _3611_/Y _3680_/X vssd1 vssd1 vccd1 vccd1 _3723_/X sky130_fd_sc_hd__o211a_2
X_3654_ _3654_/A _3654_/B vssd1 vssd1 vccd1 vccd1 _3654_/X sky130_fd_sc_hd__or2_1
XANTENNA__5816__S _5933_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4720__S _5447_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6442_ _6445_/CLK _6442_/D fanout171/X vssd1 vssd1 vccd1 vccd1 _6442_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_0_70_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3585_ _3606_/A _3584_/X _4309_/A vssd1 vssd1 vccd1 vccd1 _6124_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6373_ _6373_/CLK _6373_/D fanout169/X vssd1 vssd1 vccd1 vccd1 _6373_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_0_100_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5324_ _5324_/A _5324_/B _5324_/C _5324_/D vssd1 vssd1 vccd1 vccd1 _5327_/C sky130_fd_sc_hd__or4_1
XFILLER_0_2_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5255_ hold357/X _5254_/X _5255_/S vssd1 vssd1 vccd1 vccd1 _5255_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5551__S _6060_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4206_ _4205_/X hold201/X _4206_/S vssd1 vssd1 vccd1 vccd1 _4206_/X sky130_fd_sc_hd__mux2_1
X_5186_ _3573_/A _5193_/S _5746_/A _3065_/Y _4681_/X vssd1 vssd1 vccd1 vccd1 _5186_/X
+ sky130_fd_sc_hd__o311a_1
X_4137_ _4255_/B _4188_/C _4134_/Y _3746_/X vssd1 vssd1 vccd1 vccd1 _4137_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4068_ _6247_/Q _6248_/Q _4067_/B _5217_/A vssd1 vssd1 vccd1 vccd1 _5126_/B sky130_fd_sc_hd__o31a_1
XANTENNA__3283__D1 _3566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4614__A2 _5313_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3822__B1 _3791_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3100__A _3656_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4866__A _6324_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3770__A _3770_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4302__A1 _6270_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4838__C1 _5557_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout150 _6254_/Q vssd1 vssd1 vccd1 vccd1 _4284_/A sky130_fd_sc_hd__clkbuf_4
Xfanout161 _5077_/A vssd1 vssd1 vccd1 vccd1 _4767_/A sky130_fd_sc_hd__buf_4
Xfanout172 fanout173/X vssd1 vssd1 vccd1 vccd1 fanout172/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__6055__A1 _5557_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3813__B1 _3786_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold609 _5419_/X vssd1 vssd1 vccd1 vccd1 _6322_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6040__B _6063_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3370_ _4228_/A _4214_/B _3194_/A _5322_/A vssd1 vssd1 vccd1 vccd1 _3371_/D sky130_fd_sc_hd__a31o_1
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5040_ _6332_/Q _5039_/C _6333_/Q vssd1 vssd1 vccd1 vccd1 _5041_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_85_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4844__A2 _4843_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5942_ _3621_/A _3625_/B _5941_/Y _3623_/A _5096_/A vssd1 vssd1 vccd1 vccd1 _5942_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_19_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5873_ _6418_/Q _5872_/X _5930_/S vssd1 vssd1 vccd1 vccd1 _5873_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_7_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4824_ _6163_/Q _6171_/Q _6410_/Q _6179_/Q _5358_/A0 _4326_/B vssd1 vssd1 vccd1 vccd1
+ _4824_/X sky130_fd_sc_hd__mux4_1
X_4755_ _4755_/A _4757_/B vssd1 vssd1 vccd1 vccd1 _4796_/B sky130_fd_sc_hd__nand2_2
XANTENNA__5652__S0 _5691_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout120_A _6402_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3706_ _3700_/X _3704_/X _3701_/X vssd1 vssd1 vccd1 vccd1 _3863_/A sky130_fd_sc_hd__o21ai_4
XFILLER_0_7_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4450__S _4455_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4686_ hold397/X _4287_/A _4727_/S vssd1 vssd1 vccd1 vccd1 _4686_/X sky130_fd_sc_hd__mux2_1
X_3637_ _3630_/A _3635_/X _3636_/X vssd1 vssd1 vccd1 vccd1 _3637_/X sky130_fd_sc_hd__o21ba_1
X_6425_ _6430_/CLK _6425_/D fanout173/X vssd1 vssd1 vccd1 vccd1 _6425_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_3_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4532__A1 _4070_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3568_ _6293_/Q _4346_/A _5265_/B _3567_/X vssd1 vssd1 vccd1 vccd1 _3568_/X sky130_fd_sc_hd__a31o_1
X_6356_ _6445_/CLK hold18/X vssd1 vssd1 vccd1 vccd1 hold17/A sky130_fd_sc_hd__dfxtp_1
X_5307_ _5715_/B hold626/X _5283_/Y _5321_/S vssd1 vssd1 vccd1 vccd1 _5307_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_59_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3499_ _4223_/B _5258_/B _5256_/A _3549_/B _3498_/Y vssd1 vssd1 vccd1 vccd1 _3499_/X
+ sky130_fd_sc_hd__o311a_1
XANTENNA__3590__A _4679_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6287_ _6290_/CLK _6287_/D fanout166/X vssd1 vssd1 vccd1 vccd1 _6287_/Q sky130_fd_sc_hd__dfrtp_2
X_5238_ _6298_/Q _5149_/X _5237_/X _4182_/X _4188_/X vssd1 vssd1 vccd1 vccd1 _5238_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_98_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5169_ hold610/X _5447_/S _5167_/X _5168_/Y vssd1 vssd1 vccd1 vccd1 _5169_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_98_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_40_wb_clk_i_A clkbuf_leaf_6_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4360__S _4360_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_30_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6373_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__5720__A0 _6271_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5079__A2 _5193_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5191__S _5347_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4826__A2 _4830_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold6 hold6/A vssd1 vssd1 vccd1 vccd1 hold6/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5539__A0 _6421_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4540_ _4541_/C _5341_/B _5317_/A vssd1 vssd1 vccd1 vccd1 _4540_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_52_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3394__B _5322_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4471_ _4412_/X hold87/X _4473_/S vssd1 vssd1 vccd1 vccd1 hold88/A sky130_fd_sc_hd__mux2_1
Xhold406 _5722_/X vssd1 vssd1 vccd1 vccd1 _6366_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold417 _5718_/X vssd1 vssd1 vccd1 vccd1 _6362_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3422_ _5313_/A _3399_/X _3415_/B _5096_/B _5935_/A vssd1 vssd1 vccd1 vccd1 _3422_/X
+ sky130_fd_sc_hd__a221o_1
Xhold439 _6339_/Q vssd1 vssd1 vccd1 vccd1 _3992_/A sky130_fd_sc_hd__clkbuf_2
Xhold428 _4934_/X vssd1 vssd1 vccd1 vccd1 _6283_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6210_ _6410_/CLK _6210_/D vssd1 vssd1 vccd1 vccd1 _6210_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6141_ _6354_/CLK _6141_/D vssd1 vssd1 vccd1 vccd1 _6141_/Q sky130_fd_sc_hd__dfxtp_1
X_3353_ _4639_/C _5266_/B vssd1 vssd1 vccd1 vccd1 _3357_/C sky130_fd_sc_hd__or2_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3284_ _3290_/B _3285_/B vssd1 vssd1 vccd1 vccd1 _4541_/D sky130_fd_sc_hd__nor2_2
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6072_ _6218_/CLK _6072_/D vssd1 vssd1 vccd1 vccd1 _6072_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5023_ _5061_/A1 _5020_/X _5022_/X _4867_/B vssd1 vssd1 vccd1 vccd1 _5023_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_95_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout168_A fanout181/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4445__S _4446_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5925_ _5925_/A _5925_/B vssd1 vssd1 vccd1 vccd1 _5926_/B sky130_fd_sc_hd__xor2_1
X_5856_ _5856_/A _5926_/A vssd1 vssd1 vccd1 vccd1 _5858_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_298 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4807_ _4806_/X _4805_/X _5053_/S vssd1 vssd1 vccd1 vccd1 _4807_/X sky130_fd_sc_hd__mux2_4
XFILLER_0_8_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5787_ _6322_/Q _5852_/S _5786_/X vssd1 vssd1 vccd1 vccd1 _5787_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_9_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4738_ _5728_/D vssd1 vssd1 vccd1 vccd1 _4738_/Y sky130_fd_sc_hd__inv_2
X_4669_ _6338_/Q _6342_/Q _4674_/S vssd1 vssd1 vccd1 vccd1 _4669_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_43_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_7_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_6408_ _6408_/CLK _6408_/D vssd1 vssd1 vccd1 vccd1 _6408_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6339_ _6373_/CLK _6339_/D vssd1 vssd1 vccd1 vccd1 _6339_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__4269__B1 _5578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4863__B _4863_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4355__S _4360_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4419__S1 _3718_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6305__RESET_B fanout180/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5588__C _5603_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3971_ _3969_/B _3971_/B vssd1 vssd1 vccd1 vccd1 _3973_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_57_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5710_ hold9/X _4001_/B _6064_/S vssd1 vssd1 vccd1 vccd1 hold10/A sky130_fd_sc_hd__mux2_1
XFILLER_0_85_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3609__S _4309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5641_ _6436_/Q _5588_/X _5603_/X _5778_/A _5640_/X vssd1 vssd1 vccd1 vccd1 _5644_/A
+ sky130_fd_sc_hd__a221o_1
X_5572_ _5603_/B _5602_/B vssd1 vssd1 vccd1 vccd1 _5610_/A sky130_fd_sc_hd__nor2_1
X_4523_ _5740_/A _4523_/B vssd1 vssd1 vccd1 vccd1 _5239_/S sky130_fd_sc_hd__or2_2
Xhold214 _6176_/Q vssd1 vssd1 vccd1 vccd1 hold214/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold225 _4055_/X vssd1 vssd1 vccd1 vccd1 _6072_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold203 _6153_/Q vssd1 vssd1 vccd1 vccd1 hold203/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold247 _6251_/Q vssd1 vssd1 vccd1 vccd1 hold247/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold269 _6428_/Q vssd1 vssd1 vccd1 vccd1 hold269/X sky130_fd_sc_hd__dlygate4sd3_1
X_4454_ _4148_/X hold140/X _4455_/S vssd1 vssd1 vccd1 vccd1 _6158_/D sky130_fd_sc_hd__mux2_1
Xhold258 _4470_/X vssd1 vssd1 vccd1 vccd1 _6172_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold236 _6413_/Q vssd1 vssd1 vccd1 vccd1 hold236/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3405_ _4284_/C _5264_/B vssd1 vssd1 vccd1 vccd1 _3405_/Y sky130_fd_sc_hd__nor2_1
X_4385_ hold45/A _4382_/B _3718_/Y hold73/X _5673_/C1 vssd1 vssd1 vccd1 vccd1 _4385_/X
+ sky130_fd_sc_hd__o221a_1
X_3336_ _3336_/A _3336_/B _3336_/C vssd1 vssd1 vccd1 vccd1 _3337_/B sky130_fd_sc_hd__nor3_2
X_6124_ _6124_/CLK _6124_/D fanout176/X vssd1 vssd1 vccd1 vccd1 _6124_/Q sky130_fd_sc_hd__dfstp_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6055_ _5557_/S _5546_/X _6054_/B _6054_/Y vssd1 vssd1 vccd1 vccd1 _6056_/B sky130_fd_sc_hd__a31o_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3267_ _4255_/B _5258_/B vssd1 vssd1 vccd1 vccd1 _3267_/Y sky130_fd_sc_hd__nand2_1
X_5006_ _6383_/Q _4754_/X _4998_/X _5005_/X vssd1 vssd1 vccd1 vccd1 _5006_/X sky130_fd_sc_hd__a211o_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3198_ _3243_/B _4679_/D vssd1 vssd1 vccd1 vccd1 _5322_/A sky130_fd_sc_hd__nor2_2
XANTENNA__4897__S1 _6090_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3226__A1 _3278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5908_ _5888_/B _5892_/B _5888_/A vssd1 vssd1 vccd1 vccd1 _5909_/B sky130_fd_sc_hd__a21boi_2
X_5839_ _6326_/Q _5825_/S _5928_/B1 _5838_/X vssd1 vssd1 vccd1 vccd1 _5839_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_91_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5687__C1 _3721_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4965__B2 _4867_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4965__A1 _5061_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3768__A2 _6032_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4170_ _5217_/A _6248_/Q vssd1 vssd1 vccd1 vccd1 _5142_/A sky130_fd_sc_hd__xor2_1
X_3121_ _3293_/B _3549_/A vssd1 vssd1 vccd1 vccd1 _3121_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_93_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3052_ _6301_/Q vssd1 vssd1 vccd1 vccd1 _3755_/C sky130_fd_sc_hd__inv_2
XANTENNA__5599__B _5603_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4879__S1 _4326_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6434__SET_B fanout171/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3208__A1 _3278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3954_ _4188_/C _3953_/B _3953_/Y _3746_/X vssd1 vssd1 vccd1 vccd1 _3954_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_58_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4722__A1_N _6273_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3885_ _5088_/B _3885_/B vssd1 vssd1 vccd1 vccd1 _3885_/X sky130_fd_sc_hd__or2_1
XFILLER_0_85_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5624_ _6194_/Q _4198_/B _4200_/S _6070_/Q _5675_/C1 vssd1 vssd1 vccd1 vccd1 _5626_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_33_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4184__A2 _6248_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5555_ _5555_/A _5555_/B vssd1 vssd1 vccd1 vccd1 _5555_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5486_ _5553_/S _3067_/Y _5484_/B _3046_/A vssd1 vssd1 vccd1 vccd1 _5486_/X sky130_fd_sc_hd__a31o_1
X_4506_ hold177/X _4405_/X _4509_/S vssd1 vssd1 vccd1 vccd1 _4506_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4437_ hold165/X _4205_/X _4437_/S vssd1 vssd1 vccd1 vccd1 _4437_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_6_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6107_ _6266_/CLK _6107_/D fanout177/X vssd1 vssd1 vccd1 vccd1 _6107_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4368_ hold187/X _4367_/X _4428_/S vssd1 vssd1 vccd1 vccd1 _4368_/X sky130_fd_sc_hd__mux2_1
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3319_ _4637_/A _3311_/X _3318_/X _3269_/X _3304_/A vssd1 vssd1 vccd1 vccd1 _4758_/C
+ sky130_fd_sc_hd__o221a_2
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4299_ _4299_/A _5739_/A _4299_/C vssd1 vssd1 vccd1 vccd1 _4307_/B sky130_fd_sc_hd__and3_1
XANTENNA__4239__A3 _3952_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6038_ _6057_/B _4958_/B _5504_/Y _5992_/Y vssd1 vssd1 vccd1 vccd1 _6038_/X sky130_fd_sc_hd__o22a_1
XANTENNA__3998__A2 _3789_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4947__A1 _5061_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4947__B2 _4867_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5675__A2 _4198_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4635__B1 _5715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5060__A0 _6423_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3670_ _5096_/B _3663_/X _3668_/X vssd1 vssd1 vccd1 vccd1 _3674_/A sky130_fd_sc_hd__o21ai_4
XFILLER_0_12_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5363__A1 _4214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5340_ _5727_/S _5988_/C _5339_/X vssd1 vssd1 vccd1 vccd1 _5340_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__3913__A2 _3789_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5271_ _5480_/C _5322_/B _5322_/D _3367_/B vssd1 vssd1 vccd1 vccd1 _5272_/D sky130_fd_sc_hd__or4b_1
X_4222_ _3220_/A _4222_/B _4541_/B vssd1 vssd1 vccd1 vccd1 _5096_/D sky130_fd_sc_hd__and3b_2
X_4153_ _6098_/Q _3789_/X _3791_/X _6199_/Q vssd1 vssd1 vccd1 vccd1 _4153_/X sky130_fd_sc_hd__a22o_1
X_3104_ _6258_/Q _6257_/Q vssd1 vssd1 vccd1 vccd1 _3292_/C sky130_fd_sc_hd__nor2_2
X_4084_ _4040_/A _5206_/B _4079_/Y _4083_/X vssd1 vssd1 vccd1 vccd1 _4084_/X sky130_fd_sc_hd__a211o_1
XANTENNA__4626__B1 _4617_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3035_ _4284_/A vssd1 vssd1 vccd1 vccd1 _4679_/A sky130_fd_sc_hd__inv_2
XFILLER_0_93_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4453__S _4455_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6042__A2_N _6054_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4986_ _6382_/Q _4754_/X _4978_/X _4985_/X vssd1 vssd1 vccd1 vccd1 _4986_/X sky130_fd_sc_hd__a211o_1
X_3937_ _3939_/A _3939_/B vssd1 vssd1 vccd1 vccd1 _3938_/B sky130_fd_sc_hd__nor2_1
XANTENNA__3577__B _5956_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3868_ _3870_/B _3868_/B vssd1 vssd1 vccd1 vccd1 _4395_/A sky130_fd_sc_hd__nand2_1
XANTENNA__3593__A _4520_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5607_ _6416_/Q _5602_/X _5604_/X _5610_/A _5606_/X vssd1 vssd1 vccd1 vccd1 _5607_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_14_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3799_ _3799_/A vssd1 vssd1 vccd1 vccd1 _3877_/A sky130_fd_sc_hd__inv_2
X_5538_ hold577/X _5537_/X _5557_/S vssd1 vssd1 vccd1 vccd1 _5538_/X sky130_fd_sc_hd__mux2_1
X_5469_ hold590/X input7/X _5469_/S vssd1 vssd1 vccd1 vccd1 _5469_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5313__A _5313_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4617__B1 _4615_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout63_A _5772_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5042__A0 _6422_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3356__B1 _3611_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4840_ hold385/X _5068_/S _4838_/X _4839_/X vssd1 vssd1 vccd1 vccd1 _4840_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_23_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4771_ _4210_/A _5359_/A _3409_/B _4637_/A vssd1 vssd1 vccd1 vccd1 _4774_/A sky130_fd_sc_hd__a31o_1
XANTENNA__4387__A2 _4197_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3722_ hold233/X hold179/X hold97/X hold138/X _5676_/B1 _5676_/C1 vssd1 vssd1 vccd1
+ vccd1 _3722_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_99_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3653_ _3690_/B _5931_/S vssd1 vssd1 vccd1 vccd1 _6401_/D sky130_fd_sc_hd__and2_1
X_6441_ _6448_/CLK _6441_/D fanout171/X vssd1 vssd1 vccd1 vccd1 _6441_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA__3347__B1 _3309_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6372_ _6374_/CLK _6372_/D fanout170/X vssd1 vssd1 vccd1 vccd1 _6372_/Q sky130_fd_sc_hd__dfrtp_2
X_5323_ _5733_/A _5480_/C _5323_/C vssd1 vssd1 vccd1 vccd1 _5324_/D sky130_fd_sc_hd__or3_1
X_3584_ _4616_/A _3605_/B vssd1 vssd1 vccd1 vccd1 _3584_/X sky130_fd_sc_hd__or2_1
XFILLER_0_2_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5254_ _4115_/X _4157_/Y _5253_/X _5246_/Y _5221_/X vssd1 vssd1 vccd1 vccd1 _5254_/X
+ sky130_fd_sc_hd__o32a_1
X_5185_ _3065_/Y _5150_/Y _5184_/X _3755_/X vssd1 vssd1 vccd1 vccd1 _5185_/Y sky130_fd_sc_hd__o211ai_1
XANTENNA__4448__S _4455_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4205_ _4195_/X _4196_/X _4204_/X _4427_/S vssd1 vssd1 vccd1 vccd1 _4205_/X sky130_fd_sc_hd__a22o_2
XANTENNA__4311__A2 _4305_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4136_ _6248_/Q _3761_/A _5212_/A _3985_/A _4040_/A vssd1 vssd1 vccd1 vccd1 _4136_/X
+ sky130_fd_sc_hd__a221o_1
X_4067_ _6247_/Q _4067_/B vssd1 vssd1 vccd1 vccd1 _4072_/A sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_30_wb_clk_i_A clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_3_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3283__C1 _3183_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5575__B2 _4224_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4969_ _5929_/A1 _4968_/X _4958_/Y vssd1 vssd1 vccd1 vccd1 _4969_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_19_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3338__B1 _3654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout140 _3952_/A vssd1 vssd1 vccd1 vccd1 _3334_/C sky130_fd_sc_hd__buf_4
XANTENNA__3770__B _6390_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4358__S _4360_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4302__A2 _4316_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout151 _3566_/A vssd1 vssd1 vccd1 vccd1 _3289_/A sky130_fd_sc_hd__buf_4
Xfanout173 fanout174/X vssd1 vssd1 vccd1 vccd1 fanout173/X sky130_fd_sc_hd__buf_6
Xfanout162 hold614/X vssd1 vssd1 vccd1 vccd1 _5077_/A sky130_fd_sc_hd__buf_4
XANTENNA__5978__A _5978_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5263__B1 _6118_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4886__B1_N _4867_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4882__A _5054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4792__A _5060_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5941_ _5941_/A _5941_/B vssd1 vssd1 vccd1 vccd1 _5941_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__3201__A _3278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5872_ _5929_/A1 _5871_/X _4958_/Y vssd1 vssd1 vccd1 vccd1 _5872_/X sky130_fd_sc_hd__a21bo_1
Xclkbuf_leaf_0_wb_clk_i clkbuf_leaf_6_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6221_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4823_ hold41/A hold59/A _6131_/Q _6210_/Q _5358_/A0 _4326_/B vssd1 vssd1 vccd1 vccd1
+ _4823_/X sky130_fd_sc_hd__mux4_1
XANTENNA__5652__S1 _5690_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4731__S _4731_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4754_ _4755_/A _4757_/B vssd1 vssd1 vccd1 vccd1 _4754_/X sky130_fd_sc_hd__and2_4
XANTENNA__5309__A1 _5077_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3705_ _3700_/X _3704_/X _3701_/X vssd1 vssd1 vccd1 vccd1 _3850_/A sky130_fd_sc_hd__o21a_4
XFILLER_0_50_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4685_ _4685_/A _5715_/A _5226_/C vssd1 vssd1 vccd1 vccd1 _5240_/S sky130_fd_sc_hd__or3b_4
XANTENNA__4780__A2 _5728_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3636_ _3639_/A _3630_/X _3627_/Y vssd1 vssd1 vccd1 vccd1 _3636_/X sky130_fd_sc_hd__o21a_1
X_6424_ _6430_/CLK _6424_/D fanout172/X vssd1 vssd1 vccd1 vccd1 _6424_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_0_3_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3567_ _6293_/Q _5158_/A _3333_/S vssd1 vssd1 vccd1 vccd1 _3567_/X sky130_fd_sc_hd__o21a_1
X_6355_ _6355_/CLK hold10/X vssd1 vssd1 vccd1 vccd1 hold9/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5306_ _5715_/B _3938_/A _5321_/S _5305_/X vssd1 vssd1 vccd1 vccd1 _5306_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_59_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6286_ _6290_/CLK _6286_/D fanout166/X vssd1 vssd1 vccd1 vccd1 _6286_/Q sky130_fd_sc_hd__dfrtp_2
X_3498_ _6258_/Q _4223_/B _5258_/B vssd1 vssd1 vccd1 vccd1 _3498_/Y sky130_fd_sc_hd__o21ai_1
X_5237_ _3759_/A _5235_/X _5236_/X _3985_/A vssd1 vssd1 vccd1 vccd1 _5237_/X sky130_fd_sc_hd__a22o_1
X_5168_ _6040_/A _5243_/S _5447_/S vssd1 vssd1 vccd1 vccd1 _5168_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_98_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4119_ _4122_/B _4119_/B vssd1 vssd1 vccd1 vccd1 _4121_/A sky130_fd_sc_hd__and2b_1
X_5099_ _3759_/A _6292_/Q _3758_/Y _5150_/B _5102_/B vssd1 vssd1 vccd1 vccd1 _5099_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_78_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5472__S _5472_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold7 hold7/A vssd1 vssd1 vccd1 vccd1 hold7/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5236__A0 _6298_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5787__A1 _6322_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold418 _6424_/Q vssd1 vssd1 vccd1 vccd1 _5981_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4470_ _4405_/X hold257/X _4473_/S vssd1 vssd1 vccd1 vccd1 _4470_/X sky130_fd_sc_hd__mux2_1
Xhold407 _6080_/Q vssd1 vssd1 vccd1 vccd1 _3073_/A sky130_fd_sc_hd__dlygate4sd3_1
X_3421_ _3385_/Y _3387_/X _3417_/Y _3418_/Y _3420_/X vssd1 vssd1 vccd1 vccd1 _3421_/X
+ sky130_fd_sc_hd__a2111o_1
Xhold429 _6242_/Q vssd1 vssd1 vccd1 vccd1 hold429/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3352_ _4346_/A _4208_/B _5158_/A vssd1 vssd1 vccd1 vccd1 _5266_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__5382__S _6427_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6140_ _6218_/CLK _6140_/D vssd1 vssd1 vccd1 vccd1 _6140_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3283_ _3254_/A _3573_/A _4214_/B _3183_/B _3566_/A vssd1 vssd1 vccd1 vccd1 _3658_/B
+ sky130_fd_sc_hd__o2111ai_4
XANTENNA__4278__A1 _3566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6071_ _6354_/CLK _6071_/D vssd1 vssd1 vccd1 vccd1 _6071_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5022_ _6421_/Q _5021_/X _5060_/S vssd1 vssd1 vccd1 vccd1 _5022_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4726__S _5447_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5924_ _5915_/B _5917_/B _5915_/A vssd1 vssd1 vccd1 vccd1 _5925_/B sky130_fd_sc_hd__a21bo_1
X_5855_ _5845_/A _5854_/X _5933_/S vssd1 vssd1 vccd1 vccd1 _5855_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_63_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4806_ _6162_/Q hold43/A _6409_/Q _6178_/Q _5358_/A0 _4326_/B vssd1 vssd1 vccd1 vccd1
+ _4806_/X sky130_fd_sc_hd__mux4_1
XANTENNA__5557__S _5557_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4461__S _4464_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5786_ _5773_/A _5785_/X _4826_/X vssd1 vssd1 vccd1 vccd1 _5786_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_90_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4737_ _4767_/A _4736_/X _3631_/Y vssd1 vssd1 vccd1 vccd1 _5728_/D sky130_fd_sc_hd__a21o_4
XFILLER_0_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4668_ _6022_/A _4673_/B vssd1 vssd1 vccd1 vccd1 _4668_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_9_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3619_ _3619_/A _3619_/B vssd1 vssd1 vccd1 vccd1 _3620_/B sky130_fd_sc_hd__nor2_1
X_6407_ _6407_/CLK _6407_/D vssd1 vssd1 vccd1 vccd1 _6407_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4599_ _4599_/A _4604_/S vssd1 vssd1 vccd1 vccd1 _4599_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_101_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6338_ _6374_/CLK _6338_/D vssd1 vssd1 vccd1 vccd1 _6338_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__4269__A1 _4685_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3106__A _3502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6269_ _6271_/CLK _6269_/D fanout170/X vssd1 vssd1 vccd1 vccd1 _6269_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__4364__S1 _5673_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4441__A1 _4392_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3970_ _3970_/A _3970_/B vssd1 vssd1 vccd1 vccd1 _3971_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_15_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5640_ _6294_/Q _5587_/X _5602_/X _6419_/Q vssd1 vssd1 vccd1 vccd1 _5640_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_26_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5571_ _5571_/A vssd1 vssd1 vccd1 vccd1 _5571_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_5_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4196__B1 _5597_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4522_ _5560_/A _4522_/B _5303_/A _4522_/D vssd1 vssd1 vccd1 vccd1 _4523_/B sky130_fd_sc_hd__or4_2
XFILLER_0_25_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold215 _4475_/X vssd1 vssd1 vccd1 vccd1 _6176_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold226 _6140_/Q vssd1 vssd1 vccd1 vccd1 hold226/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold204 _4449_/X vssd1 vssd1 vccd1 vccd1 _6153_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4453_ _4102_/X hold85/X _4455_/S vssd1 vssd1 vccd1 vccd1 hold86/A sky130_fd_sc_hd__mux2_1
XFILLER_0_13_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold248 _4618_/X vssd1 vssd1 vccd1 vccd1 _6251_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3404_ _5264_/B vssd1 vssd1 vccd1 vccd1 _3404_/Y sky130_fd_sc_hd__inv_2
Xhold237 _5966_/X vssd1 vssd1 vccd1 vccd1 _6413_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5406__A _5715_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold259 _6135_/Q vssd1 vssd1 vccd1 vccd1 hold259/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4384_ hold43/A _6162_/Q _4384_/S vssd1 vssd1 vccd1 vccd1 _4384_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_21_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4310__A _4316_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6123_ _6123_/CLK _6127_/D fanout180/X vssd1 vssd1 vccd1 vccd1 _6123_/Q sky130_fd_sc_hd__dfstp_1
X_3335_ _4255_/B _5328_/C _6298_/Q vssd1 vssd1 vccd1 vccd1 _3336_/C sky130_fd_sc_hd__mux2_1
XFILLER_0_0_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3266_ _3260_/Y _3264_/X _3265_/X _4637_/A vssd1 vssd1 vccd1 vccd1 _3304_/B sky130_fd_sc_hd__a31o_1
X_6054_ _6054_/A _6054_/B vssd1 vssd1 vccd1 vccd1 _6054_/Y sky130_fd_sc_hd__nor2_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5999__A1 _5339_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6086__RESET_B fanout174/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5005_ _5061_/A1 _5000_/X _5004_/X _4867_/B vssd1 vssd1 vccd1 vccd1 _5005_/X sky130_fd_sc_hd__a22o_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3197_ _3197_/A _3197_/B _3197_/C vssd1 vssd1 vccd1 vccd1 _3247_/A sky130_fd_sc_hd__or3_1
XANTENNA__5141__A _6246_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout180_A fanout181/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3226__A2 _3369_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5907_ _5907_/A _5907_/B vssd1 vssd1 vccd1 vccd1 _5909_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_91_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5838_ _6326_/Q _6378_/Q _5849_/S vssd1 vssd1 vccd1 vccd1 _5838_/X sky130_fd_sc_hd__mux2_1
X_5769_ _5769_/A _5769_/B _5767_/X vssd1 vssd1 vccd1 vccd1 _5770_/B sky130_fd_sc_hd__or3b_1
XANTENNA__6122__D _6126_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4220__A _5317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4662__A1 _5715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3217__A2 _3502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3925__B1 _3786_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5226__A _5226_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3120_ _3289_/A _3549_/A vssd1 vssd1 vccd1 vccd1 _3534_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_93_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3051_ _6304_/Q vssd1 vssd1 vccd1 vccd1 _3759_/A sky130_fd_sc_hd__inv_2
XANTENNA__6057__A _6057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4405__B2 _4427_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3953_ _4134_/B _3953_/B vssd1 vssd1 vccd1 vccd1 _3953_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_73_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3884_ _3886_/A _3886_/B vssd1 vssd1 vccd1 vccd1 _3885_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_18_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5623_ _6293_/Q _5587_/X _5600_/X _6381_/Q _5622_/X vssd1 vssd1 vccd1 vccd1 _5631_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_5_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3392__A1 _3337_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5554_ _5554_/A _5554_/B vssd1 vssd1 vccd1 vccd1 _5555_/B sky130_fd_sc_hd__xor2_1
XANTENNA__3392__B2 _3654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5485_ _4313_/C _5377_/A _5478_/Y _5479_/Y _5558_/S vssd1 vssd1 vccd1 vccd1 _5485_/X
+ sky130_fd_sc_hd__o311a_1
X_4505_ hold161/X _4399_/X _4509_/S vssd1 vssd1 vccd1 vccd1 _4505_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_6_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4436_ hold198/X _4148_/X _4437_/S vssd1 vssd1 vccd1 vccd1 _6142_/D sky130_fd_sc_hd__mux2_1
X_4367_ _4382_/C _4364_/X _4365_/X _4366_/Y vssd1 vssd1 vccd1 vccd1 _4367_/X sky130_fd_sc_hd__a22o_2
X_3318_ _3349_/A _3318_/B _3318_/C _3318_/D vssd1 vssd1 vccd1 vccd1 _3318_/X sky130_fd_sc_hd__and4b_1
XFILLER_0_67_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6106_ _6444_/CLK _6106_/D vssd1 vssd1 vccd1 vccd1 _6106_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4892__A1 _6325_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4298_ _6078_/Q _4298_/B _6080_/Q vssd1 vssd1 vccd1 vccd1 _4299_/C sky130_fd_sc_hd__and3_1
XANTENNA__4644__A1 _6341_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3249_ _5313_/A _3686_/A vssd1 vssd1 vccd1 vccd1 _3249_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__5841__A0 _6326_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6037_ _3046_/A _6035_/X _6036_/Y hold387/X _6029_/Y vssd1 vssd1 vccd1 vccd1 _6037_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_0_83_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6440__SET_B fanout171/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold590 _6326_/Q vssd1 vssd1 vccd1 vccd1 hold590/X sky130_fd_sc_hd__buf_1
XANTENNA__4883__A1 _6325_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5596__C1 _5603_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5363__A2 _4639_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5270_ _5270_/A _5270_/B _5270_/C vssd1 vssd1 vccd1 vccd1 _5273_/C sky130_fd_sc_hd__or3_1
XFILLER_0_2_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3126__A1 _3183_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4221_ _4637_/A _4260_/A vssd1 vssd1 vccd1 vccd1 _4221_/X sky130_fd_sc_hd__or2_2
XANTENNA__3903__S _6243_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5390__S _5560_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4874__A1 _6324_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4152_ hold134/X _3779_/X _3781_/X _6106_/Q _4151_/X vssd1 vssd1 vccd1 vccd1 _4155_/A
+ sky130_fd_sc_hd__a221o_1
X_3103_ _3293_/B _3534_/A vssd1 vssd1 vccd1 vccd1 _3502_/A sky130_fd_sc_hd__or2_4
X_4083_ _4081_/S _3746_/X _3985_/A _5211_/D _4082_/X vssd1 vssd1 vccd1 vccd1 _4083_/X
+ sky130_fd_sc_hd__a221o_1
X_3034_ _3289_/A vssd1 vssd1 vccd1 vccd1 _3293_/B sky130_fd_sc_hd__inv_2
XANTENNA__5823__B1 _5932_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4985_ _5061_/A1 _4980_/X _4984_/X _4867_/B vssd1 vssd1 vccd1 vccd1 _4985_/X sky130_fd_sc_hd__a22o_1
XANTENNA_fanout143_A _5226_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3936_ _3938_/A _6338_/Q vssd1 vssd1 vccd1 vccd1 _3939_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__3113__D_N _3183_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3867_ _4389_/A _5249_/C vssd1 vssd1 vccd1 vccd1 _3868_/B sky130_fd_sc_hd__or2_1
XFILLER_0_5_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5606_ _4070_/A _5587_/X _5589_/X _6267_/Q _5605_/X vssd1 vssd1 vccd1 vccd1 _5606_/X
+ sky130_fd_sc_hd__a221o_1
X_3798_ _4111_/A _3798_/B vssd1 vssd1 vccd1 vccd1 _3799_/A sky130_fd_sc_hd__xnor2_1
X_5537_ hold577/X _5377_/X _5536_/Y _5441_/A vssd1 vssd1 vccd1 vccd1 _5537_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_14_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5468_ hold590/X _5377_/X _5467_/Y _5377_/A vssd1 vssd1 vccd1 vccd1 _5468_/Y sky130_fd_sc_hd__o2bb2ai_1
X_5399_ _5399_/A _5399_/B vssd1 vssd1 vccd1 vccd1 _5400_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4419_ hold81/X hold136/X hold89/X hold159/X _5673_/C1 _3718_/Y vssd1 vssd1 vccd1
+ vccd1 _4419_/X sky130_fd_sc_hd__mux4_1
XANTENNA__4617__A1 _5371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout56_A _5977_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_24_wb_clk_i _6404_/CLK vssd1 vssd1 vccd1 vccd1 _6270_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_37_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5593__A2 _6313_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4599__B _4604_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6118__RESET_B fanout173/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4305__A0 _6271_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6058__B1 _6063_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4608__A1 _6402_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5281__A1 _3656_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6054__B _6054_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4770_ _4637_/B _3512_/Y _4769_/X vssd1 vssd1 vccd1 vccd1 _5060_/S sky130_fd_sc_hd__o21ai_4
XFILLER_0_55_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3721_ _6077_/Q _4382_/C _3719_/X vssd1 vssd1 vccd1 vccd1 _3721_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_0_28_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3652_ _4309_/A _3652_/B vssd1 vssd1 vccd1 vccd1 _6125_/D sky130_fd_sc_hd__or2_1
XFILLER_0_43_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6440_ _6440_/CLK _6440_/D fanout171/X vssd1 vssd1 vccd1 vccd1 _6440_/Q sky130_fd_sc_hd__dfstp_1
X_3583_ _3583_/A _3583_/B _3605_/B _3583_/D vssd1 vssd1 vccd1 vccd1 _3606_/A sky130_fd_sc_hd__or4_1
X_6371_ _6374_/CLK _6371_/D fanout170/X vssd1 vssd1 vccd1 vccd1 _6371_/Q sky130_fd_sc_hd__dfrtp_1
X_5322_ _5322_/A _5322_/B _5322_/C _5322_/D vssd1 vssd1 vccd1 vccd1 _5482_/A sky130_fd_sc_hd__or4_1
X_5253_ _5253_/A _5253_/B _5253_/C _4022_/Y vssd1 vssd1 vccd1 vccd1 _5253_/X sky130_fd_sc_hd__or4b_1
X_5184_ _5209_/A _4025_/B _5183_/X _6304_/Q vssd1 vssd1 vccd1 vccd1 _5184_/X sky130_fd_sc_hd__o22a_1
X_4204_ _5690_/S _4201_/X _4202_/X _4203_/X vssd1 vssd1 vccd1 vccd1 _4204_/X sky130_fd_sc_hd__o31a_1
X_4135_ _6247_/Q _5217_/A _4135_/S vssd1 vssd1 vccd1 vccd1 _5212_/A sky130_fd_sc_hd__mux2_1
X_4066_ _4066_/A _4066_/B vssd1 vssd1 vccd1 vccd1 _4067_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_64_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4464__S _4464_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3588__B _4679_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3822__A2 _3789_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5024__A1 _6384_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4968_ _6329_/Q _5928_/A2 _5928_/B1 _4967_/X vssd1 vssd1 vccd1 vccd1 _4968_/X sky130_fd_sc_hd__a22o_1
X_3919_ _3919_/A _3919_/B vssd1 vssd1 vccd1 vccd1 _5251_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_34_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4899_ _4898_/X _4897_/X _6085_/Q vssd1 vssd1 vccd1 vccd1 _4900_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_61_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6282__RESET_B fanout169/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5308__B _5313_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3754__D _6304_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3109__A _4255_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4838__A1 _6322_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout130 _4309_/A vssd1 vssd1 vccd1 vccd1 _3337_/A sky130_fd_sc_hd__clkbuf_4
Xfanout141 hold671/X vssd1 vssd1 vccd1 vccd1 _3952_/A sky130_fd_sc_hd__clkbuf_4
Xfanout152 _3566_/A vssd1 vssd1 vccd1 vccd1 _4744_/B sky130_fd_sc_hd__buf_2
Xfanout174 fanout181/X vssd1 vssd1 vccd1 vccd1 fanout174/X sky130_fd_sc_hd__buf_6
Xfanout163 _4326_/B vssd1 vssd1 vccd1 vccd1 _5052_/S1 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_88_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6055__A3 _6054_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4882__B _4882_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3813__A2 _3784_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3329__A1 _6293_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5933__S _5933_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4829__A1 _6322_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5940_ _3081_/Y _5936_/B _5937_/B _5935_/A vssd1 vssd1 vccd1 vccd1 _5941_/B sky130_fd_sc_hd__o31a_1
XANTENNA__3265__B1 _3654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5254__B2 _5221_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5871_ hold558/X _5928_/A2 _5928_/B1 _5870_/X vssd1 vssd1 vccd1 vccd1 _5871_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_34_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4822_ hold338/X _4821_/Y _5068_/S vssd1 vssd1 vccd1 vccd1 _4822_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_90_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3568__A1 _6293_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4753_ _6389_/Q _6400_/Q _6223_/Q vssd1 vssd1 vccd1 vccd1 _5784_/S sky130_fd_sc_hd__nand3_2
XFILLER_0_62_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3704_ _6317_/Q hold1/A _3704_/S vssd1 vssd1 vccd1 vccd1 _3704_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4313__A _6064_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4860__S0 _5051_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6423_ _6423_/CLK _6423_/D fanout175/X vssd1 vssd1 vccd1 vccd1 _6423_/Q sky130_fd_sc_hd__dfrtp_4
X_4684_ _5226_/A _5553_/S _5226_/C vssd1 vssd1 vccd1 vccd1 _5102_/A sky130_fd_sc_hd__and3_2
XFILLER_0_70_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3635_ _3631_/Y _3634_/Y hold422/X vssd1 vssd1 vccd1 vccd1 _3635_/X sky130_fd_sc_hd__o21a_1
XANTENNA__5843__S _5932_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3566_ _3566_/A _3566_/B _5158_/B vssd1 vssd1 vccd1 vccd1 _5320_/B sky130_fd_sc_hd__or3_1
XANTENNA_fanout106_A _5472_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6354_ _6354_/CLK hold20/X vssd1 vssd1 vccd1 vccd1 hold19/A sky130_fd_sc_hd__dfxtp_1
X_5305_ _5313_/A _5296_/X _5304_/X _3530_/D _5301_/X vssd1 vssd1 vccd1 vccd1 _5305_/X
+ sky130_fd_sc_hd__a221o_1
X_3497_ _4070_/A _3100_/B _3277_/A _3496_/Y vssd1 vssd1 vccd1 vccd1 _3497_/X sky130_fd_sc_hd__a31o_1
XANTENNA__4459__S _4464_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6285_ _6376_/CLK _6285_/D fanout166/X vssd1 vssd1 vccd1 vccd1 _6285_/Q sky130_fd_sc_hd__dfrtp_2
X_5236_ _6298_/Q _5212_/B _5236_/S vssd1 vssd1 vccd1 vccd1 _5236_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_52_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5493__A1 _6057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5167_ hold357/X _5158_/A _5158_/B _5243_/S _5166_/X vssd1 vssd1 vccd1 vccd1 _5167_/X
+ sky130_fd_sc_hd__o311a_1
X_4118_ _4130_/A _4118_/B vssd1 vssd1 vccd1 vccd1 _4119_/B sky130_fd_sc_hd__nand2_1
X_5098_ _5098_/A _5242_/S _5178_/A vssd1 vssd1 vccd1 vccd1 _5098_/Y sky130_fd_sc_hd__nor3_1
XANTENNA__5245__A1 _3473_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4049_ _6048_/A vssd1 vssd1 vccd1 vccd1 _4049_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_78_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3731__A1 _6242_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3781__B _3850_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5054__A _5054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold8 hold8/A vssd1 vssd1 vccd1 vccd1 hold8/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5229__A _6417_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4842__S0 _5051_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold408 _4296_/X vssd1 vssd1 vccd1 vccd1 _6080_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3420_ _3654_/A _4347_/C _3391_/Y _5270_/A _3419_/X vssd1 vssd1 vccd1 vccd1 _3420_/X
+ sky130_fd_sc_hd__a221o_1
Xhold419 _3626_/X vssd1 vssd1 vccd1 vccd1 _6415_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3351_ _5096_/A _4541_/B vssd1 vssd1 vccd1 vccd1 _4346_/B sky130_fd_sc_hd__nand2_4
XFILLER_0_0_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3282_ _5303_/B _3573_/A _4214_/B vssd1 vssd1 vccd1 vccd1 _5323_/C sky130_fd_sc_hd__and3b_2
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6070_ _6194_/CLK _6070_/D vssd1 vssd1 vccd1 vccd1 _6070_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5021_ _6332_/Q _5039_/C vssd1 vssd1 vccd1 vccd1 _5021_/X sky130_fd_sc_hd__xor2_1
XANTENNA__5227__A1 _5240_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5923_ _5914_/A _5742_/A _5922_/X _5731_/X vssd1 vssd1 vccd1 vccd1 _5923_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_61_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5854_ _5848_/Y _5853_/X _5932_/S vssd1 vssd1 vccd1 vccd1 _5854_/X sky130_fd_sc_hd__mux2_1
X_4805_ hold39/A hold55/A hold45/A hold73/A _5358_/A0 _4326_/B vssd1 vssd1 vccd1 vccd1
+ _4805_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_8_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4202__A2 _4198_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5785_ _6322_/Q _5772_/S _5850_/B1 _5784_/X vssd1 vssd1 vccd1 vccd1 _5785_/X sky130_fd_sc_hd__a22o_1
X_4736_ _3511_/D _3773_/B _4734_/X _4735_/X vssd1 vssd1 vccd1 vccd1 _4736_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_71_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4667_ _5715_/B _4663_/Y _4666_/X hold355/X _4635_/Y vssd1 vssd1 vccd1 vccd1 _4667_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_0_31_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6406_ _6406_/CLK _6406_/D fanout180/X vssd1 vssd1 vccd1 vccd1 _6406_/Q sky130_fd_sc_hd__dfrtp_1
X_3618_ _4214_/A _3686_/A hold357/X _3426_/A _4750_/B vssd1 vssd1 vccd1 vccd1 _3619_/B
+ sky130_fd_sc_hd__a41o_1
XFILLER_0_43_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4598_ _5695_/A1 hold500/X _4546_/Y _4597_/X vssd1 vssd1 vccd1 vccd1 _4598_/X sky130_fd_sc_hd__a22o_1
X_6337_ _6343_/CLK _6337_/D vssd1 vssd1 vccd1 vccd1 _6337_/Q sky130_fd_sc_hd__dfxtp_2
X_3549_ _3549_/A _3549_/B vssd1 vssd1 vccd1 vccd1 _5324_/C sky130_fd_sc_hd__nor2_1
X_6268_ _6271_/CLK _6268_/D fanout170/X vssd1 vssd1 vccd1 vccd1 _6268_/Q sky130_fd_sc_hd__dfstp_4
X_5219_ _5219_/A _5219_/B _5219_/C _5219_/D vssd1 vssd1 vccd1 vccd1 _5219_/X sky130_fd_sc_hd__or4_1
XANTENNA__3477__B1 _5339_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6199_ _6354_/CLK _6199_/D vssd1 vssd1 vccd1 vccd1 _6199_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5602__A _5603_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4824__S0 _5358_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4901__A0 _6378_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3032__A _5935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3235__A3 _3566_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5090__C1 _6304_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5570_ _5599_/A _5603_/B _5603_/C _5339_/A vssd1 vssd1 vccd1 vccd1 _5571_/A sky130_fd_sc_hd__a31o_1
XFILLER_0_80_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4521_ _5447_/S _5371_/A _5075_/B vssd1 vssd1 vccd1 vccd1 _4539_/S sky130_fd_sc_hd__and3_4
XFILLER_0_13_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold216 _6093_/Q vssd1 vssd1 vccd1 vccd1 hold216/X sky130_fd_sc_hd__dlygate4sd3_1
X_4452_ _4054_/X hold235/X _4455_/S vssd1 vssd1 vccd1 vccd1 _6156_/D sky130_fd_sc_hd__mux2_1
Xhold205 _6069_/Q vssd1 vssd1 vccd1 vccd1 hold205/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold249 _6087_/Q vssd1 vssd1 vccd1 vccd1 hold249/X sky130_fd_sc_hd__dlygate4sd3_1
X_3403_ _3572_/A _3403_/B vssd1 vssd1 vccd1 vccd1 _5264_/B sky130_fd_sc_hd__or2_1
Xhold238 _6193_/Q vssd1 vssd1 vccd1 vccd1 hold238/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold227 _4434_/X vssd1 vssd1 vccd1 vccd1 _6140_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5406__B _6419_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4383_ hold55/A _4384_/S _5673_/C1 _4382_/X vssd1 vssd1 vccd1 vccd1 _4383_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_0_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6122_ _6122_/CLK _6126_/D fanout180/X vssd1 vssd1 vccd1 vccd1 _6122_/Q sky130_fd_sc_hd__dfstp_1
X_3334_ _4284_/A _5226_/A _3334_/C vssd1 vssd1 vccd1 vccd1 _5328_/C sky130_fd_sc_hd__and3_2
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3265_ _3611_/A _4346_/A _3654_/A _5097_/B _3546_/B vssd1 vssd1 vccd1 vccd1 _3265_/X
+ sky130_fd_sc_hd__o221a_1
X_6053_ _3046_/A _6051_/X _6052_/Y hold508/X _6029_/Y vssd1 vssd1 vccd1 vccd1 _6053_/X
+ sky130_fd_sc_hd__o32a_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5004_ _6420_/Q _5060_/S _5003_/Y vssd1 vssd1 vccd1 vccd1 _5004_/X sky130_fd_sc_hd__o21a_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5141__B _6247_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3196_ _3196_/A _3196_/B _3510_/B _5291_/A vssd1 vssd1 vccd1 vccd1 _3197_/C sky130_fd_sc_hd__or4_1
XANTENNA_fanout173_A fanout174/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4959__B1 _4958_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5906_ _5906_/A vssd1 vssd1 vccd1 vccd1 _5907_/B sky130_fd_sc_hd__inv_2
XANTENNA__4472__S _4473_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4806__S0 _5358_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5837_ _5846_/B _5837_/B vssd1 vssd1 vccd1 vccd1 _5837_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_36_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4187__A1 _6343_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5768_ _5769_/A _5769_/B _5767_/X vssd1 vssd1 vccd1 vccd1 _5782_/B sky130_fd_sc_hd__o21ba_1
XFILLER_0_71_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4719_ _4087_/Y _4718_/X _4731_/S vssd1 vssd1 vccd1 vccd1 _4719_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5136__B1 _5077_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5699_ _5699_/A vssd1 vssd1 vccd1 vccd1 _6345_/D sky130_fd_sc_hd__inv_2
XFILLER_0_4_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_49_wb_clk_i clkbuf_leaf_6_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6194_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__3117__A _3254_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3698__B1 _3365_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5611__A1 _6268_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5375__A0 _6416_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5226__B _6427_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3050_ _6305_/Q vssd1 vssd1 vccd1 vccd1 _5247_/A sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_10_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__6057__B _6057_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4102__B2 _4427_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3952_ _3952_/A _3952_/B vssd1 vssd1 vccd1 vccd1 _3953_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_73_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3883_ _5088_/B _6337_/Q vssd1 vssd1 vccd1 vccd1 _3886_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_73_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5622_ _6418_/Q _5602_/X _5603_/X _6373_/Q vssd1 vssd1 vccd1 vccd1 _5622_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_5_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5553_ _6448_/Q _5054_/B _5553_/S vssd1 vssd1 vccd1 vccd1 _5554_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_26_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5118__A0 _6293_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4504_ hold73/X _4392_/X _4509_/S vssd1 vssd1 vccd1 vccd1 hold74/A sky130_fd_sc_hd__mux2_1
XFILLER_0_41_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5484_ _5553_/S _5484_/B vssd1 vssd1 vccd1 vccd1 _5558_/S sky130_fd_sc_hd__nand2_4
XANTENNA__5669__A1 _6272_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4435_ hold282/X _4102_/X _4437_/S vssd1 vssd1 vccd1 vccd1 _6141_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_13_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4366_ _3079_/Y _3700_/B _4382_/C vssd1 vssd1 vccd1 vccd1 _4366_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_6_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3317_ _3186_/B _3316_/X _3369_/B vssd1 vssd1 vccd1 vccd1 _3318_/B sky130_fd_sc_hd__a21o_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6105_ _6194_/CLK hold80/X vssd1 vssd1 vccd1 vccd1 hold79/A sky130_fd_sc_hd__dfxtp_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4467__S _4473_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4297_ _6078_/Q _6079_/Q _6080_/Q _4287_/B _4299_/A vssd1 vssd1 vccd1 vccd1 _4297_/X
+ sky130_fd_sc_hd__a41o_1
X_3248_ _6392_/Q _3362_/B _3247_/X _5313_/A vssd1 vssd1 vccd1 vccd1 _3304_/A sky130_fd_sc_hd__a22oi_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6036_ _6036_/A _6063_/S vssd1 vssd1 vccd1 vccd1 _6036_/Y sky130_fd_sc_hd__nor2_1
X_3179_ _3220_/A _3243_/B vssd1 vssd1 vccd1 vccd1 _3277_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_83_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4801__C1 _5740_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4580__A1 _6418_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4580__B2 _6269_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold580 _5392_/X vssd1 vssd1 vccd1 vccd1 _6320_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold591 _5472_/X vssd1 vssd1 vccd1 vccd1 _6326_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4883__A2 _4752_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4399__A1 _4427_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4571__B2 _6267_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4571__A1 _6416_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4220_ _5317_/A _4220_/B vssd1 vssd1 vccd1 vccd1 _4260_/B sky130_fd_sc_hd__or2_1
X_4151_ _6222_/Q _3784_/X _3786_/X _6159_/Q vssd1 vssd1 vccd1 vccd1 _4151_/X sky130_fd_sc_hd__a22o_1
X_3102_ _3293_/B _3534_/A vssd1 vssd1 vccd1 vccd1 _3642_/C sky130_fd_sc_hd__nor2_1
X_4082_ _3746_/X _4081_/X _6341_/Q vssd1 vssd1 vccd1 vccd1 _4082_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_37_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4626__A2 _4615_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3033_ _3183_/B vssd1 vssd1 vccd1 vccd1 _3136_/B sky130_fd_sc_hd__inv_2
XANTENNA__3204__B _4679_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4984_ _6419_/Q _4983_/Y _5060_/S vssd1 vssd1 vccd1 vccd1 _4984_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4316__A _6064_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3935_ _3935_/A _3935_/B vssd1 vssd1 vccd1 vccd1 _5252_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_6_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5605_ _5594_/Y _5596_/X _5598_/X _5588_/X _6433_/Q vssd1 vssd1 vccd1 vccd1 _5605_/X
+ sky130_fd_sc_hd__a32o_1
X_3866_ _4394_/A _3866_/B vssd1 vssd1 vccd1 vccd1 _5249_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__6000__A1 _6057_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3797_ _3797_/A _3797_/B vssd1 vssd1 vccd1 vccd1 _3798_/B sky130_fd_sc_hd__nand2_2
X_5536_ _5536_/A vssd1 vssd1 vccd1 vccd1 _5536_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_14_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5467_ _5467_/A _5467_/B vssd1 vssd1 vccd1 vccd1 _5467_/Y sky130_fd_sc_hd__xnor2_1
X_4418_ hold3/X _4425_/A2 _5597_/B vssd1 vssd1 vccd1 vccd1 _4418_/X sky130_fd_sc_hd__o21a_1
X_5398_ _5367_/Y _5385_/B _5383_/X vssd1 vssd1 vccd1 vccd1 _5399_/B sky130_fd_sc_hd__a21o_1
X_4349_ _5560_/A _5327_/A _4349_/C _4748_/C vssd1 vssd1 vccd1 vccd1 _4349_/X sky130_fd_sc_hd__or4b_1
X_6019_ _3046_/A _6017_/X _6018_/Y hold540/X _5995_/Y vssd1 vssd1 vccd1 vccd1 _6019_/X
+ sky130_fd_sc_hd__o32a_1
XANTENNA__5290__A2 _5578_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3784__B _3850_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6294__SET_B fanout177/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5281__A2 _6118_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3816__B1 _3794_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3720_ _6077_/Q _4382_/C _3719_/X vssd1 vssd1 vccd1 vccd1 _3720_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_7_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3651_ _5715_/A _5975_/S _4541_/B vssd1 vssd1 vccd1 vccd1 _6241_/D sky130_fd_sc_hd__a21o_2
X_3582_ _3580_/Y _5315_/A _4767_/A vssd1 vssd1 vccd1 vccd1 _3583_/D sky130_fd_sc_hd__o21a_1
X_6370_ _6428_/CLK hold22/X vssd1 vssd1 vccd1 vccd1 hold21/A sky130_fd_sc_hd__dfxtp_1
X_5321_ hold128/X _5320_/Y _5321_/S vssd1 vssd1 vccd1 vccd1 _5321_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_51_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5252_ _5252_/A _5252_/B _4424_/B vssd1 vssd1 vccd1 vccd1 _5253_/C sky130_fd_sc_hd__or3b_1
X_5183_ _5087_/A _5087_/B _5182_/A _5182_/Y _3759_/B vssd1 vssd1 vccd1 vccd1 _5183_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4203_ _6314_/Q _5597_/B _5675_/C1 _4200_/X _4199_/X vssd1 vssd1 vccd1 vccd1 _4203_/X
+ sky130_fd_sc_hd__a221o_1
X_4134_ _4255_/B _4134_/B vssd1 vssd1 vccd1 vccd1 _4134_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__5257__C1 _5258_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4065_ _5087_/A _6247_/Q _6341_/Q _3740_/Y _4064_/X vssd1 vssd1 vccd1 vccd1 _5206_/B
+ sky130_fd_sc_hd__o41a_2
XANTENNA__3807__B1 _3781_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3283__A1 _3254_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4232__B1 _5315_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4480__S _4482_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4967_ _6362_/Q _4966_/X _5927_/S vssd1 vssd1 vccd1 vccd1 _4967_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3918_ _4394_/A _3798_/B _3876_/X vssd1 vssd1 vccd1 vccd1 _3919_/B sky130_fd_sc_hd__o21ai_1
X_4898_ _6167_/Q _6175_/Q _6414_/Q _6183_/Q _6318_/Q _6090_/Q vssd1 vssd1 vccd1 vccd1
+ _4898_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_61_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3849_ hold115/X hold239/X _3861_/S vssd1 vssd1 vccd1 vccd1 _3850_/C sky130_fd_sc_hd__mux2_1
XFILLER_0_27_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5732__B1 _4214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4535__A1 _6294_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5519_ _5554_/A _5520_/B vssd1 vssd1 vccd1 vccd1 _5519_/X sky130_fd_sc_hd__and2_1
XANTENNA__6251__RESET_B fanout179/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout131 hold666/X vssd1 vssd1 vccd1 vccd1 _4309_/A sky130_fd_sc_hd__buf_4
Xfanout120 _6402_/Q vssd1 vssd1 vccd1 vccd1 _5695_/A1 sky130_fd_sc_hd__buf_4
Xfanout153 hold674/X vssd1 vssd1 vccd1 vccd1 _3566_/A sky130_fd_sc_hd__clkbuf_4
Xfanout142 _3482_/A vssd1 vssd1 vccd1 vccd1 _4228_/A sky130_fd_sc_hd__buf_4
Xfanout164 hold656/X vssd1 vssd1 vccd1 vccd1 _4326_/B sky130_fd_sc_hd__buf_6
Xfanout175 fanout178/X vssd1 vssd1 vccd1 vccd1 fanout175/X sky130_fd_sc_hd__clkbuf_8
XANTENNA_hold632_A _6417_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3779__B _3850_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5971__A0 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5723__A0 _6274_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4526__A1 _6269_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3035__A _4284_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4565__S _4604_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3265__A1 _3611_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3265__B2 _5097_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5870_ _6362_/Q _6381_/Q _5927_/S vssd1 vssd1 vccd1 vccd1 _5870_/X sky130_fd_sc_hd__mux2_1
X_4821_ _3073_/Y _5557_/S _4820_/X vssd1 vssd1 vccd1 vccd1 _4821_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4752_ _6389_/Q _6400_/Q _6223_/Q vssd1 vssd1 vccd1 vccd1 _4752_/X sky130_fd_sc_hd__and3_2
XFILLER_0_50_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5962__A0 _4392_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3703_ _3473_/A _3697_/X _3674_/B _3669_/X vssd1 vssd1 vccd1 vccd1 _3704_/S sky130_fd_sc_hd__o211ai_4
XFILLER_0_50_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4683_ _5740_/A _4682_/X _4681_/X _3072_/Y vssd1 vssd1 vccd1 vccd1 _4683_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_43_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4860__S1 _5052_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3634_ _6405_/Q _3634_/B vssd1 vssd1 vccd1 vccd1 _3634_/Y sky130_fd_sc_hd__nor2_1
X_6422_ _6423_/CLK _6422_/D fanout175/X vssd1 vssd1 vccd1 vccd1 _6422_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_43_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3565_ _4637_/A _4745_/B vssd1 vssd1 vccd1 vccd1 _5158_/B sky130_fd_sc_hd__or2_2
XFILLER_0_59_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6353_ _6355_/CLK hold14/X vssd1 vssd1 vccd1 vccd1 hold13/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5304_ _3482_/A _5302_/X _5303_/Y _3426_/A vssd1 vssd1 vccd1 vccd1 _5304_/X sky130_fd_sc_hd__a211o_1
X_3496_ _3496_/A _3496_/B vssd1 vssd1 vccd1 vccd1 _3496_/Y sky130_fd_sc_hd__nor2_1
X_6284_ _6290_/CLK _6284_/D fanout166/X vssd1 vssd1 vccd1 vccd1 _6284_/Q sky130_fd_sc_hd__dfrtp_2
X_5235_ _6298_/Q _5109_/B _5347_/B vssd1 vssd1 vccd1 vccd1 _5235_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5493__A2 _5377_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5166_ _5154_/X _5157_/X _5165_/Y _5242_/S _5158_/Y vssd1 vssd1 vccd1 vccd1 _5166_/X
+ sky130_fd_sc_hd__a221o_1
X_4117_ _4130_/A _4118_/B vssd1 vssd1 vccd1 vccd1 _4122_/B sky130_fd_sc_hd__nor2_1
X_5097_ _5097_/A _5097_/B _5158_/B vssd1 vssd1 vccd1 vccd1 _5178_/A sky130_fd_sc_hd__nor3_2
XANTENNA__5160__A _6417_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4475__S _4482_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4048_ _4029_/B _4047_/Y _4142_/S vssd1 vssd1 vccd1 vccd1 _6048_/A sky130_fd_sc_hd__mux2_4
XANTENNA__5650__C1 _5673_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5999_ _5339_/A _5997_/X _5998_/Y hold498/X _5995_/Y vssd1 vssd1 vccd1 vccd1 _5999_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_0_19_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6432__RESET_B fanout178/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3731__A2 _6336_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3781__C _3838_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3495__B2 _4070_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold9 hold9/A vssd1 vssd1 vccd1 vccd1 hold9/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5229__B _6416_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4842__S1 _5052_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold409 _6289_/Q vssd1 vssd1 vccd1 vccd1 hold409/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3350_ _4210_/A _5578_/A vssd1 vssd1 vccd1 vccd1 _4208_/B sky130_fd_sc_hd__nor2_2
XANTENNA__3400__C_N _5313_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3281_ _3281_/A _3281_/B vssd1 vssd1 vccd1 vccd1 _3281_/Y sky130_fd_sc_hd__nor2_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5020_ _5016_/B _5019_/X _5058_/S vssd1 vssd1 vccd1 vccd1 _5020_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_29_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4295__S _4305_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5922_ _5932_/S _5917_/Y _5921_/X _5747_/A vssd1 vssd1 vccd1 vccd1 _5922_/X sky130_fd_sc_hd__o22a_1
X_5853_ _5852_/X _5845_/A _5931_/S vssd1 vssd1 vccd1 vccd1 _5853_/X sky130_fd_sc_hd__mux2_1
X_5784_ _6322_/Q _5778_/A _5784_/S vssd1 vssd1 vccd1 vccd1 _5784_/X sky130_fd_sc_hd__mux2_1
X_4804_ _6321_/Q _4752_/X _4751_/B vssd1 vssd1 vccd1 vccd1 _4804_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_90_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4735_ _3367_/B _4745_/B _6389_/Q _5270_/C vssd1 vssd1 vccd1 vccd1 _4735_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_8_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5854__S _5932_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4666_ _3691_/B _4665_/X _4673_/B vssd1 vssd1 vccd1 vccd1 _4666_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_43_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3961__A2 _6040_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3617_ _4541_/A hold249/X hold118/X _6391_/Q _3616_/X vssd1 vssd1 vccd1 vccd1 _4750_/B
+ sky130_fd_sc_hd__a221o_2
X_6405_ _6423_/CLK _6405_/D fanout178/X vssd1 vssd1 vccd1 vccd1 _6405_/Q sky130_fd_sc_hd__dfrtp_4
X_4597_ _6438_/Q _4567_/Y _4568_/X _6446_/Q _4596_/X vssd1 vssd1 vccd1 vccd1 _4597_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_101_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3548_ _4639_/C _4767_/B _4224_/C _3546_/Y _3547_/Y vssd1 vssd1 vccd1 vccd1 _3548_/Y
+ sky130_fd_sc_hd__a221oi_2
X_6336_ _6373_/CLK _6336_/D vssd1 vssd1 vccd1 vccd1 _6336_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__4910__A1 _6378_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3479_ _4767_/A _3479_/B vssd1 vssd1 vccd1 vccd1 _3505_/A sky130_fd_sc_hd__and2_1
X_6267_ _6271_/CLK _6267_/D fanout170/X vssd1 vssd1 vccd1 vccd1 _6267_/Q sky130_fd_sc_hd__dfstp_2
XANTENNA__4674__A0 _6339_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5218_ _3761_/Y _5216_/X _5217_/X _5148_/X _5150_/Y vssd1 vssd1 vccd1 vccd1 _5218_/X
+ sky130_fd_sc_hd__o311a_1
XANTENNA__3477__A1 _5975_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6198_ _6221_/CLK _6198_/D vssd1 vssd1 vccd1 vccd1 _6198_/Q sky130_fd_sc_hd__dfxtp_1
X_5149_ _6304_/Q _5150_/B vssd1 vssd1 vccd1 vccd1 _5149_/X sky130_fd_sc_hd__and2_1
XANTENNA__4933__S _5557_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4977__A1 _6270_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4729__B2 _5371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4729__A1 _6274_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4824__S1 _4326_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3792__B _3850_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4901__A1 _6326_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3313__A _4228_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5614__C1 _5676_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4843__S _5053_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3967__B _6339_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6008__A2_N _6054_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4520_ _5077_/A _4520_/B vssd1 vssd1 vccd1 vccd1 _4520_/Y sky130_fd_sc_hd__nand2_2
XANTENNA__5145__B2 _6336_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5145__A1 _6341_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold217 _4331_/X vssd1 vssd1 vccd1 vccd1 _6093_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4451_ _4007_/X hold271/X _4455_/S vssd1 vssd1 vccd1 vccd1 _6155_/D sky130_fd_sc_hd__mux2_1
Xhold206 _3924_/X vssd1 vssd1 vccd1 vccd1 _6069_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3402_ _4679_/D _3594_/A _4222_/B vssd1 vssd1 vccd1 vccd1 _4284_/C sky130_fd_sc_hd__and3b_2
Xhold239 _6408_/Q vssd1 vssd1 vccd1 vccd1 hold239/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold228 _6165_/Q vssd1 vssd1 vccd1 vccd1 hold228/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6121_ _6291_/CLK _6124_/D fanout176/X vssd1 vssd1 vccd1 vccd1 _6121_/Q sky130_fd_sc_hd__dfstp_1
X_4382_ hold39/A _4382_/B _4382_/C vssd1 vssd1 vccd1 vccd1 _4382_/X sky130_fd_sc_hd__or3_1
XFILLER_0_21_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3333_ _3896_/S _3332_/Y _3333_/S vssd1 vssd1 vccd1 vccd1 _3336_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_0_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3264_ _3611_/A _3501_/B _3654_/A _5265_/B _3632_/B vssd1 vssd1 vccd1 vccd1 _3264_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_56_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6052_ _6052_/A _6063_/S vssd1 vssd1 vccd1 vccd1 _6052_/Y sky130_fd_sc_hd__nor2_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5003_ _5039_/C _5002_/Y _5060_/S vssd1 vssd1 vccd1 vccd1 _5003_/Y sky130_fd_sc_hd__o21ai_1
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3195_ _3549_/A _3195_/B vssd1 vssd1 vccd1 vccd1 _5291_/A sky130_fd_sc_hd__nor2_2
XANTENNA__3223__A _3278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4959__A1 _6269_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5905_ _5905_/A _5926_/A vssd1 vssd1 vccd1 vccd1 _5906_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_36_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4806__S1 _4326_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5836_ _5836_/A _5836_/B _5834_/X vssd1 vssd1 vccd1 vccd1 _5837_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_63_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5767_ _5782_/A _5767_/B vssd1 vssd1 vccd1 vccd1 _5767_/X sky130_fd_sc_hd__or2_1
X_4718_ _4716_/X _4717_/X _5102_/A vssd1 vssd1 vccd1 vccd1 _4718_/X sky130_fd_sc_hd__mux2_1
X_5698_ _3080_/Y _4574_/A _5727_/S vssd1 vssd1 vccd1 vccd1 _5698_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_16_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4649_ _4648_/X _6342_/Q _4675_/S vssd1 vssd1 vccd1 vccd1 _4649_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5687__A2 _6313_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3084__1 _6406_/CLK vssd1 vssd1 vccd1 vccd1 _6122_/CLK sky130_fd_sc_hd__inv_2
XANTENNA__3698__A1 _3473_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3117__B _3183_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6319_ _6326_/CLK _6319_/D fanout175/X vssd1 vssd1 vccd1 vccd1 _6319_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_12_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_18_wb_clk_i _6404_/CLK vssd1 vssd1 vccd1 vccd1 _6403_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA_fanout79_A _4321_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3787__B _3862_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3925__A2 _3784_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5127__A1 _6292_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3308__A _3611_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4638__A0 _6242_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3310__B1 _5096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6057__C _6057_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_6_wb_clk_i_A clkbuf_leaf_6_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_3951_ _3761_/A _5216_/C _5211_/A _3985_/A _4040_/A vssd1 vssd1 vccd1 vccd1 _3951_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_58_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3882_ _3881_/X hold298/X _4206_/S vssd1 vssd1 vccd1 vccd1 _3882_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4169__A2 _5217_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5621_ _5695_/A1 _3907_/A _5571_/Y _5620_/X vssd1 vssd1 vccd1 vccd1 _5621_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5366__A1 _5715_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5552_ _5544_/B _5546_/B _5542_/X vssd1 vssd1 vccd1 vccd1 _5555_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_26_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4503_ hold57/X _4380_/X _4509_/S vssd1 vssd1 vccd1 vccd1 hold58/A sky130_fd_sc_hd__mux2_1
XFILLER_0_26_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5483_ _5480_/D _3512_/Y _4748_/X _5482_/Y vssd1 vssd1 vccd1 vccd1 _5484_/B sky130_fd_sc_hd__a2bb2o_2
XANTENNA__4321__B _4321_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4434_ hold226/X _4054_/X _4437_/S vssd1 vssd1 vccd1 vccd1 _4434_/X sky130_fd_sc_hd__mux2_1
X_4365_ _3724_/A _5249_/B _3768_/Y vssd1 vssd1 vccd1 vccd1 _4365_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_6_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3316_ _4679_/C _3309_/Y _3315_/Y _3590_/B vssd1 vssd1 vccd1 vccd1 _3316_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_67_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6104_ _6444_/CLK _6104_/D vssd1 vssd1 vccd1 vccd1 _6104_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6035_ _4313_/C _6034_/X _6063_/S vssd1 vssd1 vccd1 vccd1 _6035_/X sky130_fd_sc_hd__o21a_1
X_4296_ _3073_/A _4295_/X _4296_/S vssd1 vssd1 vccd1 vccd1 _4296_/X sky130_fd_sc_hd__mux2_1
X_3247_ _3247_/A _3247_/B _3247_/C vssd1 vssd1 vccd1 vccd1 _3247_/X sky130_fd_sc_hd__or3_1
XANTENNA__4049__A _6048_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3178_ _4522_/B _5303_/A _4522_/D vssd1 vssd1 vccd1 vccd1 _4520_/B sky130_fd_sc_hd__nor3_4
XFILLER_0_95_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3478__B1_N _3477_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6276__RESET_B fanout169/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6205__RESET_B fanout174/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3604__A1 _4637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3400__B _3400_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5819_ _6377_/Q _5819_/B vssd1 vssd1 vccd1 vccd1 _5820_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_44_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3128__A _4685_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4350__A2_N _5317_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold581 _6312_/Q vssd1 vssd1 vccd1 vccd1 _3066_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold570 _6431_/Q vssd1 vssd1 vccd1 vccd1 _3630_/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_hold662_A _6270_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold592 _6324_/Q vssd1 vssd1 vccd1 vccd1 hold592/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4393__S _4428_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5596__A1 _5690_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5348__A1 _5077_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4150_ _4115_/A _4115_/B _4112_/A vssd1 vssd1 vccd1 vccd1 _4157_/A sky130_fd_sc_hd__a21o_1
X_3101_ _3183_/B _3254_/A vssd1 vssd1 vccd1 vccd1 _3534_/A sky130_fd_sc_hd__nand2b_4
X_4081_ _3748_/Y _4188_/C _4081_/S vssd1 vssd1 vccd1 vccd1 _4081_/X sky130_fd_sc_hd__mux2_1
X_3032_ _5935_/A vssd1 vssd1 vccd1 vccd1 _5952_/A sky130_fd_sc_hd__clkinv_4
XFILLER_0_78_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3501__A _4637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3220__B _3566_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4983_ _5002_/B _4983_/B vssd1 vssd1 vccd1 vccd1 _4983_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__4316__B _4316_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3934_ _4009_/A _3934_/B _3934_/C vssd1 vssd1 vccd1 vccd1 _3935_/B sky130_fd_sc_hd__and3_1
XFILLER_0_73_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3865_ _3853_/Y _3864_/A _3864_/B _3855_/A vssd1 vssd1 vccd1 vccd1 _4389_/A sky130_fd_sc_hd__o31a_1
XFILLER_0_6_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3647__S input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5604_ _6441_/Q _5610_/B _5602_/C vssd1 vssd1 vccd1 vccd1 _5604_/X sky130_fd_sc_hd__a21o_1
XANTENNA__6000__A2 _4788_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout129_A _3337_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3796_ hold298/X _4474_/A _4501_/A hold278/X _3793_/X vssd1 vssd1 vccd1 vccd1 _3797_/B
+ sky130_fd_sc_hd__o221a_1
X_5535_ _5535_/A _5535_/B vssd1 vssd1 vccd1 vccd1 _5536_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5466_ _5464_/Y _5466_/B vssd1 vssd1 vccd1 vccd1 _5467_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__4478__S _4482_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4417_ _3724_/A _5251_/B _4144_/X vssd1 vssd1 vccd1 vccd1 _4417_/X sky130_fd_sc_hd__a21bo_1
X_5397_ _5395_/X _5397_/B vssd1 vssd1 vccd1 vccd1 _5399_/A sky130_fd_sc_hd__and2b_1
X_4348_ _4348_/A _5326_/C vssd1 vssd1 vccd1 vccd1 _4748_/C sky130_fd_sc_hd__nor2_1
X_4279_ _4279_/A _5603_/B vssd1 vssd1 vccd1 vccd1 _5349_/B sky130_fd_sc_hd__nand2_1
X_6018_ _6052_/A _6026_/B vssd1 vssd1 vccd1 vccd1 _6018_/Y sky130_fd_sc_hd__nor2_1
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4250__A1 _4214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3130__B _3952_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4941__S _6315_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4250__B2 _3337_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4242__A _4568_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5772__S _5772_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_33_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6271_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_20_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4936__S0 _5051_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6058__A2 _5557_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3650_ _6126_/Q _6122_/Q input1/X vssd1 vssd1 vccd1 vccd1 _3650_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_82_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3581_ _3581_/A _3581_/B vssd1 vssd1 vccd1 vccd1 _5315_/A sky130_fd_sc_hd__nor2_4
XFILLER_0_70_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5741__A1 _5931_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5320_ _6399_/Q _5320_/B vssd1 vssd1 vccd1 vccd1 _5320_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5251_ _5251_/A _5251_/B _5251_/C _4409_/B vssd1 vssd1 vccd1 vccd1 _5252_/A sky130_fd_sc_hd__or4b_1
X_4202_ hold286/X _4198_/B _4200_/S hold201/X _5675_/C1 vssd1 vssd1 vccd1 vccd1 _4202_/X
+ sky130_fd_sc_hd__o221a_1
X_5182_ _5182_/A _5182_/B vssd1 vssd1 vccd1 vccd1 _5182_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__3215__B _4224_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4133_ _6292_/Q _4132_/Y _4129_/X vssd1 vssd1 vccd1 vccd1 _5120_/A sky130_fd_sc_hd__a21oi_2
X_4064_ _3740_/Y _4060_/X _4061_/X _4063_/X vssd1 vssd1 vccd1 vccd1 _4064_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3283__A2 _3573_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4761__S _6315_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4232__A1 _3656_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4966_ _6381_/Q _4754_/X _4960_/X _4965_/X vssd1 vssd1 vccd1 vccd1 _4966_/X sky130_fd_sc_hd__a211o_1
XANTENNA__3991__A0 _6419_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5158__A _5158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3917_ _4394_/A _3917_/B vssd1 vssd1 vccd1 vccd1 _3919_/A sky130_fd_sc_hd__xnor2_2
X_4897_ hold71/A hold65/A _6135_/Q _6214_/Q _6318_/Q _6090_/Q vssd1 vssd1 vccd1 vccd1
+ _4897_/X sky130_fd_sc_hd__mux4_1
XANTENNA__4783__A2 _4752_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3848_ _3850_/A _3862_/S _3848_/C vssd1 vssd1 vccd1 vccd1 _3852_/C sky130_fd_sc_hd__or3_1
XFILLER_0_6_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3779_ _3850_/A _3850_/B _3861_/S vssd1 vssd1 vccd1 vccd1 _3779_/X sky130_fd_sc_hd__and3_4
XANTENNA__4569__A_N _4604_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5518_ _6445_/Q _4996_/B _5518_/S vssd1 vssd1 vccd1 vccd1 _5520_/B sky130_fd_sc_hd__mux2_1
XANTENNA__4918__S0 _5052_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5449_ _6439_/Q _4882_/B _5553_/S vssd1 vssd1 vccd1 vccd1 _5450_/C sky130_fd_sc_hd__mux2_1
Xfanout121 _5560_/B vssd1 vssd1 vccd1 vccd1 _5715_/B sky130_fd_sc_hd__clkbuf_8
Xfanout110 _3046_/Y vssd1 vssd1 vccd1 vccd1 _4732_/S sky130_fd_sc_hd__clkbuf_8
Xfanout143 _5226_/A vssd1 vssd1 vccd1 vccd1 _3525_/B sky130_fd_sc_hd__buf_4
Xfanout154 hold659/X vssd1 vssd1 vccd1 vccd1 _3254_/A sky130_fd_sc_hd__buf_6
Xfanout165 hold630/X vssd1 vssd1 vccd1 vccd1 _5053_/S sky130_fd_sc_hd__buf_8
Xfanout132 _5358_/A0 vssd1 vssd1 vccd1 vccd1 _5051_/S0 sky130_fd_sc_hd__buf_6
XANTENNA__5248__B1 _5560_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout176 fanout177/X vssd1 vssd1 vccd1 vccd1 fanout176/X sky130_fd_sc_hd__clkbuf_8
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3795__B _3850_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5723__A1 hold560/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6379__RESET_B fanout168/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6308__RESET_B fanout173/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3051__A _6304_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4820_ _4809_/A _5728_/D _4818_/Y _4819_/Y _4313_/C vssd1 vssd1 vccd1 vccd1 _4820_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3422__C1 _5935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4751_ _5825_/S _4751_/B vssd1 vssd1 vccd1 vccd1 _4751_/Y sky130_fd_sc_hd__nor2_1
X_3702_ _3473_/A _3697_/X _3674_/B _3669_/X vssd1 vssd1 vccd1 vccd1 _3702_/X sky130_fd_sc_hd__o211a_1
X_4682_ _6225_/Q _4520_/Y _4680_/X _3072_/Y vssd1 vssd1 vccd1 vccd1 _4682_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_7_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3633_ _5715_/A _3633_/B _3629_/B vssd1 vssd1 vccd1 vccd1 _3641_/A sky130_fd_sc_hd__or3b_1
X_6421_ _6421_/CLK _6421_/D fanout175/X vssd1 vssd1 vccd1 vccd1 _6421_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__4313__C _4313_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3564_ _6487_/A vssd1 vssd1 vccd1 vccd1 _3583_/A sky130_fd_sc_hd__inv_2
XFILLER_0_51_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6352_ _6408_/CLK _6352_/D vssd1 vssd1 vccd1 vccd1 _6352_/Q sky130_fd_sc_hd__dfxtp_1
X_5303_ _5303_/A _5303_/B vssd1 vssd1 vccd1 vccd1 _5303_/Y sky130_fd_sc_hd__nor2_1
X_3495_ _3333_/S _5715_/C _3537_/A _4070_/A _3494_/X vssd1 vssd1 vccd1 vccd1 _3496_/B
+ sky130_fd_sc_hd__o221a_1
X_6283_ _6290_/CLK _6283_/D fanout166/X vssd1 vssd1 vccd1 vccd1 _6283_/Q sky130_fd_sc_hd__dfrtp_2
X_5234_ hold652/X _5233_/X _5447_/S vssd1 vssd1 vccd1 vccd1 _6297_/D sky130_fd_sc_hd__mux2_1
X_5165_ _5165_/A _5165_/B vssd1 vssd1 vccd1 vccd1 _5165_/Y sky130_fd_sc_hd__xnor2_1
X_4116_ _5088_/B _6342_/Q vssd1 vssd1 vccd1 vccd1 _4118_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5441__A _5441_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5096_ _5096_/A _5096_/B _5979_/A _5096_/D vssd1 vssd1 vccd1 vccd1 _5242_/S sky130_fd_sc_hd__and4_2
X_4047_ _5247_/A _6420_/Q _4046_/X vssd1 vssd1 vccd1 vccd1 _4047_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__5160__B _6416_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4491__S _4491_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5998_ _6032_/A _6026_/B vssd1 vssd1 vccd1 vccd1 _5998_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__4205__B2 _4427_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4949_ _6361_/Q _4948_/X _5927_/S vssd1 vssd1 vccd1 vccd1 _4949_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_61_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3835__S _3838_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4520__A _5077_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3136__A _3254_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6401__RESET_B fanout178/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3495__A2 _5715_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4692__A1 _6268_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4692__B2 _5029_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6446__SET_B fanout171/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5229__C _6421_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3707__B1 _4382_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5172__A2 _5075_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3280_ _3280_/A _3600_/C _3386_/B _3592_/A vssd1 vssd1 vccd1 vccd1 _3281_/B sky130_fd_sc_hd__or4_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5921_ _6422_/Q _5920_/X _5930_/S vssd1 vssd1 vccd1 vccd1 _5921_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_75_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5852_ _6416_/Q _5851_/X _5852_/S vssd1 vssd1 vccd1 vccd1 _5852_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_75_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4199__B1 _5673_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4803_ hold373/X _4802_/X _5068_/S vssd1 vssd1 vccd1 vccd1 _4803_/X sky130_fd_sc_hd__mux2_1
X_5783_ _5795_/B _5783_/B vssd1 vssd1 vccd1 vccd1 _5783_/X sky130_fd_sc_hd__and2b_1
XANTENNA__3946__A0 _6292_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4734_ _3337_/B _4734_/B _4734_/C vssd1 vssd1 vccd1 vccd1 _4734_/X sky130_fd_sc_hd__and3b_1
XFILLER_0_16_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4665_ _4664_/X _6243_/Q _4675_/S vssd1 vssd1 vccd1 vccd1 _4665_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_9_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6404_ _6404_/CLK _6404_/D fanout180/X vssd1 vssd1 vccd1 vccd1 _6404_/Q sky130_fd_sc_hd__dfrtp_1
X_3616_ _6390_/Q _6086_/Q _6089_/Q _6389_/Q _3615_/Y vssd1 vssd1 vccd1 vccd1 _3616_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout111_A _5236_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4596_ _6421_/Q _4569_/X _4570_/X _6272_/Q _4595_/X vssd1 vssd1 vccd1 vccd1 _4596_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3225__C_N _3254_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3547_ _4257_/B _5256_/A _4346_/B _5096_/B vssd1 vssd1 vccd1 vccd1 _3547_/Y sky130_fd_sc_hd__o31ai_1
X_6335_ _6433_/CLK _6335_/D fanout174/X vssd1 vssd1 vccd1 vccd1 _6335_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_0_12_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6266_ _6266_/CLK _6266_/D fanout177/X vssd1 vssd1 vccd1 vccd1 _6266_/Q sky130_fd_sc_hd__dfrtp_1
X_3478_ _4323_/A _5560_/D _3477_/X vssd1 vssd1 vccd1 vccd1 _3484_/B sky130_fd_sc_hd__o21bai_1
XANTENNA__4674__A1 _6343_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5217_ _5217_/A _6246_/Q _6247_/Q _6248_/Q vssd1 vssd1 vccd1 vccd1 _5217_/X sky130_fd_sc_hd__or4_1
XANTENNA__4486__S _4491_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3477__A2 _5560_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6197_ _6354_/CLK _6197_/D vssd1 vssd1 vccd1 vccd1 _6197_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5148_ _6340_/Q _4042_/A _5144_/X _5147_/X vssd1 vssd1 vccd1 vccd1 _5148_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_98_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5079_ _4070_/A _5193_/S _5078_/Y _5076_/A vssd1 vssd1 vccd1 vccd1 _5079_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_79_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3792__C _3838_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4362__B1 _5339_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4665__A1 _6243_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3468__A2 _6389_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5081__A _5977_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5862__A0 _6417_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3313__B _5578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5614__B1 _5676_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5020__S _5058_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3928__B1 _3794_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4160__A _5217_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6394__RESET_B fanout179/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4450_ _3965_/X hold183/X _4455_/S vssd1 vssd1 vccd1 vccd1 _4450_/X sky130_fd_sc_hd__mux2_1
Xhold207 _6091_/Q vssd1 vssd1 vccd1 vccd1 hold207/X sky130_fd_sc_hd__dlygate4sd3_1
X_3401_ _3401_/A vssd1 vssd1 vccd1 vccd1 _3434_/B sky130_fd_sc_hd__inv_2
XANTENNA__6323__RESET_B fanout173/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4381_ hold75/X _4380_/X _4428_/S vssd1 vssd1 vccd1 vccd1 hold76/A sky130_fd_sc_hd__mux2_1
Xhold229 _6139_/Q vssd1 vssd1 vccd1 vccd1 hold229/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold218 _6180_/Q vssd1 vssd1 vccd1 vccd1 hold218/X sky130_fd_sc_hd__dlygate4sd3_1
X_3332_ _3525_/A _3525_/B _3334_/C vssd1 vssd1 vccd1 vccd1 _3332_/Y sky130_fd_sc_hd__nor3_1
X_6120_ _6270_/CLK _6125_/D fanout176/X vssd1 vssd1 vccd1 vccd1 _6120_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA__5690__S _5690_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3263_ _5265_/B _3654_/A vssd1 vssd1 vccd1 vccd1 _3263_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__4105__B1 _3786_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6051_ _6057_/A _6050_/X _6063_/S vssd1 vssd1 vccd1 vccd1 _6051_/X sky130_fd_sc_hd__o21a_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3194_ _3194_/A _3194_/B vssd1 vssd1 vccd1 vccd1 _3195_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_56_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5002_ _6331_/Q _5002_/B vssd1 vssd1 vccd1 vccd1 _5002_/Y sky130_fd_sc_hd__nor2_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3223__B _3566_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5904_ _5905_/A _5926_/A vssd1 vssd1 vccd1 vccd1 _5907_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_48_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5835_ _5836_/A _5836_/B _5834_/X vssd1 vssd1 vccd1 vccd1 _5846_/B sky130_fd_sc_hd__o21ba_1
XFILLER_0_91_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6030__B1 _6057_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5766_ _6373_/Q _5766_/B vssd1 vssd1 vccd1 vccd1 _5767_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_71_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5697_ _5697_/A vssd1 vssd1 vccd1 vccd1 _6344_/D sky130_fd_sc_hd__inv_2
X_4717_ hold534/X _4313_/B _4727_/S vssd1 vssd1 vccd1 vccd1 _4717_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4070__A _4070_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4648_ _6244_/Q _6338_/Q _4674_/S vssd1 vssd1 vccd1 vccd1 _4648_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_71_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4579_ _3930_/B _3841_/Y _4604_/S vssd1 vssd1 vccd1 vccd1 _4579_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_97_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6318_ _6433_/CLK _6318_/D vssd1 vssd1 vccd1 vccd1 _6318_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__4647__A1 _5715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6249_ _6421_/CLK _6249_/D vssd1 vssd1 vccd1 vccd1 _6249_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_hold538_A _6378_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3308__B _5158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4886__A1 _6325_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4638__A1 _6336_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5015__S _5053_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold90 hold90/A vssd1 vssd1 vccd1 vccd1 hold90/X sky130_fd_sc_hd__dlygate4sd3_1
X_3950_ _6243_/Q _6245_/Q _4135_/S vssd1 vssd1 vccd1 vccd1 _5211_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_58_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3881_ _4427_/S _3722_/X _3879_/X _3880_/Y vssd1 vssd1 vccd1 vccd1 _3881_/X sky130_fd_sc_hd__a22o_2
XANTENNA__6012__B1 _6057_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3994__A _6044_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4169__A3 _6343_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5620_ _5620_/A _5620_/B vssd1 vssd1 vccd1 vccd1 _5620_/X sky130_fd_sc_hd__or2_1
XFILLER_0_38_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5551_ _5548_/A _5550_/X _6060_/S vssd1 vssd1 vccd1 vccd1 _5551_/X sky130_fd_sc_hd__mux2_1
X_4502_ hold124/X _4367_/X _4509_/S vssd1 vssd1 vccd1 vccd1 _4502_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_26_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5482_ _5482_/A _5482_/B vssd1 vssd1 vccd1 vccd1 _5482_/Y sky130_fd_sc_hd__nor2_1
X_4433_ hold229/X _4007_/X _4437_/S vssd1 vssd1 vccd1 vccd1 _4433_/X sky130_fd_sc_hd__mux2_1
X_4364_ hold53/X hold95/X hold91/X hold105/X _4384_/S _5673_/C1 vssd1 vssd1 vccd1
+ vccd1 _4364_/X sky130_fd_sc_hd__mux4_1
X_3315_ _3573_/A _4214_/A _5574_/A vssd1 vssd1 vccd1 vccd1 _3315_/Y sky130_fd_sc_hd__a21oi_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6103_ _6331_/CLK hold78/X vssd1 vssd1 vccd1 vccd1 hold77/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4295_ _6269_/Q _3073_/Y _4305_/S vssd1 vssd1 vccd1 vccd1 _4295_/X sky130_fd_sc_hd__mux2_1
X_3246_ _5294_/B _5322_/C _3246_/C _3244_/X vssd1 vssd1 vccd1 vccd1 _3247_/C sky130_fd_sc_hd__or4b_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6034_ _5492_/Y _6054_/B _6057_/B _4938_/B vssd1 vssd1 vccd1 vccd1 _6034_/X sky130_fd_sc_hd__o2bb2a_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3177_ _3177_/A _3177_/B _3177_/C _3177_/D vssd1 vssd1 vccd1 vccd1 _3197_/B sky130_fd_sc_hd__or4_1
XFILLER_0_83_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5818_ _6377_/Q _5819_/B vssd1 vssd1 vccd1 vccd1 _5836_/A sky130_fd_sc_hd__and2_1
XFILLER_0_91_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5749_ _6319_/Q _5825_/S _5850_/B1 _5748_/X _4319_/X vssd1 vssd1 vccd1 vccd1 _5749_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_32_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4868__A1 _6324_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold571 _3637_/X vssd1 vssd1 vccd1 vccd1 _3638_/C sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout91_A _5029_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold560 _6367_/Q vssd1 vssd1 vccd1 vccd1 hold560/X sky130_fd_sc_hd__buf_1
Xhold582 _5348_/X vssd1 vssd1 vccd1 vccd1 _6312_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold593 _5447_/X vssd1 vssd1 vccd1 vccd1 _6324_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5817__B1 _5735_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4674__S _4674_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5348__A2 _5347_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4849__S _5058_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3531__A1 _5560_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3531__B2 _3528_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3054__A _6243_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3100_ _3656_/A _3100_/B vssd1 vssd1 vccd1 vccd1 _4223_/B sky130_fd_sc_hd__nand2_4
XANTENNA__5808__B1 _5735_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4080_ _6246_/Q _6248_/Q _4135_/S vssd1 vssd1 vccd1 vccd1 _5211_/D sky130_fd_sc_hd__mux2_2
XANTENNA__4584__S _4604_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4982_ _6329_/Q _4981_/C _6330_/Q vssd1 vssd1 vccd1 vccd1 _4983_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_92_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_3_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6414_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_3933_ _3934_/B _3934_/C _4009_/A vssd1 vssd1 vccd1 vccd1 _3935_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__4613__A input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3864_ _3864_/A _3864_/B vssd1 vssd1 vccd1 vccd1 _5249_/B sky130_fd_sc_hd__or2_2
X_5603_ _5603_/A _5603_/B _5603_/C _5603_/D vssd1 vssd1 vccd1 vccd1 _5603_/X sky130_fd_sc_hd__and4_2
X_3795_ _3863_/A _3850_/B _3861_/S vssd1 vssd1 vccd1 vccd1 _4501_/A sky130_fd_sc_hd__or3_4
X_5534_ _5521_/B _5524_/B _5519_/X vssd1 vssd1 vccd1 vccd1 _5535_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_5_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5465_ _5554_/A _5465_/B vssd1 vssd1 vccd1 vccd1 _5466_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_41_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4416_ _4416_/A _4416_/B vssd1 vssd1 vccd1 vccd1 _5251_/B sky130_fd_sc_hd__xnor2_1
X_5396_ _5450_/A _5395_/B _5395_/C vssd1 vssd1 vccd1 vccd1 _5397_/B sky130_fd_sc_hd__a21o_1
X_4347_ _5270_/A _5270_/B _4347_/C vssd1 vssd1 vccd1 vccd1 _5326_/C sky130_fd_sc_hd__or3_1
XANTENNA__5356__A1_N _5578_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5275__A1 _5096_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4278_ _3566_/A _4247_/X _4277_/X _5952_/A vssd1 vssd1 vccd1 vccd1 _5603_/B sky130_fd_sc_hd__a22o_4
XFILLER_0_94_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3229_ _3281_/A _5293_/A _5294_/A _3212_/X vssd1 vssd1 vccd1 vccd1 _3247_/B sky130_fd_sc_hd__or4b_1
XANTENNA__4361__C_N _4633_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4494__S _4500_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6017_ _6057_/A _6016_/X _6026_/B vssd1 vssd1 vccd1 vccd1 _6017_/X sky130_fd_sc_hd__o21a_1
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4523__A _5740_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3838__S _3838_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_hold403_A _6288_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4553__A3 _4767_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5750__A2 _5728_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4669__S _4674_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4936__S1 _5052_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold390 _4992_/X vssd1 vssd1 vccd1 vccd1 _6286_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3602__A _5560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3816__A2 _3715_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3580_ _3580_/A vssd1 vssd1 vccd1 vccd1 _3580_/Y sky130_fd_sc_hd__inv_2
XANTENNA__5741__A2 _5932_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3752__A1 _5217_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4579__S _4604_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5264__A _5317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5250_ _5250_/A _5250_/B _5250_/C _4396_/B vssd1 vssd1 vccd1 vccd1 _5251_/C sky130_fd_sc_hd__or4b_1
X_4201_ hold169/X _4198_/B _4200_/S hold165/X _5676_/C1 vssd1 vssd1 vccd1 vccd1 _4201_/X
+ sky130_fd_sc_hd__o221a_1
X_5181_ hold599/X _5180_/X _5447_/S vssd1 vssd1 vccd1 vccd1 _6294_/D sky130_fd_sc_hd__mux2_1
X_4132_ _4177_/B _4132_/B vssd1 vssd1 vccd1 vccd1 _4132_/Y sky130_fd_sc_hd__xnor2_1
X_4063_ _3741_/X _4061_/A _4062_/X _5087_/B vssd1 vssd1 vccd1 vccd1 _4063_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3512__A _4639_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5203__S _5347_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3807__A2 _3779_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4965_ _5061_/A1 _4962_/X _4964_/X _4867_/B vssd1 vssd1 vccd1 vccd1 _4965_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_19_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3916_ _3917_/B vssd1 vssd1 vccd1 vccd1 _3916_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_80_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4896_ hold371/X _4895_/X _4916_/S vssd1 vssd1 vccd1 vccd1 _4896_/X sky130_fd_sc_hd__mux2_1
X_3847_ hold67/X hold167/X _3861_/S vssd1 vssd1 vccd1 vccd1 _3848_/C sky130_fd_sc_hd__mux2_1
XFILLER_0_6_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5193__A0 _6272_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3778_ _4394_/A vssd1 vssd1 vccd1 vccd1 _4156_/A sky130_fd_sc_hd__inv_2
X_5517_ _5514_/A _5516_/X _6060_/S vssd1 vssd1 vccd1 vccd1 _5517_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4489__S _4491_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4918__S1 _5358_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5448_ _5715_/A _6422_/Q vssd1 vssd1 vccd1 vccd1 _5450_/B sky130_fd_sc_hd__or2_1
Xfanout100 _4639_/B vssd1 vssd1 vccd1 vccd1 _5584_/A1 sky130_fd_sc_hd__buf_2
Xfanout111 _5236_/S vssd1 vssd1 vccd1 vccd1 _5560_/A sky130_fd_sc_hd__clkbuf_8
Xfanout122 hold612/X vssd1 vssd1 vccd1 vccd1 _5560_/B sky130_fd_sc_hd__buf_4
X_5379_ _5472_/S _5375_/X _5378_/X hold573/X vssd1 vssd1 vccd1 vccd1 _5379_/X sky130_fd_sc_hd__a22o_1
Xfanout144 _3482_/A vssd1 vssd1 vccd1 vccd1 _5226_/A sky130_fd_sc_hd__buf_4
Xfanout155 hold659/X vssd1 vssd1 vccd1 vccd1 _4744_/A sky130_fd_sc_hd__buf_2
Xfanout133 hold663/X vssd1 vssd1 vccd1 vccd1 _5358_/A0 sky130_fd_sc_hd__buf_6
Xfanout177 fanout178/X vssd1 vssd1 vccd1 vccd1 fanout177/X sky130_fd_sc_hd__clkbuf_8
Xfanout166 fanout167/X vssd1 vssd1 vccd1 vccd1 fanout166/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_96_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6260__RESET_B fanout177/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5863__A1_N _5932_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5349__A _5603_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3982__A1 _6292_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5031__S0 _5051_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3498__B1 _5258_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5239__A1 _6298_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output35_A _6289_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4862__S _5053_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4750_ _6405_/Q _4750_/B vssd1 vssd1 vccd1 vccd1 _4751_/B sky130_fd_sc_hd__and2_2
XFILLER_0_55_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3701_ _4197_/B _4391_/A2 _3699_/Y _6335_/Q vssd1 vssd1 vccd1 vccd1 _3701_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_55_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4681_ _4520_/Y _4680_/X _5740_/A vssd1 vssd1 vccd1 vccd1 _4681_/X sky130_fd_sc_hd__a21o_2
X_3632_ _6432_/Q _3632_/B _5158_/B _3473_/A vssd1 vssd1 vccd1 vccd1 _3638_/A sky130_fd_sc_hd__or4b_1
X_6420_ _6432_/CLK _6420_/D fanout175/X vssd1 vssd1 vccd1 vccd1 _6420_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_3_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6351_ _6351_/CLK hold8/X vssd1 vssd1 vccd1 vccd1 hold7/A sky130_fd_sc_hd__dfxtp_1
X_5302_ _3581_/A _4347_/C _4349_/C _5273_/X vssd1 vssd1 vccd1 vccd1 _5302_/X sky130_fd_sc_hd__a211o_1
X_3563_ _3562_/X _3561_/X _3548_/Y _3544_/X vssd1 vssd1 vccd1 vccd1 _6487_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_70_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3494_ _6297_/Q _3494_/B vssd1 vssd1 vccd1 vccd1 _3494_/X sky130_fd_sc_hd__or2_1
XFILLER_0_3_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6282_ _6368_/CLK _6282_/D fanout169/X vssd1 vssd1 vccd1 vccd1 _6282_/Q sky130_fd_sc_hd__dfrtp_1
X_5233_ _4143_/Y _5232_/X _5243_/S vssd1 vssd1 vccd1 vccd1 _5233_/X sky130_fd_sc_hd__mux2_1
X_5164_ _5164_/A _5164_/B vssd1 vssd1 vccd1 vccd1 _5165_/B sky130_fd_sc_hd__xnor2_1
X_4115_ _4115_/A _4115_/B vssd1 vssd1 vccd1 vccd1 _4115_/X sky130_fd_sc_hd__xor2_1
XANTENNA__6089__RESET_B fanout174/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5095_ _4070_/A _5094_/X _5447_/S vssd1 vssd1 vccd1 vccd1 _6291_/D sky130_fd_sc_hd__mux2_1
XANTENNA__4057__B _6341_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4046_ _6305_/Q _4046_/B _4046_/C vssd1 vssd1 vccd1 vccd1 _4046_/X sky130_fd_sc_hd__and3_1
XFILLER_0_78_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5402__A1 input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5997_ _5560_/D _5996_/X _6026_/B vssd1 vssd1 vccd1 vccd1 _5997_/X sky130_fd_sc_hd__o21a_1
XANTENNA__4073__A _6246_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3413__B1 _4767_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4948_ _6380_/Q _4754_/X _4940_/X _4947_/X vssd1 vssd1 vccd1 vccd1 _4948_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_74_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4879_ _6190_/Q _6150_/Q _6134_/Q _6213_/Q _5358_/A0 _4326_/B vssd1 vssd1 vccd1 vccd1
+ _4879_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_61_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4520__B _4520_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5469__A1 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5013__S0 _5358_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold470_A _6245_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4248__A _4255_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3955__B2 _6338_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5229__D _6420_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5526__B _6057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4380__A1 _4382_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5632__A1 _5695_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5920_ _5929_/A1 _5919_/X _5034_/Y vssd1 vssd1 vccd1 vccd1 _5920_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_88_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5851_ _5929_/A1 _5850_/X _4920_/Y vssd1 vssd1 vccd1 vccd1 _5851_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_8_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4802_ _4298_/B _4313_/C _4801_/X vssd1 vssd1 vccd1 vccd1 _4802_/X sky130_fd_sc_hd__a21bo_1
X_5782_ _5782_/A _5782_/B _5780_/X vssd1 vssd1 vccd1 vccd1 _5783_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_71_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4733_ _5931_/S _5029_/S _3477_/X vssd1 vssd1 vccd1 vccd1 _4916_/S sky130_fd_sc_hd__a21oi_2
XANTENNA__4621__A input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6403_ _6403_/CLK _6403_/D fanout180/X vssd1 vssd1 vccd1 vccd1 _6403_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4664_ _6337_/Q _6341_/Q _4674_/S vssd1 vssd1 vccd1 vccd1 _4664_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_43_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3615_ _4541_/B _3615_/B vssd1 vssd1 vccd1 vccd1 _3615_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_71_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4595_ _4094_/Y _4604_/S _4564_/A _4594_/Y vssd1 vssd1 vccd1 vccd1 _4595_/X sky130_fd_sc_hd__o211a_1
X_3546_ _4224_/A _3546_/B vssd1 vssd1 vccd1 vccd1 _3546_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_10_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6334_ _6383_/CLK _6334_/D fanout168/X vssd1 vssd1 vccd1 vccd1 _6334_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_0_3_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout104_A _6064_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6265_ _6291_/CLK _6265_/D fanout177/X vssd1 vssd1 vccd1 vccd1 _6265_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5216_ _5216_/A _5216_/B _5216_/C _5216_/D vssd1 vssd1 vccd1 vccd1 _5216_/X sky130_fd_sc_hd__or4_1
X_3477_ _5975_/S _5560_/D _5339_/A vssd1 vssd1 vccd1 vccd1 _3477_/X sky130_fd_sc_hd__a21o_2
XFILLER_0_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6196_ _6218_/CLK _6196_/D vssd1 vssd1 vccd1 vccd1 _6196_/Q sky130_fd_sc_hd__dfxtp_1
X_5147_ _6343_/Q _5328_/C _3755_/X _5146_/X vssd1 vssd1 vccd1 vccd1 _5147_/X sky130_fd_sc_hd__a211o_1
X_5078_ _4284_/A _4070_/A _5193_/S vssd1 vssd1 vccd1 vccd1 _5078_/Y sky130_fd_sc_hd__a21oi_1
X_4029_ _5088_/B _4029_/B vssd1 vssd1 vccd1 vccd1 _4031_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_79_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5623__B2 _6381_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5623__A1 _6293_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3700__A _4427_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4831__C1 _5061_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_hold316_A _6249_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5081__B _5740_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5378__B1 _5339_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5971__S _5975_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold208 _4329_/X vssd1 vssd1 vccd1 vccd1 _6091_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3057__A _6245_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3400_ _5265_/A _3400_/B _5313_/A vssd1 vssd1 vccd1 vccd1 _3401_/A sky130_fd_sc_hd__or3b_1
X_4380_ _4382_/C _4375_/X _4378_/X _4379_/Y vssd1 vssd1 vccd1 vccd1 _4380_/X sky130_fd_sc_hd__a22o_2
Xhold219 _4479_/X vssd1 vssd1 vccd1 vccd1 _6180_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3331_ _3525_/B _3334_/C _4135_/S vssd1 vssd1 vccd1 vccd1 _3896_/S sky130_fd_sc_hd__nor3b_2
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3262_ _4541_/A _5578_/A vssd1 vssd1 vccd1 vccd1 _3654_/A sky130_fd_sc_hd__or2_4
X_6050_ _6057_/B _5016_/B _5536_/Y _5992_/Y vssd1 vssd1 vccd1 vccd1 _6050_/X sky130_fd_sc_hd__o22a_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3193_ _3278_/A _3193_/B vssd1 vssd1 vccd1 vccd1 _5270_/B sky130_fd_sc_hd__nor2_2
X_5001_ _6331_/Q _5002_/B vssd1 vssd1 vccd1 vccd1 _5039_/C sky130_fd_sc_hd__and2_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5903_ _6421_/Q _5902_/X _5930_/S vssd1 vssd1 vccd1 vccd1 _5903_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_76_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5834_ _5846_/A _5834_/B vssd1 vssd1 vccd1 vccd1 _5834_/X sky130_fd_sc_hd__or2_1
XFILLER_0_91_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6030__B2 _4920_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5765_ _5765_/A _5766_/B vssd1 vssd1 vccd1 vccd1 _5782_/A sky130_fd_sc_hd__and2_1
XFILLER_0_98_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4716_ _6272_/Q _4681_/X _4715_/X _5371_/A vssd1 vssd1 vccd1 vccd1 _4716_/X sky130_fd_sc_hd__a22o_1
X_5696_ _3079_/Y _5249_/B _5727_/S vssd1 vssd1 vccd1 vccd1 _5697_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_16_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4647_ _5715_/B _4645_/Y _4646_/X hold312/X _4635_/Y vssd1 vssd1 vccd1 vccd1 _4647_/X
+ sky130_fd_sc_hd__o32a_1
XANTENNA__3552__C1 _6389_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6317_ _6399_/CLK _6317_/D fanout173/X vssd1 vssd1 vccd1 vccd1 _6317_/Q sky130_fd_sc_hd__dfrtp_2
X_4578_ _5695_/A1 hold549/X _4546_/Y _4577_/X vssd1 vssd1 vccd1 vccd1 _4578_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4497__S _4500_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3529_ _5347_/A _4639_/B vssd1 vssd1 vccd1 vccd1 _3529_/Y sky130_fd_sc_hd__nand2_1
X_6248_ _6421_/CLK _6248_/D vssd1 vssd1 vccd1 vccd1 _6248_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__3414__B _4284_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6179_ _6410_/CLK _6179_/D vssd1 vssd1 vccd1 vccd1 _6179_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_hold433_A _6314_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_27_wb_clk_i _6404_/CLK vssd1 vssd1 vccd1 vccd1 _6423_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__6021__A1 _6057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold600_A _6296_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4583__A1 _5695_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3605__A _6487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold91 hold91/A vssd1 vssd1 vccd1 vccd1 hold91/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold80 hold80/A vssd1 vssd1 vccd1 vccd1 hold80/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6012__B2 _4843_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3880_ _3078_/Y _3700_/B _4382_/C vssd1 vssd1 vccd1 vccd1 _3880_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_42_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5550_ _6422_/Q _5558_/S _5549_/X vssd1 vssd1 vccd1 vccd1 _5550_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5481_ _5481_/A _5481_/B _5481_/C _5481_/D vssd1 vssd1 vccd1 vccd1 _5482_/B sky130_fd_sc_hd__or4_1
X_4501_ _4501_/A _5959_/B vssd1 vssd1 vccd1 vccd1 _4509_/S sky130_fd_sc_hd__nor2_4
X_4432_ hold220/X _3965_/X _4437_/S vssd1 vssd1 vccd1 vccd1 _4432_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4363_ _4363_/A _5959_/B vssd1 vssd1 vccd1 vccd1 _4428_/S sky130_fd_sc_hd__nor2_4
X_3314_ _3549_/B _3313_/X _3299_/X vssd1 vssd1 vccd1 vccd1 _3318_/C sky130_fd_sc_hd__o21a_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6102_ _6218_/CLK _6102_/D vssd1 vssd1 vccd1 vccd1 _6102_/Q sky130_fd_sc_hd__dfxtp_1
X_4294_ _6064_/S _4294_/B vssd1 vssd1 vccd1 vccd1 _4296_/S sky130_fd_sc_hd__and2_1
X_3245_ _3126_/X _3628_/B _3143_/X _3683_/C vssd1 vssd1 vccd1 vccd1 _3246_/C sky130_fd_sc_hd__a2bb2o_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6033_ _3046_/A _6031_/X _6032_/Y hold520/X _6029_/Y vssd1 vssd1 vccd1 vccd1 _6033_/X
+ sky130_fd_sc_hd__o32a_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3176_ _3216_/A _3373_/A _3171_/Y _3170_/X vssd1 vssd1 vccd1 vccd1 _3177_/D sky130_fd_sc_hd__a31o_1
XFILLER_0_96_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3250__A _5313_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout171_A fanout181/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4801__A2 _5728_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6003__A1 _5339_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4014__B1 _3786_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5817_ _5236_/S _6422_/Q _3580_/A _5735_/X vssd1 vssd1 vccd1 vccd1 _5819_/B sky130_fd_sc_hd__o31a_1
XFILLER_0_44_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5748_ _6319_/Q _5745_/A _5849_/S vssd1 vssd1 vccd1 vccd1 _5748_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_32_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4317__A1 _6064_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5679_ _6385_/Q _5600_/X _5602_/X _6422_/Q vssd1 vssd1 vccd1 vccd1 _5679_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4317__B2 _6273_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold572 _3638_/X vssd1 vssd1 vccd1 vccd1 _6431_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold550 _4578_/X vssd1 vssd1 vccd1 vccd1 _6243_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold561 _5723_/X vssd1 vssd1 vccd1 vccd1 _6367_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold583 _6381_/Q vssd1 vssd1 vccd1 vccd1 _5865_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold594 _6448_/Q vssd1 vssd1 vccd1 vccd1 hold594/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout84_A _4197_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5817__A1 _5236_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3828__B1 _3781_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold648_A _6269_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4690__S _4732_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5348__A3 _5315_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4005__B1 _5597_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4556__A1 _4224_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5753__B1 _5735_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4308__A1 _4309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5808__A1 _5236_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4981_ _6329_/Q _6330_/Q _4981_/C vssd1 vssd1 vccd1 vccd1 _5002_/B sky130_fd_sc_hd__and3_1
XANTENNA__4795__A1 _6417_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3932_ _4394_/A _3917_/B _3876_/X vssd1 vssd1 vccd1 vccd1 _3934_/C sky130_fd_sc_hd__a21o_1
XANTENNA__4613__B _4631_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3863_ _3863_/A _3863_/B vssd1 vssd1 vccd1 vccd1 _3864_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_61_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5602_ _5603_/B _5602_/B _5602_/C vssd1 vssd1 vccd1 vccd1 _5602_/X sky130_fd_sc_hd__and3_2
XFILLER_0_6_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5533_ _5531_/X _5533_/B vssd1 vssd1 vccd1 vccd1 _5535_/A sky130_fd_sc_hd__and2b_1
X_3794_ _3850_/A _3862_/S _3838_/S vssd1 vssd1 vccd1 vccd1 _3794_/X sky130_fd_sc_hd__and3_4
XFILLER_0_81_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5725__A _5725_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5464_ _5554_/A _5465_/B vssd1 vssd1 vccd1 vccd1 _5464_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_41_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5395_ _5450_/A _5395_/B _5395_/C vssd1 vssd1 vccd1 vccd1 _5395_/X sky130_fd_sc_hd__and3_1
X_4415_ _4416_/A _4416_/B vssd1 vssd1 vccd1 vccd1 _4415_/X sky130_fd_sc_hd__and2b_1
X_4346_ _4346_/A _4346_/B vssd1 vssd1 vccd1 vccd1 _5317_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_1_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4277_ _3530_/D _4274_/X _4276_/X _5584_/A1 vssd1 vssd1 vccd1 vccd1 _4277_/X sky130_fd_sc_hd__a22o_1
X_3228_ _3228_/A _3253_/A _3219_/X _3215_/X vssd1 vssd1 vccd1 vccd1 _5294_/A sky130_fd_sc_hd__or4bb_1
X_6016_ _5441_/B _6054_/B _6057_/B _4863_/B vssd1 vssd1 vccd1 vccd1 _6016_/X sky130_fd_sc_hd__o2bb2a_1
X_3159_ _6258_/Q _6257_/Q vssd1 vssd1 vccd1 vccd1 _3159_/Y sky130_fd_sc_hd__nand2b_1
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4235__B1 _3725_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3589__A2 _5733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4523__B _4523_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4538__A1 _6297_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3139__B _4228_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4710__A1 _6271_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold380 _5776_/X vssd1 vssd1 vccd1 vccd1 _6373_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4710__B2 _5029_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold391 _6084_/Q vssd1 vssd1 vccd1 vccd1 _4314_/S sky130_fd_sc_hd__buf_1
XANTENNA__5370__A _6392_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_42_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6440_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_87_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4226__B1 _4221_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5974__A0 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4529__A1 _6272_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3065__A _6295_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4200_ hold149/X hold122/X _4200_/S vssd1 vssd1 vccd1 vccd1 _4200_/X sky130_fd_sc_hd__mux2_1
X_5180_ _3994_/Y _5179_/X _5243_/S vssd1 vssd1 vccd1 vccd1 _5180_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3215__D _3566_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4131_ _4179_/A _4177_/A vssd1 vssd1 vccd1 vccd1 _4132_/B sky130_fd_sc_hd__or2_1
X_4062_ _6247_/Q _6341_/Q _5088_/B vssd1 vssd1 vccd1 vccd1 _4062_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_3_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5662__C1 _5675_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4964_ _6418_/Q _4963_/X _5060_/S vssd1 vssd1 vccd1 vccd1 _4964_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_19_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4232__A3 _3952_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3915_ _3915_/A _3915_/B vssd1 vssd1 vccd1 vccd1 _3917_/B sky130_fd_sc_hd__nor2_2
XANTENNA__5717__A0 _6268_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4895_ _6084_/Q _4894_/X _5029_/S vssd1 vssd1 vccd1 vccd1 _4895_/X sky130_fd_sc_hd__mux2_1
X_3846_ _3862_/S _3844_/X _3845_/X _3863_/A vssd1 vssd1 vccd1 vccd1 _3852_/B sky130_fd_sc_hd__a211o_1
XANTENNA_fanout134_A _4382_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3777_ _5380_/B _5380_/C vssd1 vssd1 vccd1 vccd1 _4394_/A sky130_fd_sc_hd__nor2_8
XFILLER_0_42_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5516_ _6419_/Q _5558_/S _5515_/X vssd1 vssd1 vccd1 vccd1 _5516_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_100_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5447_ hold592/X _5446_/X _5447_/S vssd1 vssd1 vccd1 vccd1 _5447_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_14_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout112 _3040_/Y vssd1 vssd1 vccd1 vccd1 _5236_/S sky130_fd_sc_hd__clkbuf_4
Xfanout101 _3249_/Y vssd1 vssd1 vccd1 vccd1 _4639_/B sky130_fd_sc_hd__buf_4
X_5378_ _5371_/A _5471_/S _5377_/X _5339_/A vssd1 vssd1 vccd1 vccd1 _5378_/X sky130_fd_sc_hd__a31o_1
Xfanout145 hold514/X vssd1 vssd1 vccd1 vccd1 _3482_/A sky130_fd_sc_hd__buf_4
Xfanout156 _6251_/Q vssd1 vssd1 vccd1 vccd1 _3183_/B sky130_fd_sc_hd__buf_6
Xfanout123 hold587/X vssd1 vssd1 vccd1 vccd1 _5935_/A sky130_fd_sc_hd__buf_4
Xfanout134 _4382_/B vssd1 vssd1 vccd1 vccd1 _4198_/B sky130_fd_sc_hd__buf_4
X_4329_ hold207/X _3881_/X _4336_/S vssd1 vssd1 vccd1 vccd1 _4329_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5248__A2 _5247_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout178 fanout181/X vssd1 vssd1 vccd1 vccd1 fanout178/X sky130_fd_sc_hd__buf_4
Xfanout167 fanout168/X vssd1 vssd1 vccd1 vccd1 fanout167/X sky130_fd_sc_hd__buf_4
XFILLER_0_96_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4759__A1 _5365_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4759__B2 _6416_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5184__B2 _6304_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5365__A _5553_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5031__S1 _5052_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3613__A _5560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3670__A1 _5096_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6317__RESET_B fanout173/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3422__A1 _5313_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3422__B2 _5096_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5974__S _5975_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5355__A1_N _3656_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3700_ _4427_/S _3700_/B _3700_/C vssd1 vssd1 vccd1 vccd1 _3700_/X sky130_fd_sc_hd__or3_2
XFILLER_0_83_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4680_ _5931_/S _5192_/S vssd1 vssd1 vccd1 vccd1 _4680_/X sky130_fd_sc_hd__or2_2
XFILLER_0_83_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5175__A1 _6339_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3631_ _3632_/B _5158_/B vssd1 vssd1 vccd1 vccd1 _3631_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_24_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3562_ _5941_/A _4734_/B _3524_/X _5096_/B vssd1 vssd1 vccd1 vccd1 _3562_/X sky130_fd_sc_hd__a31o_1
X_6350_ _6350_/CLK hold4/X vssd1 vssd1 vccd1 vccd1 hold3/A sky130_fd_sc_hd__dfxtp_1
X_5301_ _5317_/A _5298_/X _5300_/X _5584_/A1 vssd1 vssd1 vccd1 vccd1 _5301_/X sky130_fd_sc_hd__o31a_1
XFILLER_0_51_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3493_ _4767_/A _3374_/A _3591_/B _3492_/X vssd1 vssd1 vccd1 vccd1 _3493_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6281_ _6368_/CLK _6281_/D fanout169/X vssd1 vssd1 vccd1 vccd1 _6281_/Q sky130_fd_sc_hd__dfrtp_1
X_5232_ _5242_/S _5228_/X _5231_/Y vssd1 vssd1 vccd1 vccd1 _5232_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_11_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4619__A input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5163_ _5163_/A _5163_/B vssd1 vssd1 vccd1 vccd1 _5164_/B sky130_fd_sc_hd__xnor2_1
X_4114_ _4022_/A _4022_/B _4098_/A _4113_/Y vssd1 vssd1 vccd1 vccd1 _4115_/B sky130_fd_sc_hd__a31o_1
XFILLER_0_75_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5094_ _5243_/S _5085_/Y _5093_/X _5072_/Y vssd1 vssd1 vccd1 vccd1 _5094_/X sky130_fd_sc_hd__a31o_1
X_4045_ _3758_/Y _5219_/A _4044_/X vssd1 vssd1 vccd1 vccd1 _4046_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_78_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5650__A2 _4382_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5996_ _5368_/Y _6054_/B _6057_/B _5365_/C vssd1 vssd1 vccd1 vccd1 _5996_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_19_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5884__S _5932_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4947_ _5061_/A1 _4942_/X _4946_/X _4867_/B vssd1 vssd1 vccd1 vccd1 _4947_/X sky130_fd_sc_hd__a22o_1
X_4878_ hold381/X _4877_/X _5068_/S vssd1 vssd1 vccd1 vccd1 _4878_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5166__B2 _5242_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3829_ _6131_/Q _3789_/X _3791_/X _6410_/Q vssd1 vssd1 vccd1 vccd1 _3829_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_30_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5013__S1 _4326_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4141__A2 _6422_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold630_A _6085_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4264__A _5603_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5969__S _5975_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5632__A2 _3061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4174__A _5217_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5850_ _6327_/Q _5928_/A2 _5850_/B1 _5849_/X vssd1 vssd1 vccd1 vccd1 _5850_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_61_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4801_ _3076_/Y _5728_/D _4799_/Y _4800_/Y _5740_/A vssd1 vssd1 vccd1 vccd1 _4801_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_0_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5781_ _5782_/A _5782_/B _5780_/X vssd1 vssd1 vccd1 vccd1 _5795_/B sky130_fd_sc_hd__o21ba_1
XFILLER_0_44_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4732_ hold619/X _4731_/X _4732_/S vssd1 vssd1 vccd1 vccd1 _6274_/D sky130_fd_sc_hd__mux2_1
XANTENNA__5148__A1 _6340_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4663_ _6052_/A _4673_/B vssd1 vssd1 vccd1 vccd1 _4663_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_56_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4621__B _4631_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3614_ _6087_/Q _6086_/Q _6088_/Q _6089_/Q vssd1 vssd1 vccd1 vccd1 _3615_/B sky130_fd_sc_hd__or4_1
XFILLER_0_71_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6402_ _6423_/CLK _6402_/D fanout178/X vssd1 vssd1 vccd1 vccd1 _6402_/Q sky130_fd_sc_hd__dfrtp_4
X_4594_ _4594_/A _4604_/S vssd1 vssd1 vccd1 vccd1 _4594_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_101_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3545_ _3581_/A _3545_/B vssd1 vssd1 vccd1 vccd1 _4224_/C sky130_fd_sc_hd__and2_1
X_6333_ _6447_/CLK _6333_/D fanout171/X vssd1 vssd1 vccd1 vccd1 _6333_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_12_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4659__A0 _6336_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5733__A _5733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6264_ _6291_/CLK _6264_/D fanout177/X vssd1 vssd1 vccd1 vccd1 _6264_/Q sky130_fd_sc_hd__dfrtp_1
X_3476_ _5553_/S _6425_/Q _3473_/A _4309_/A vssd1 vssd1 vccd1 vccd1 _3476_/Y sky130_fd_sc_hd__o31ai_1
X_5215_ _5215_/A _5215_/B vssd1 vssd1 vccd1 vccd1 _5215_/X sky130_fd_sc_hd__or2_1
XFILLER_0_86_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4349__A _5560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6195_ _6354_/CLK _6195_/D vssd1 vssd1 vccd1 vccd1 _6195_/Q sky130_fd_sc_hd__dfxtp_1
X_5146_ _6342_/Q _4255_/B _3988_/B _6339_/Q _5145_/X vssd1 vssd1 vccd1 vccd1 _5146_/X
+ sky130_fd_sc_hd__a221o_1
X_5077_ _5077_/A _5077_/B vssd1 vssd1 vccd1 vccd1 _5193_/S sky130_fd_sc_hd__nand2_4
X_4028_ _5087_/A _6340_/Q vssd1 vssd1 vccd1 vccd1 _4031_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_66_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5979_ _5979_/A _5982_/S vssd1 vssd1 vccd1 vccd1 _5979_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_19_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3862__S _3862_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4362__A2 _5597_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4993__S0 _5051_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3570__B1 _4637_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5311__A1 _5258_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3163__A _3573_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4693__S _4727_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5614__A2 _4198_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5378__A1 _5371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3928__A2 _3715_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5029__S _5029_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5550__A1 _6422_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold209 _6216_/Q vssd1 vssd1 vccd1 vccd1 hold209/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4868__S _6315_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3330_ _5715_/C _3494_/B _6297_/Q vssd1 vssd1 vccd1 vccd1 _3330_/X sky130_fd_sc_hd__mux2_1
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3261_ _5096_/A _5265_/A vssd1 vssd1 vccd1 vccd1 _4270_/B sky130_fd_sc_hd__nor2_2
XANTENNA__4105__A2 _3784_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5000_ _4996_/B _4999_/X _5058_/S vssd1 vssd1 vccd1 vccd1 _5000_/X sky130_fd_sc_hd__mux2_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3192_ _3525_/A _4522_/B _5303_/A _3220_/A vssd1 vssd1 vccd1 vccd1 _3510_/B sky130_fd_sc_hd__nor4_4
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3632__D_N _3473_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5066__A0 _6423_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6332__RESET_B fanout168/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3616__B2 _6389_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3616__A1 _6390_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5902_ _5929_/A1 _5901_/X _5016_/Y vssd1 vssd1 vccd1 vccd1 _5902_/X sky130_fd_sc_hd__a21bo_1
X_5833_ _6378_/Q _5833_/B vssd1 vssd1 vccd1 vccd1 _5834_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_63_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5764_ _5236_/S _6418_/Q _3580_/A _5735_/X vssd1 vssd1 vccd1 vccd1 _5766_/B sky130_fd_sc_hd__o31a_1
XFILLER_0_71_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4715_ _6272_/Q _4680_/X _5075_/B hold466/X vssd1 vssd1 vccd1 vccd1 _4715_/X sky130_fd_sc_hd__a2bb2o_1
X_5695_ _5695_/A1 _4158_/A _5571_/Y _5694_/X vssd1 vssd1 vccd1 vccd1 _5695_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_71_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4646_ _3691_/B _4644_/X _4673_/B vssd1 vssd1 vccd1 vccd1 _4646_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_44_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4577_ hold437/X _4567_/Y _4568_/X hold387/X _4576_/X vssd1 vssd1 vccd1 vccd1 _4577_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_12_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5541__A1 _6057_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6316_ _6399_/CLK _6316_/D fanout173/X vssd1 vssd1 vccd1 vccd1 _6316_/Q sky130_fd_sc_hd__dfrtp_1
X_3528_ _5560_/B _4637_/A vssd1 vssd1 vccd1 vccd1 _3528_/Y sky130_fd_sc_hd__nor2_1
X_3459_ _5935_/A _3459_/B vssd1 vssd1 vccd1 vccd1 _3459_/Y sky130_fd_sc_hd__nand2_1
X_6247_ _6297_/CLK _6247_/D vssd1 vssd1 vccd1 vccd1 _6247_/Q sky130_fd_sc_hd__dfxtp_4
X_6178_ _6414_/CLK _6178_/D vssd1 vssd1 vccd1 vccd1 _6178_/Q sky130_fd_sc_hd__dfxtp_1
X_5129_ _5212_/A _5212_/B vssd1 vssd1 vccd1 vccd1 _5135_/A sky130_fd_sc_hd__xor2_1
XANTENNA__5057__A0 _6386_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3324__C _4070_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3846__A1 _3862_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold70 hold70/A vssd1 vssd1 vccd1 vccd1 hold70/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold92 hold92/A vssd1 vssd1 vccd1 vccd1 hold92/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5048__A0 _6422_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold81 hold81/A vssd1 vssd1 vccd1 vccd1 hold81/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4271__A1 _3656_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3068__A _6418_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5480_ _5560_/A _5733_/A _5480_/C _5480_/D vssd1 vssd1 vccd1 vccd1 _5481_/D sky130_fd_sc_hd__or4_1
X_4500_ _4205_/X hold286/X _4500_/S vssd1 vssd1 vccd1 vccd1 _4500_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_1 _5360_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4431_ hold185/X _3923_/X _4437_/S vssd1 vssd1 vccd1 vccd1 _4431_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4362_ _3682_/X _5597_/B _4391_/A2 _4361_/X _5339_/A vssd1 vssd1 vccd1 vccd1 _5959_/B
+ sky130_fd_sc_hd__a41o_4
X_3313_ _4228_/A _5578_/A vssd1 vssd1 vccd1 vccd1 _3313_/X sky130_fd_sc_hd__or2_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6101_ _6218_/CLK hold64/X vssd1 vssd1 vccd1 vccd1 hold63/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4293_ _4298_/B _4292_/X _6064_/S vssd1 vssd1 vccd1 vccd1 _4293_/X sky130_fd_sc_hd__mux2_1
X_3244_ _3116_/A _4522_/D _3122_/X _3633_/B _3590_/B vssd1 vssd1 vccd1 vccd1 _3244_/X
+ sky130_fd_sc_hd__a41o_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6032_ _6032_/A _6063_/S vssd1 vssd1 vccd1 vccd1 _6032_/Y sky130_fd_sc_hd__nor2_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4627__A input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3175_ _3600_/A _4765_/A _3175_/C vssd1 vssd1 vccd1 vccd1 _3177_/C sky130_fd_sc_hd__or3_1
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5816_ hold552/X _5815_/X _5933_/S vssd1 vssd1 vccd1 vccd1 _5816_/X sky130_fd_sc_hd__mux2_1
X_5747_ _5747_/A vssd1 vssd1 vccd1 vccd1 _5747_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_8_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5762__A1 _5932_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5678_ _5677_/X _5674_/X _4147_/X _4419_/X _5691_/S _5690_/S vssd1 vssd1 vccd1 vccd1
+ _5678_/X sky130_fd_sc_hd__mux4_2
X_4629_ input5/X _4631_/B vssd1 vssd1 vccd1 vccd1 _4629_/X sky130_fd_sc_hd__and2_1
Xhold551 _6425_/Q vssd1 vssd1 vccd1 vccd1 _3577_/A sky130_fd_sc_hd__clkbuf_2
Xhold562 _6437_/Q vssd1 vssd1 vccd1 vccd1 hold562/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold540 _6438_/Q vssd1 vssd1 vccd1 vccd1 hold540/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold573 _6319_/Q vssd1 vssd1 vccd1 vccd1 hold573/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold584 _5875_/X vssd1 vssd1 vccd1 vccd1 _6381_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_49_wb_clk_i_A clkbuf_leaf_6_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold595 _6379_/Q vssd1 vssd1 vccd1 vccd1 _5845_/A sky130_fd_sc_hd__buf_1
XFILLER_0_12_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6254__RESET_B fanout179/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5817__A2 _6422_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout77_A _3718_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4789__C1 _5061_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4971__S _5557_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4253__A1 _5578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5753__A1 _5236_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5505__B2 _5441_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5808__A2 _6421_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3351__A _5096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5042__S _5060_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4447__A _4510_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5977__S _5977_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4881__S _5053_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4980_ _4976_/B _4979_/X _5058_/S vssd1 vssd1 vccd1 vccd1 _4980_/X sky130_fd_sc_hd__mux2_1
X_3931_ _3798_/B _3917_/B _4394_/A vssd1 vssd1 vccd1 vccd1 _3934_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_73_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3862_ _3860_/X _3861_/X _3862_/S vssd1 vssd1 vccd1 vccd1 _3863_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_61_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5601_ _5603_/A _5691_/S vssd1 vssd1 vccd1 vccd1 _5602_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5532_ _5554_/A _5532_/B vssd1 vssd1 vccd1 vccd1 _5533_/B sky130_fd_sc_hd__or2_1
XFILLER_0_14_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3793_ hold207/X _4363_/A _5959_/A hold292/X vssd1 vssd1 vccd1 vccd1 _3793_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_14_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5463_ _6440_/Q _4900_/B _5518_/S vssd1 vssd1 vccd1 vccd1 _5465_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_78_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5394_ _6435_/Q _4807_/X _5553_/S vssd1 vssd1 vccd1 vccd1 _5395_/C sky130_fd_sc_hd__mux2_1
X_4414_ _4111_/A _3818_/Y _3825_/X _3872_/Y vssd1 vssd1 vccd1 vccd1 _4416_/B sky130_fd_sc_hd__a211o_1
XFILLER_0_1_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4345_ hold173/X _4205_/X _4345_/S vssd1 vssd1 vccd1 vccd1 _4345_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_1_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4276_ _3132_/B _4258_/X _4260_/X _4275_/X vssd1 vssd1 vccd1 vccd1 _4276_/X sky130_fd_sc_hd__a211o_1
X_3227_ _3289_/A _3566_/B vssd1 vssd1 vccd1 vccd1 _3253_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_94_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3261__A _5096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6015_ _3046_/A _6013_/X _6014_/Y hold562/X _5995_/Y vssd1 vssd1 vccd1 vccd1 _6015_/X
+ sky130_fd_sc_hd__o32a_1
X_3158_ _6258_/Q _6257_/Q vssd1 vssd1 vccd1 vccd1 _4222_/B sky130_fd_sc_hd__and2b_4
XFILLER_0_96_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3089_ _3525_/B _3334_/C vssd1 vssd1 vccd1 vccd1 _4522_/B sky130_fd_sc_hd__or2_4
XANTENNA__4235__A1 _6256_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5432__A0 _6420_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5983__B2 _3577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5983__A1 _3473_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5735__A1 _5077_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3436__A _5518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_5_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_32_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4171__A0 _5217_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold370 _4312_/X vssd1 vssd1 vccd1 vccd1 _6083_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold381 _6280_/Q vssd1 vssd1 vccd1 vccd1 hold381/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold392 _4317_/X vssd1 vssd1 vccd1 vccd1 _6084_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5370__B _5518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4226__A1 _4228_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6482__A _6487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_11_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6344_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_43_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5037__S _6315_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4130_ _4130_/A _4174_/C vssd1 vssd1 vccd1 vccd1 _4177_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_48_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4061_ _4061_/A _4061_/B vssd1 vssd1 vccd1 vccd1 _4061_/X sky130_fd_sc_hd__or2_1
XFILLER_0_3_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5414__A0 _4284_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4963_ _6329_/Q _4981_/C vssd1 vssd1 vccd1 vccd1 _4963_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_80_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3914_ _6069_/Q _3715_/X _3794_/X _6137_/Q _3913_/X vssd1 vssd1 vccd1 vccd1 _3915_/B
+ sky130_fd_sc_hd__a221o_1
X_4894_ _6325_/Q _4893_/X _5852_/S vssd1 vssd1 vccd1 vccd1 _4894_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_73_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3845_ _6185_/Q _3838_/S _3843_/X _3850_/B vssd1 vssd1 vccd1 vccd1 _3845_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_46_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout127_A _3611_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3776_ _3263_/Y _3677_/Y _3775_/X _5096_/B vssd1 vssd1 vccd1 vccd1 _5380_/C sky130_fd_sc_hd__o211a_2
XFILLER_0_54_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5515_ _6057_/A _5513_/X _5514_/Y _5558_/S vssd1 vssd1 vccd1 vccd1 _5515_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_14_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3256__A _3278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5446_ _6421_/Q _5445_/X _5471_/S vssd1 vssd1 vccd1 vccd1 _5446_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_42_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4786__S _5053_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4153__B1 _3791_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout102 _3725_/B vssd1 vssd1 vccd1 vccd1 _5256_/A sky130_fd_sc_hd__clkbuf_8
Xfanout113 _3039_/Y vssd1 vssd1 vccd1 vccd1 _4541_/B sky130_fd_sc_hd__clkbuf_8
X_5377_ _5377_/A _5442_/S vssd1 vssd1 vccd1 vccd1 _5377_/X sky130_fd_sc_hd__and2_4
XFILLER_0_10_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout146 _4224_/A vssd1 vssd1 vccd1 vccd1 _3549_/A sky130_fd_sc_hd__clkbuf_8
XANTENNA__3900__B1 _6245_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout124 _4214_/A vssd1 vssd1 vccd1 vccd1 _5096_/A sky130_fd_sc_hd__clkbuf_8
Xfanout135 hold667/X vssd1 vssd1 vccd1 vccd1 _4382_/B sky130_fd_sc_hd__clkbuf_8
X_4328_ _4510_/A _4363_/A vssd1 vssd1 vccd1 vccd1 _4336_/S sky130_fd_sc_hd__nor2_4
Xfanout157 _6249_/Q vssd1 vssd1 vccd1 vccd1 _5217_/A sky130_fd_sc_hd__buf_4
X_4259_ _3594_/A _4258_/X _4257_/Y vssd1 vssd1 vccd1 vccd1 _4259_/X sky130_fd_sc_hd__a21o_1
Xfanout179 fanout180/X vssd1 vssd1 vccd1 vccd1 fanout179/X sky130_fd_sc_hd__clkbuf_8
Xfanout168 fanout181/X vssd1 vssd1 vccd1 vccd1 fanout168/X sky130_fd_sc_hd__buf_4
XANTENNA__4087__A _6052_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6435__SET_B fanout171/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4550__A _5578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5365__B _6416_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3166__A _4685_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5381__A _5715_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4696__S _5447_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5175__A2 _3502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3630_ _3630_/A _6404_/Q _3634_/B vssd1 vssd1 vccd1 vccd1 _3630_/X sky130_fd_sc_hd__and3_1
XFILLER_0_50_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4907__C1 _4867_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3561_ _3686_/A _3561_/B _3561_/C vssd1 vssd1 vccd1 vccd1 _3561_/X sky130_fd_sc_hd__and3_1
XANTENNA__4383__B1 _5673_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5300_ _3226_/Y _3313_/X _4260_/A _3573_/A _5299_/X vssd1 vssd1 vccd1 vccd1 _5300_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_11_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4135__A0 _6247_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3492_ _4767_/A _3487_/Y _3505_/B _3491_/X vssd1 vssd1 vccd1 vccd1 _3492_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_59_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6280_ _6368_/CLK _6280_/D fanout169/X vssd1 vssd1 vccd1 vccd1 _6280_/Q sky130_fd_sc_hd__dfrtp_1
X_5231_ _5229_/X _5230_/X _5242_/S vssd1 vssd1 vccd1 vccd1 _5231_/Y sky130_fd_sc_hd__o21ai_1
X_5162_ _6419_/Q _6418_/Q vssd1 vssd1 vccd1 vccd1 _5163_/B sky130_fd_sc_hd__xor2_1
XANTENNA__4619__B _4631_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5093_ _3758_/Y _4172_/C _5089_/X _3759_/A _5092_/X vssd1 vssd1 vccd1 vccd1 _5093_/X
+ sky130_fd_sc_hd__a221o_1
X_4113_ _4019_/B _4095_/B _4394_/A vssd1 vssd1 vccd1 vccd1 _4113_/Y sky130_fd_sc_hd__a21oi_1
X_4044_ _6246_/Q _3761_/A _4043_/X _6340_/Q _4041_/X vssd1 vssd1 vccd1 vccd1 _4044_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3949__A0 _6338_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5995_ _6026_/B _5994_/A _3046_/A vssd1 vssd1 vccd1 vccd1 _5995_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__3413__A2 _3654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4946_ _6417_/Q _4945_/Y _5060_/S vssd1 vssd1 vccd1 vccd1 _4946_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_19_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4877_ _4313_/B _4876_/X _5029_/S vssd1 vssd1 vccd1 vccd1 _4877_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_46_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3828_ hold41/A _3779_/X _3781_/X hold59/A vssd1 vssd1 vccd1 vccd1 _3831_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_6_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4374__B1 _5675_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3759_ _3759_/A _3759_/B vssd1 vssd1 vccd1 vccd1 _5209_/A sky130_fd_sc_hd__or2_1
XANTENNA__4677__A1 _5715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5429_ _5441_/A _5428_/X _5371_/A vssd1 vssd1 vccd1 vccd1 _5429_/X sky130_fd_sc_hd__o21a_1
XANTENNA__5405__S _5447_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4545__A _5725_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6051__B1 _6063_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4601__A1 _6422_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4601__B2 _6273_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5376__A _5975_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3624__A _4901_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4174__B _6248_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4800_ _5054_/A _4788_/B _5728_/D vssd1 vssd1 vccd1 vccd1 _4800_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__6042__B1 _6057_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5780_ _5795_/A _5780_/B vssd1 vssd1 vccd1 vccd1 _5780_/X sky130_fd_sc_hd__or2_1
X_4731_ _4193_/Y _4730_/X _4731_/S vssd1 vssd1 vccd1 vccd1 _4731_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5286__A _5715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4662_ _5715_/B _4658_/Y _4661_/X hold344/X _4635_/Y vssd1 vssd1 vccd1 vccd1 _4662_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_0_43_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6401_ _6401_/CLK _6401_/D fanout178/X vssd1 vssd1 vccd1 vccd1 _6401_/Q sky130_fd_sc_hd__dfrtp_1
X_3613_ _5560_/A _4270_/B _3426_/A vssd1 vssd1 vccd1 vccd1 _5247_/B sky130_fd_sc_hd__or3b_4
XFILLER_0_43_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4593_ _5695_/A1 hold420/X _4546_/Y _4592_/X vssd1 vssd1 vccd1 vccd1 _4593_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3544_ _5097_/B _5265_/B _4745_/B vssd1 vssd1 vccd1 vccd1 _3544_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_10_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6332_ _6383_/CLK _6332_/D fanout168/X vssd1 vssd1 vccd1 vccd1 _6332_/Q sky130_fd_sc_hd__dfrtp_4
X_6263_ _6291_/CLK _6263_/D fanout177/X vssd1 vssd1 vccd1 vccd1 _6263_/Q sky130_fd_sc_hd__dfrtp_1
X_3475_ _5553_/S _6425_/Q _3473_/A _4309_/A vssd1 vssd1 vccd1 vccd1 _3475_/X sky130_fd_sc_hd__o31a_1
XFILLER_0_12_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5214_ _5560_/A _6297_/Q _3985_/A vssd1 vssd1 vccd1 vccd1 _5215_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_86_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4659__A1 _6340_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6194_ _6194_/CLK _6194_/D vssd1 vssd1 vccd1 vccd1 _6194_/Q sky130_fd_sc_hd__dfxtp_1
X_5145_ _6341_/Q _4081_/S _3332_/Y _6336_/Q vssd1 vssd1 vccd1 vccd1 _5145_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_98_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5076_ _5076_/A vssd1 vssd1 vccd1 vccd1 _5076_/Y sky130_fd_sc_hd__inv_2
X_4027_ _6245_/Q _6247_/Q _4135_/S vssd1 vssd1 vccd1 vccd1 _5211_/C sky130_fd_sc_hd__mux2_1
XANTENNA__5084__B2 _5371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4831__A1 _3365_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5978_ _5978_/A _5978_/B vssd1 vssd1 vccd1 vccd1 _5982_/S sky130_fd_sc_hd__or2_4
XFILLER_0_19_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4929_ _6360_/Q _4928_/X _5927_/S vssd1 vssd1 vccd1 vccd1 _4929_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_74_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4993__S1 _4326_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3570__A1 _5097_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3444__A _4901_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5311__A2 _4222_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6024__B1 _6057_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3389__A1 _5096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4050__A2 _6048_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4889__A1 _6422_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4889__B2 _5061_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3354__A _3611_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5838__A0 _6326_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3260_ _4639_/C _3581_/A _3257_/X vssd1 vssd1 vccd1 vccd1 _3260_/Y sky130_fd_sc_hd__a21oi_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3191_ _3137_/Y _3143_/X _3628_/B vssd1 vssd1 vccd1 vccd1 _3196_/B sky130_fd_sc_hd__o21ba_1
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4884__S _4901_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5605__A3 _5598_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5901_ _6332_/Q _5928_/A2 _5928_/B1 _5900_/X vssd1 vssd1 vccd1 vccd1 _5901_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4813__B2 _5061_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4813__A1 _6418_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5832_ _6378_/Q _5926_/A vssd1 vssd1 vccd1 vccd1 _5846_/A sky130_fd_sc_hd__and2_1
XANTENNA__6301__RESET_B fanout179/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5763_ _5755_/A _5742_/Y _5762_/Y _5933_/S vssd1 vssd1 vccd1 vccd1 _5763_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3529__A _5347_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4714_ hold646/X _4713_/X _4732_/S vssd1 vssd1 vccd1 vccd1 _6271_/D sky130_fd_sc_hd__mux2_1
X_5694_ _5694_/A _5694_/B _5694_/C vssd1 vssd1 vccd1 vccd1 _5694_/X sky130_fd_sc_hd__or3_1
X_4645_ _6036_/A _4673_/B vssd1 vssd1 vccd1 vccd1 _4645_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_4_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4576_ _6417_/Q _4569_/X _4570_/X _6268_/Q _4575_/X vssd1 vssd1 vccd1 vccd1 _4576_/X
+ sky130_fd_sc_hd__a221o_1
X_3527_ _3522_/X _3523_/X _3526_/X hold101/X _5472_/S vssd1 vssd1 vccd1 vccd1 _3527_/X
+ sky130_fd_sc_hd__o32a_1
X_6315_ _6399_/CLK _6315_/D fanout173/X vssd1 vssd1 vccd1 vccd1 _6315_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_clkbuf_leaf_39_wb_clk_i_A clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_3458_ hold47/X _3449_/X _3457_/X vssd1 vssd1 vccd1 vccd1 hold48/A sky130_fd_sc_hd__a21o_1
X_6246_ _6297_/CLK _6246_/D vssd1 vssd1 vccd1 vccd1 _6246_/Q sky130_fd_sc_hd__dfxtp_4
X_3389_ _5096_/A _3654_/B _3343_/Y vssd1 vssd1 vccd1 vccd1 _3389_/Y sky130_fd_sc_hd__o21ai_1
X_6177_ _6408_/CLK _6177_/D vssd1 vssd1 vccd1 vccd1 _6177_/Q sky130_fd_sc_hd__dfxtp_1
X_5128_ _5128_/A _5128_/B vssd1 vssd1 vccd1 vccd1 _5128_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_98_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5059_ _6334_/Q _5059_/B vssd1 vssd1 vccd1 vccd1 _5059_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_94_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_36_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6290_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__6485__A _6487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3902__A _6245_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold60 hold60/A vssd1 vssd1 vccd1 vccd1 hold60/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 hold82/A vssd1 vssd1 vccd1 vccd1 hold82/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 hold71/A vssd1 vssd1 vccd1 vccd1 hold71/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold93 hold93/A vssd1 vssd1 vccd1 vccd1 hold93/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5548__B _6057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_2 _3501_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4430_ hold278/X _3881_/X _4437_/S vssd1 vssd1 vccd1 vccd1 _4430_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4731__A0 _4193_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4361_ _5069_/A _4361_/B _4633_/C vssd1 vssd1 vccd1 vccd1 _4361_/X sky130_fd_sc_hd__or3b_1
X_6100_ _6217_/CLK hold52/X vssd1 vssd1 vccd1 vccd1 hold51/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__5287__A1 _5715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3312_ _4214_/A _3195_/B _3281_/Y vssd1 vssd1 vccd1 vccd1 _3349_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_67_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4292_ _4290_/Y _4294_/B _6268_/Q _4316_/B vssd1 vssd1 vccd1 vccd1 _4292_/X sky130_fd_sc_hd__a2bb2o_1
X_3243_ _4685_/A _3243_/B vssd1 vssd1 vccd1 vccd1 _3590_/B sky130_fd_sc_hd__or2_2
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6031_ _4313_/C _6030_/X _6063_/S vssd1 vssd1 vccd1 vccd1 _6031_/X sky130_fd_sc_hd__o21a_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3174_ _3148_/X _3152_/Y _3683_/C _3137_/Y vssd1 vssd1 vccd1 vccd1 _3175_/C sky130_fd_sc_hd__a2bb2o_1
XANTENNA__4627__B _4631_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5739__A _5739_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout157_A _6249_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5815_ _5814_/X _5807_/X _5815_/S vssd1 vssd1 vccd1 vccd1 _5815_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_91_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3259__A _5096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4014__A2 _3784_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5746_ _5746_/A _5746_/B vssd1 vssd1 vccd1 vccd1 _5747_/A sky130_fd_sc_hd__or2_4
XFILLER_0_72_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4970__A0 _6418_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5677_ _5677_/A _5677_/B vssd1 vssd1 vccd1 vccd1 _5677_/X sky130_fd_sc_hd__or2_1
XFILLER_0_17_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4628_ _3952_/A _4615_/X _4617_/Y _4627_/X vssd1 vssd1 vccd1 vccd1 _4628_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_44_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold530 _6333_/Q vssd1 vssd1 vccd1 vccd1 _5548_/A sky130_fd_sc_hd__dlygate4sd3_1
X_4559_ _5341_/B _5574_/B _4558_/Y _4556_/X _5096_/A vssd1 vssd1 vccd1 vccd1 _4559_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_12_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold552 _6376_/Q vssd1 vssd1 vccd1 vccd1 hold552/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold541 _6019_/X vssd1 vssd1 vccd1 vccd1 _6438_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold563 _6015_/X vssd1 vssd1 vccd1 vccd1 _6437_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4722__B1 _5075_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold574 _5379_/X vssd1 vssd1 vccd1 vccd1 _6319_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold585 _6321_/Q vssd1 vssd1 vccd1 vccd1 hold585/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold596 _5855_/X vssd1 vssd1 vccd1 vccd1 _6379_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6229_ _6271_/CLK _6229_/D fanout170/X vssd1 vssd1 vccd1 vccd1 _6229_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA__5817__A3 _3580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3828__A2 _3779_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3160__C _4222_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6223__RESET_B fanout179/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4410__C1 _5597_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5753__A2 _6417_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4961__A0 _6381_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5505__A2 _5377_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput50 _6241_/Q vssd1 vssd1 vccd1 vccd1 io_out[5] sky130_fd_sc_hd__buf_12
XANTENNA__5808__A3 _3580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3351__B _4541_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3930_ _4111_/A _3930_/B vssd1 vssd1 vccd1 vccd1 _4009_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_85_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3861_ _6207_/Q _6128_/Q _3861_/S vssd1 vssd1 vccd1 vccd1 _3861_/X sky130_fd_sc_hd__mux2_1
X_5600_ _5603_/B _5603_/C _5610_/B vssd1 vssd1 vccd1 vccd1 _5600_/X sky130_fd_sc_hd__and3_2
XFILLER_0_6_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3792_ _3850_/A _3850_/B _3838_/S vssd1 vssd1 vccd1 vccd1 _5959_/A sky130_fd_sc_hd__or3_1
X_5531_ _5554_/A _5532_/B vssd1 vssd1 vccd1 vccd1 _5531_/X sky130_fd_sc_hd__and2_1
XANTENNA__4952__A0 _6417_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5052__S0 _5358_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5462_ _5715_/A _6423_/Q _5450_/A vssd1 vssd1 vccd1 vccd1 _5475_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_78_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5393_ _6427_/Q _5393_/B vssd1 vssd1 vccd1 vccd1 _5395_/B sky130_fd_sc_hd__nand2_1
X_4413_ hold251/X _4412_/X _4428_/S vssd1 vssd1 vccd1 vccd1 _6133_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_22_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4344_ hold79/X _4148_/X _4345_/S vssd1 vssd1 vccd1 vccd1 hold80/A sky130_fd_sc_hd__mux2_1
XFILLER_0_94_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4275_ _3226_/Y _4208_/B _4257_/Y _3656_/A vssd1 vssd1 vccd1 vccd1 _4275_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5233__S _5243_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6014_ _6048_/A _6026_/B vssd1 vssd1 vccd1 vccd1 _6014_/Y sky130_fd_sc_hd__nor2_1
X_3226_ _3278_/A _3369_/B _3566_/B vssd1 vssd1 vccd1 vccd1 _3226_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__5680__A1 _6297_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3157_ _3290_/B _3220_/A vssd1 vssd1 vccd1 vccd1 _3600_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_27_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4235__A2 _3952_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3088_ _5226_/A _3952_/A vssd1 vssd1 vccd1 vccd1 _3216_/A sky130_fd_sc_hd__nor2_2
XANTENNA__6064__S _6064_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5196__A0 _6341_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5735__A2 _4734_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5729_ _5077_/A _3597_/A _3771_/Y _4748_/X _5728_/X vssd1 vssd1 vccd1 vccd1 _5729_/X
+ sky130_fd_sc_hd__a41o_2
XANTENNA__3717__A _4510_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4312__S _5447_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5499__A1 _4958_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold360 _3540_/X vssd1 vssd1 vccd1 vccd1 _6223_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold371 _6281_/Q vssd1 vssd1 vccd1 vccd1 hold371/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold393 _6082_/Q vssd1 vssd1 vccd1 vccd1 _4304_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold382 _4878_/X vssd1 vssd1 vccd1 vccd1 _6280_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6404__RESET_B fanout180/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold653_A _6268_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5671__A1 _5695_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4283__A _4639_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5098__B _5242_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_51_wb_clk_i clkbuf_leaf_6_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6181_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_23_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3362__A _3611_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5053__S _5053_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4060_ _4059_/A _4059_/B _4061_/A vssd1 vssd1 vccd1 vccd1 _4060_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_3_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5414__A1 _6322_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4905__B _6322_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4962_ _4958_/B _4961_/X _5058_/S vssd1 vssd1 vccd1 vccd1 _4962_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4193__A _6026_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3913_ _6092_/Q _3789_/X _3791_/X _6193_/Q vssd1 vssd1 vccd1 vccd1 _3913_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_19_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4893_ _5773_/A _4892_/X _4882_/Y vssd1 vssd1 vccd1 vccd1 _4893_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_80_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3844_ hold57/A hold75/A _3861_/S vssd1 vssd1 vccd1 vccd1 _3844_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_6_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3775_ _4224_/A _3770_/A _5265_/A vssd1 vssd1 vccd1 vccd1 _3775_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_6_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5514_ _5514_/A _6057_/A vssd1 vssd1 vccd1 vccd1 _5514_/Y sky130_fd_sc_hd__nand2_1
X_5445_ _5441_/Y _5443_/X _5444_/X _5740_/A vssd1 vssd1 vccd1 vccd1 _5445_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_14_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5350__A0 _4382_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout103 _3159_/Y vssd1 vssd1 vccd1 vccd1 _3725_/B sky130_fd_sc_hd__buf_4
XANTENNA__3900__A1 _6243_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5376_ _5975_/S _5376_/B vssd1 vssd1 vccd1 vccd1 _5442_/S sky130_fd_sc_hd__or2_2
XFILLER_0_1_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout147 _6254_/Q vssd1 vssd1 vccd1 vccd1 _4224_/A sky130_fd_sc_hd__clkbuf_8
Xfanout136 _3938_/A vssd1 vssd1 vccd1 vccd1 _5088_/B sky130_fd_sc_hd__clkbuf_8
Xfanout125 _4214_/A vssd1 vssd1 vccd1 vccd1 _4541_/A sky130_fd_sc_hd__clkbuf_8
Xfanout114 _4679_/A vssd1 vssd1 vccd1 vccd1 _3573_/A sky130_fd_sc_hd__buf_8
X_4327_ _5339_/A _4757_/B _4323_/X _4326_/X vssd1 vssd1 vccd1 vccd1 _4327_/X sky130_fd_sc_hd__o31a_1
XFILLER_0_10_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4258_ _3572_/A _3770_/A _3309_/Y _3546_/Y vssd1 vssd1 vccd1 vccd1 _4258_/X sky130_fd_sc_hd__a22o_1
Xfanout158 hold670/X vssd1 vssd1 vccd1 vccd1 _5313_/A sky130_fd_sc_hd__buf_4
Xfanout169 fanout181/X vssd1 vssd1 vccd1 vccd1 fanout169/X sky130_fd_sc_hd__clkbuf_8
X_3209_ _3594_/A _3292_/C vssd1 vssd1 vccd1 vccd1 _3241_/B sky130_fd_sc_hd__nand2_1
XANTENNA__5653__B2 _6420_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5653__A1 _6295_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5898__S _5932_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4189_ _3985_/A _5212_/B _4187_/X _4188_/X vssd1 vssd1 vccd1 vccd1 _4189_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_96_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3416__B1 _5935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold401_A _6287_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3447__A _5935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5365__C _5365_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4392__A1 _4427_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3166__B _3594_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5381__B _6417_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold190 _4507_/X vssd1 vssd1 vccd1 vccd1 _6212_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3655__B1 _5560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4080__A0 _6246_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3560_ _3502_/A _3297_/X _5256_/A vssd1 vssd1 vccd1 vccd1 _3561_/C sky130_fd_sc_hd__a21o_1
XANTENNA__6397__RESET_B fanout174/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6441__SET_B fanout171/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4135__A1 _5217_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3491_ _5313_/A _3491_/B _3541_/A _3639_/B vssd1 vssd1 vccd1 vccd1 _3491_/X sky130_fd_sc_hd__or4b_1
X_5230_ _6419_/Q _6418_/Q _6423_/Q _6422_/Q vssd1 vssd1 vccd1 vccd1 _5230_/X sky130_fd_sc_hd__or4_1
XANTENNA__5572__A _5603_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3894__A0 _6242_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4188__A _6343_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5161_ _6423_/Q _6422_/Q vssd1 vssd1 vccd1 vccd1 _5163_/A sky130_fd_sc_hd__xor2_1
X_5092_ _3985_/A _5091_/X _5241_/S hold304/X _5090_/X vssd1 vssd1 vccd1 vccd1 _5092_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_75_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4112_ _4112_/A _4112_/B vssd1 vssd1 vccd1 vccd1 _4115_/A sky130_fd_sc_hd__nor2_1
X_4043_ _4042_/A _4188_/C _4042_/Y _3746_/X vssd1 vssd1 vccd1 vccd1 _4043_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_38_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3646__B1 _5931_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5994_ _5994_/A vssd1 vssd1 vccd1 vccd1 _5994_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_93_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3949__A1 _6342_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4945_ _4981_/C _4945_/B vssd1 vssd1 vccd1 vccd1 _4945_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_86_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5747__A _5747_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4876_ _6324_/Q _4875_/X _5852_/S vssd1 vssd1 vccd1 vccd1 _4876_/X sky130_fd_sc_hd__mux2_1
X_3827_ _6163_/Q _3784_/X _3786_/X _6171_/Q vssd1 vssd1 vccd1 vccd1 _3831_/A sky130_fd_sc_hd__a22o_1
XANTENNA__3267__A _4255_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3758_ _3759_/A _3759_/B vssd1 vssd1 vccd1 vccd1 _3758_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__4374__A1 _6314_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3689_ _6303_/Q _6301_/Q _5088_/B vssd1 vssd1 vccd1 vccd1 _5196_/S sky130_fd_sc_hd__nand3_4
X_5428_ _5226_/A _6323_/Q _5442_/S vssd1 vssd1 vccd1 vccd1 _5428_/X sky130_fd_sc_hd__mux2_1
X_5359_ _5359_/A _5359_/B vssd1 vssd1 vccd1 vccd1 _5359_/X sky130_fd_sc_hd__or2_1
XANTENNA__5874__B2 _5747_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5874__A1 _5932_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5421__S _5518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4545__B _4568_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6051__A1 _6057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold616_A _6304_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5562__B1 _5315_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4500__S _4500_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output33_A _6288_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3800__B1 _3781_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4730_ _4727_/X _4729_/X _5240_/S vssd1 vssd1 vccd1 vccd1 _4730_/X sky130_fd_sc_hd__mux2_1
X_4661_ _3691_/B _4660_/X _4673_/B vssd1 vssd1 vccd1 vccd1 _4661_/X sky130_fd_sc_hd__o21a_1
X_3612_ _4309_/A _5715_/A _3584_/X _3610_/Y vssd1 vssd1 vccd1 vccd1 _6126_/D sky130_fd_sc_hd__a31o_1
XFILLER_0_71_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6400_ _6423_/CLK _6400_/D fanout178/X vssd1 vssd1 vccd1 vccd1 _6400_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6331_ _6331_/CLK _6331_/D fanout171/X vssd1 vssd1 vccd1 vccd1 _6331_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_3_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4592_ _4564_/A _4589_/X _4591_/X vssd1 vssd1 vccd1 vccd1 _4592_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_101_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3543_ _4541_/B _4734_/B vssd1 vssd1 vccd1 vccd1 _4745_/B sky130_fd_sc_hd__nand2_2
XANTENNA_clkbuf_leaf_29_wb_clk_i_A clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_10_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5506__S _5557_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6262_ _6291_/CLK _6262_/D fanout177/X vssd1 vssd1 vccd1 vccd1 _6262_/Q sky130_fd_sc_hd__dfrtp_1
X_3474_ _5560_/B _5975_/S vssd1 vssd1 vccd1 vccd1 _4615_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_10_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5213_ _5130_/A _5130_/B _5212_/X _5560_/A vssd1 vssd1 vccd1 vccd1 _5215_/A sky130_fd_sc_hd__o31a_1
XFILLER_0_86_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6193_ _6217_/CLK _6193_/D vssd1 vssd1 vccd1 vccd1 _6193_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_2_2__f_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5144_ _6337_/Q _3896_/S _3953_/B _6338_/Q vssd1 vssd1 vccd1 vccd1 _5144_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5608__A1 _6379_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5075_ _5931_/S _5075_/B vssd1 vssd1 vccd1 vccd1 _5076_/A sky130_fd_sc_hd__or2_1
X_4026_ _5122_/A vssd1 vssd1 vccd1 vccd1 _5219_/A sky130_fd_sc_hd__inv_2
XFILLER_0_79_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4292__B1 _6268_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5977_ _3443_/A _5976_/X _5977_/S vssd1 vssd1 vccd1 vccd1 _5977_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_59_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4928_ _6379_/Q _4754_/X _4922_/X _4927_/X vssd1 vssd1 vccd1 vccd1 _4928_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_74_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4859_ hold319/X _5068_/S _4857_/X _4858_/X vssd1 vssd1 vccd1 vccd1 _4859_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_34_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3725__A _5560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6024__B2 _4900_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5378__A3 _5377_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3354__B _3632_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5838__A1 _6378_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3190_ _4685_/A _3594_/A _3290_/B vssd1 vssd1 vccd1 vccd1 _3628_/B sky130_fd_sc_hd__or3_2
XANTENNA__6272__SET_B fanout177/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5900_ _6365_/Q _6384_/Q _5927_/S vssd1 vssd1 vccd1 vccd1 _5900_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_88_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5831_ _5236_/S _6423_/Q _3580_/A _5735_/X vssd1 vssd1 vccd1 vccd1 _5833_/B sky130_fd_sc_hd__o31a_1
XFILLER_0_8_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5762_ _5932_/S _5756_/X _5769_/B _5761_/X vssd1 vssd1 vccd1 vccd1 _5762_/Y sky130_fd_sc_hd__o31ai_1
XANTENNA__3529__B _4639_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4713_ _4049_/Y _4712_/X _4731_/S vssd1 vssd1 vccd1 vccd1 _4713_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_8_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_6_wb_clk_i clkbuf_leaf_6_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6350_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_71_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5693_ _6386_/Q _5600_/X _5602_/X _6423_/Q _5692_/X vssd1 vssd1 vccd1 vccd1 _5694_/C
+ sky130_fd_sc_hd__a221o_1
X_4644_ _4643_/X _6341_/Q _4675_/S vssd1 vssd1 vccd1 vccd1 _4644_/X sky130_fd_sc_hd__mux2_1
X_4575_ _3916_/Y _4604_/S _4564_/A _4574_/Y vssd1 vssd1 vccd1 vccd1 _4575_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_12_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout102_A _3725_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3526_ _4541_/A _3277_/A _3525_/X _3524_/X _5560_/B vssd1 vssd1 vccd1 vccd1 _3526_/X
+ sky130_fd_sc_hd__a311o_1
XANTENNA__5236__S _5236_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6314_ _6351_/CLK _6314_/D vssd1 vssd1 vccd1 vccd1 _6314_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_4_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6245_ _6297_/CLK _6245_/D vssd1 vssd1 vccd1 vccd1 _6245_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5829__B2 _5932_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3457_ _3457_/A _4558_/A _3457_/C vssd1 vssd1 vccd1 vccd1 _3457_/X sky130_fd_sc_hd__and3_1
X_3388_ _4558_/A _6391_/Q _6389_/Q vssd1 vssd1 vccd1 vccd1 _3654_/B sky130_fd_sc_hd__a21oi_2
X_6176_ _6407_/CLK _6176_/D vssd1 vssd1 vccd1 vccd1 _6176_/Q sky130_fd_sc_hd__dfxtp_1
X_5127_ _6292_/Q _4178_/Y _5126_/Y _4179_/A vssd1 vssd1 vccd1 vccd1 _5128_/B sky130_fd_sc_hd__a211o_1
X_5058_ _5054_/B _5057_/X _5058_/S vssd1 vssd1 vccd1 vccd1 _5058_/X sky130_fd_sc_hd__mux2_1
X_4009_ _4009_/A _4009_/B vssd1 vssd1 vccd1 vccd1 _4009_/X sky130_fd_sc_hd__or2_1
XANTENNA__4804__A2 _4752_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3776__C1 _5096_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5935__A _5935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6082__RESET_B fanout169/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3902__B _6295_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4286__A _5226_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold50 hold50/A vssd1 vssd1 vccd1 vccd1 hold50/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3190__A _4685_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold72 hold72/A vssd1 vssd1 vccd1 vccd1 hold72/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 hold83/A vssd1 vssd1 vccd1 vccd1 hold83/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold61 hold61/A vssd1 vssd1 vccd1 vccd1 hold61/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4256__B1 _3725_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold94 hold94/A vssd1 vssd1 vccd1 vccd1 hold94/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4559__B2 _5096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6006__A _6040_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3231__A1 _3183_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_3 _3513_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4360_ hold134/X _4205_/X _4360_/S vssd1 vssd1 vccd1 vccd1 _4360_/X sky130_fd_sc_hd__mux2_1
X_3311_ _3546_/B _3309_/Y _3308_/X _3264_/X _3260_/Y vssd1 vssd1 vccd1 vccd1 _3311_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_0_1_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4895__S _5029_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4291_ _6078_/Q _4298_/B _4287_/B _4316_/B vssd1 vssd1 vccd1 vccd1 _4294_/B sky130_fd_sc_hd__a31o_1
X_3242_ _5292_/B _3242_/B vssd1 vssd1 vccd1 vccd1 _5322_/C sky130_fd_sc_hd__or2_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6030_ _5478_/Y _6054_/B _6057_/B _4920_/B vssd1 vssd1 vccd1 vccd1 _6030_/X sky130_fd_sc_hd__o2bb2a_1
X_3173_ _4210_/A _3502_/A _4222_/B _5941_/A vssd1 vssd1 vccd1 vccd1 _3177_/B sky130_fd_sc_hd__o31a_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5814_ _5821_/B _5814_/B vssd1 vssd1 vccd1 vccd1 _5814_/X sky130_fd_sc_hd__and2b_1
XANTENNA__3259__B _6389_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5745_ _5745_/A _5745_/B vssd1 vssd1 vccd1 vccd1 _5745_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_96_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5676_ _6097_/Q _4198_/B _5676_/B1 _6142_/Q _5676_/C1 vssd1 vssd1 vccd1 vccd1 _5677_/B
+ sky130_fd_sc_hd__o221a_1
X_4627_ input4/X _4631_/B vssd1 vssd1 vccd1 vccd1 _4627_/X sky130_fd_sc_hd__and2_1
Xhold520 _6441_/Q vssd1 vssd1 vccd1 vccd1 hold520/X sky130_fd_sc_hd__dlygate4sd3_1
X_4558_ _4558_/A _5578_/B vssd1 vssd1 vccd1 vccd1 _4558_/Y sky130_fd_sc_hd__nand2_1
Xhold531 _5551_/X vssd1 vssd1 vccd1 vccd1 _6333_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold542 _6386_/Q vssd1 vssd1 vccd1 vccd1 _5925_/A sky130_fd_sc_hd__buf_1
Xhold553 _5816_/X vssd1 vssd1 vccd1 vccd1 _6376_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold597 _6257_/Q vssd1 vssd1 vccd1 vccd1 hold597/X sky130_fd_sc_hd__dlygate4sd3_1
X_3509_ _3337_/B _4734_/B _3418_/A vssd1 vssd1 vccd1 vccd1 _3511_/C sky130_fd_sc_hd__a21oi_1
Xhold564 _6395_/Q vssd1 vssd1 vccd1 vccd1 _5949_/C sky130_fd_sc_hd__buf_1
Xhold586 _5405_/X vssd1 vssd1 vccd1 vccd1 _6321_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold575 _6382_/Q vssd1 vssd1 vccd1 vccd1 _5876_/A sky130_fd_sc_hd__buf_1
X_4489_ hold141/X _4412_/X _4491_/S vssd1 vssd1 vccd1 vccd1 _4489_/X sky130_fd_sc_hd__mux2_1
X_6228_ _6295_/CLK _6228_/D fanout176/X vssd1 vssd1 vccd1 vccd1 _6228_/Q sky130_fd_sc_hd__dfstp_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6159_ _6444_/CLK _6159_/D vssd1 vssd1 vccd1 vccd1 _6159_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4789__A1 _3365_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3169__B _3369_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6263__RESET_B fanout177/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5738__B1 _5735_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3749__C1 _6336_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5753__A3 _3580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5910__B1 _5932_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput40 _6265_/Q vssd1 vssd1 vccd1 vccd1 io_out[25] sky130_fd_sc_hd__buf_12
Xoutput51 _6279_/Q vssd1 vssd1 vccd1 vccd1 io_out[6] sky130_fd_sc_hd__buf_12
XANTENNA__5269__A2 _5715_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4477__A0 _4392_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3632__B _3632_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5977__A0 _3443_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3860_ hold91/A _6184_/Q _3861_/S vssd1 vssd1 vccd1 vccd1 _3860_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3447__D_N _6392_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3791_ _3863_/A _3862_/S _3861_/S vssd1 vssd1 vccd1 vccd1 _3791_/X sky130_fd_sc_hd__and3_4
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5530_ _6446_/Q _5016_/B _5553_/S vssd1 vssd1 vccd1 vccd1 _5532_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_81_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5461_ _5452_/B _5454_/B _5450_/X vssd1 vssd1 vccd1 vccd1 _5467_/A sky130_fd_sc_hd__a21oi_2
XANTENNA__3095__A _3573_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5052__S1 _5052_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4412_ _4427_/S _4411_/X _4410_/X vssd1 vssd1 vccd1 vccd1 _4412_/X sky130_fd_sc_hd__a21o_2
XANTENNA__4704__A1 _6270_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4704__B2 _5371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5392_ hold579/X _5391_/X _5447_/S vssd1 vssd1 vccd1 vccd1 _5392_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_22_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4343_ hold143/X _4102_/X _4345_/S vssd1 vssd1 vccd1 vccd1 _4343_/X sky130_fd_sc_hd__mux2_1
X_4274_ _4274_/A _4274_/B vssd1 vssd1 vccd1 vccd1 _4274_/X sky130_fd_sc_hd__or2_1
XANTENNA__4468__A0 _4392_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3225_ _3566_/A _3566_/B _3254_/A vssd1 vssd1 vccd1 vccd1 _5265_/B sky130_fd_sc_hd__or3b_4
X_6013_ _4313_/C _6012_/X _6026_/B vssd1 vssd1 vccd1 vccd1 _6013_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_94_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3156_ _5325_/A _5560_/C vssd1 vssd1 vccd1 vccd1 _4765_/A sky130_fd_sc_hd__nand2_1
X_3087_ _6258_/Q _6257_/Q vssd1 vssd1 vccd1 vccd1 _3290_/B sky130_fd_sc_hd__nand2_8
XANTENNA__5968__A0 input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3989_ _3992_/A _3987_/X _3988_/X _3746_/X _3985_/X vssd1 vssd1 vccd1 vccd1 _3989_/X
+ sky130_fd_sc_hd__a221o_1
X_5728_ _5728_/A _5728_/B _5728_/C _5728_/D vssd1 vssd1 vccd1 vccd1 _5728_/X sky130_fd_sc_hd__or4_1
XFILLER_0_9_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5659_ _6412_/Q _4198_/B _5676_/B1 _6181_/Q _5675_/C1 vssd1 vssd1 vccd1 vccd1 _5661_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_32_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold350 hold682/X vssd1 vssd1 vccd1 vccd1 _3443_/A sky130_fd_sc_hd__buf_2
Xhold361 _6079_/Q vssd1 vssd1 vccd1 vccd1 _4298_/B sky130_fd_sc_hd__clkbuf_2
Xhold383 _6328_/Q vssd1 vssd1 vccd1 vccd1 hold383/X sky130_fd_sc_hd__buf_1
Xhold394 _4306_/X vssd1 vssd1 vccd1 vccd1 _6082_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold372 _4896_/X vssd1 vssd1 vccd1 vccd1 _6281_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4459__A0 _4392_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_hold646_A _6271_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3419__D1 _5322_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4283__B _4284_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4503__S _4509_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3627__B _3639_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4698__B1 _5075_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3643__A _5931_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5647__C1 _5676_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3673__A1 _5096_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5662__A2 _4382_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4622__B1 _4617_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4961_ _6381_/Q _6329_/Q _6315_/Q vssd1 vssd1 vccd1 vccd1 _4961_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3976__A2 _6245_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3912_ _6109_/Q _3779_/X _3781_/X hold51/A _3911_/X vssd1 vssd1 vccd1 vccd1 _3915_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_19_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4892_ _4891_/X _6325_/Q _5825_/S vssd1 vssd1 vccd1 vccd1 _4892_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_86_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3843_ _3699_/Y _3704_/S _3711_/Y _3712_/X _6145_/Q vssd1 vssd1 vccd1 vccd1 _3843_/X
+ sky130_fd_sc_hd__a311o_1
XANTENNA__4386__C1 _5675_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5509__S _5518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4413__S _4428_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3818__A _4594_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3774_ _3659_/X _3661_/X _3769_/X _3773_/X _3686_/A vssd1 vssd1 vccd1 vccd1 _5380_/B
+ sky130_fd_sc_hd__o311a_2
XFILLER_0_42_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5513_ _6330_/Q _5377_/X _5512_/Y _5377_/A vssd1 vssd1 vccd1 vccd1 _5513_/X sky130_fd_sc_hd__o2bb2a_1
X_5444_ hold592/X input4/X _5469_/S vssd1 vssd1 vccd1 vccd1 _5444_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4153__A2 _3789_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3553__A _5578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5375_ _6416_/Q _5374_/X _5471_/S vssd1 vssd1 vccd1 vccd1 _5375_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4784__S0 _4326_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout104 _6064_/S vssd1 vssd1 vccd1 vccd1 _6060_/S sky130_fd_sc_hd__buf_6
XANTENNA__5244__S _5347_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout137 hold633/X vssd1 vssd1 vccd1 vccd1 _3938_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__3900__A2 _6244_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout126 hold650/X vssd1 vssd1 vccd1 vccd1 _4214_/A sky130_fd_sc_hd__buf_6
Xfanout115 _5553_/S vssd1 vssd1 vccd1 vccd1 _5518_/S sky130_fd_sc_hd__buf_8
X_4326_ _5727_/S _4326_/B vssd1 vssd1 vccd1 vccd1 _4326_/X sky130_fd_sc_hd__or2_1
Xfanout148 _4284_/A vssd1 vssd1 vccd1 vccd1 _3525_/A sky130_fd_sc_hd__buf_4
X_4257_ _4541_/B _4257_/B _5256_/A vssd1 vssd1 vccd1 vccd1 _4257_/Y sky130_fd_sc_hd__nor3_2
Xfanout159 _6116_/Q vssd1 vssd1 vccd1 vccd1 _3686_/A sky130_fd_sc_hd__buf_4
X_3208_ _3278_/A _3220_/A _4679_/C _3525_/A vssd1 vssd1 vccd1 vccd1 _3208_/X sky130_fd_sc_hd__a211o_1
X_4188_ _6343_/Q _5328_/C _4188_/C vssd1 vssd1 vccd1 vccd1 _4188_/X sky130_fd_sc_hd__and3_1
X_3139_ _3656_/A _4228_/A vssd1 vssd1 vccd1 vccd1 _3152_/A sky130_fd_sc_hd__and2b_2
XANTENNA__3664__A1 _3164_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3530__A_N _5560_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3728__A _6304_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5419__S _5447_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3447__B _3451_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4144__A2 _6022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3352__B1 _5158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold180 _4511_/X vssd1 vssd1 vccd1 vccd1 _6215_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold191 hold683/X vssd1 vssd1 vccd1 vccd1 _3507_/C sky130_fd_sc_hd__buf_1
XANTENNA__4294__A _6064_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4080__A1 _6248_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4907__A1 _4809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6014__A _6048_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5580__A1 _3183_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_19_wb_clk_i_A _6404_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3490_ _5472_/S _4287_/B vssd1 vssd1 vccd1 vccd1 _5354_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_59_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3894__A1 _6244_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5160_ _6417_/Q _6416_/Q vssd1 vssd1 vccd1 vccd1 _5164_/A sky130_fd_sc_hd__xor2_1
XANTENNA__3092__B _3183_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5091_ _3573_/A _5217_/A _4183_/Y vssd1 vssd1 vccd1 vccd1 _5091_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_45_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4111_ _4111_/A _4111_/B vssd1 vssd1 vccd1 vccd1 _4112_/B sky130_fd_sc_hd__nor2_1
X_4042_ _4042_/A _4134_/B vssd1 vssd1 vccd1 vccd1 _4042_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_91_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5993_ _6057_/B _5992_/Y _4313_/C vssd1 vssd1 vccd1 vccd1 _5994_/A sky130_fd_sc_hd__a21o_2
X_4944_ _6327_/Q _4943_/C _6328_/Q vssd1 vssd1 vccd1 vccd1 _4945_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_86_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4875_ _5773_/A _4874_/X _4863_/Y vssd1 vssd1 vccd1 vccd1 _4875_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_61_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout132_A _5358_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3826_ _4111_/A _3826_/B vssd1 vssd1 vccd1 vccd1 _4401_/A sky130_fd_sc_hd__xnor2_1
X_3757_ _6303_/Q _3757_/B vssd1 vssd1 vccd1 vccd1 _3759_/B sky130_fd_sc_hd__nand2_2
XANTENNA__3267__B _5258_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4374__A2 _4197_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3688_ _6301_/Q _5088_/B vssd1 vssd1 vccd1 vccd1 _3740_/B sky130_fd_sc_hd__nand2_1
X_5427_ _5441_/A _5427_/B vssd1 vssd1 vccd1 vccd1 _5427_/Y sky130_fd_sc_hd__nand2_1
X_5358_ _5358_/A0 _5357_/Y _5727_/S vssd1 vssd1 vccd1 vccd1 _5358_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_10_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4309_ _4309_/A _4313_/B _4313_/D vssd1 vssd1 vccd1 vccd1 _4310_/C sky130_fd_sc_hd__and3_1
X_5289_ _3237_/A _3135_/X _3246_/C vssd1 vssd1 vccd1 vccd1 _5289_/Y sky130_fd_sc_hd__o21bai_1
XANTENNA__5702__S _6060_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3730__B _6336_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4062__A1 _6247_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3193__A _3278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5078__B1 _5193_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4752__A _6389_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4660_ _4659_/X _6242_/Q _4675_/S vssd1 vssd1 vccd1 vccd1 _4660_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_9_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6295__SET_B fanout177/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3611_ _3611_/A _5715_/A vssd1 vssd1 vccd1 vccd1 _3611_/Y sky130_fd_sc_hd__nand2_1
X_6330_ _6331_/CLK _6330_/D fanout171/X vssd1 vssd1 vccd1 vccd1 _6330_/Q sky130_fd_sc_hd__dfrtp_4
X_4591_ _6437_/Q _4567_/Y _4568_/X hold399/X _4590_/X vssd1 vssd1 vccd1 vccd1 _4591_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_101_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3542_ _5353_/A _5354_/A _5354_/B _5313_/A _3484_/C vssd1 vssd1 vccd1 vccd1 _6118_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_101_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5305__A1 _5313_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6261_ _6291_/CLK _6261_/D fanout177/X vssd1 vssd1 vccd1 vccd1 _6261_/Q sky130_fd_sc_hd__dfrtp_1
X_3473_ _3473_/A _3473_/B vssd1 vssd1 vccd1 vccd1 _5975_/S sky130_fd_sc_hd__nand2_8
XANTENNA__4739__S0 _4326_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5212_ _5212_/A _5212_/B _5212_/C vssd1 vssd1 vccd1 vccd1 _5212_/X sky130_fd_sc_hd__or3_1
X_6192_ _6413_/CLK _6192_/D vssd1 vssd1 vccd1 vccd1 _6192_/Q sky130_fd_sc_hd__dfxtp_1
X_5143_ _5143_/A _5143_/B vssd1 vssd1 vccd1 vccd1 _5143_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_86_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5074_ _3906_/S _5247_/B _4188_/C vssd1 vssd1 vccd1 vccd1 _5102_/B sky130_fd_sc_hd__a21o_2
X_4025_ _4066_/A _4025_/B vssd1 vssd1 vccd1 vccd1 _5122_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_79_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4292__B2 _4316_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4044__A1 _6246_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4044__B2 _6340_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5976_ _6398_/Q _3645_/B _3424_/X _3049_/Y vssd1 vssd1 vccd1 vccd1 _5976_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3278__A _3278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4927_ _5061_/A1 _4924_/X _4926_/X _4867_/B vssd1 vssd1 vccd1 vccd1 _4927_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4595__A2 _4604_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4858_ _6082_/Q _4313_/C _5068_/S vssd1 vssd1 vccd1 vccd1 _4858_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_35_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3809_ _6182_/Q _3715_/X _3794_/X _6213_/Q _3808_/X vssd1 vssd1 vccd1 vccd1 _3810_/B
+ sky130_fd_sc_hd__a221o_1
X_4789_ _3365_/B _4787_/X _4788_/X _5061_/A1 vssd1 vssd1 vccd1 vccd1 _4789_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_15_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3725__B _3725_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3858__A1 _3862_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold461_A _6343_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3188__A _5733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4511__S _4518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5471__A0 _6423_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5578__A _5578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5830_ hold504/X _5829_/X _5933_/S vssd1 vssd1 vccd1 vccd1 _5830_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5728__D _5728_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5761_ _3076_/Y _5728_/D _4800_/Y _5760_/Y _5747_/A vssd1 vssd1 vccd1 vccd1 _5761_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_29_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3098__A _3573_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4712_ _4710_/X _4711_/X _5102_/A vssd1 vssd1 vccd1 vccd1 _4712_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_44_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5692_ _6378_/Q _5603_/X _5691_/X _5594_/Y vssd1 vssd1 vccd1 vccd1 _5692_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_71_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4643_ _6243_/Q _6337_/Q _4674_/S vssd1 vssd1 vccd1 vccd1 _4643_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5517__S _6060_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4574_ _4574_/A _4604_/S vssd1 vssd1 vccd1 vccd1 _4574_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__4421__S _4428_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3525_ _3525_/A _3525_/B _5077_/A _4070_/A vssd1 vssd1 vccd1 vccd1 _3525_/X sky130_fd_sc_hd__and4_1
X_6313_ _6351_/CLK _6313_/D vssd1 vssd1 vccd1 vccd1 _6313_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_24_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6244_ _6421_/CLK _6244_/D vssd1 vssd1 vccd1 vccd1 _6244_/Q sky130_fd_sc_hd__dfxtp_4
X_3456_ _3507_/B _3449_/X _3453_/B _6391_/Q vssd1 vssd1 vccd1 vccd1 _3456_/X sky130_fd_sc_hd__a22o_1
XANTENNA__6310__RESET_B fanout173/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3387_ _3426_/A _3599_/C vssd1 vssd1 vccd1 vccd1 _3387_/X sky130_fd_sc_hd__or2_1
XFILLER_0_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6175_ _6414_/CLK _6175_/D vssd1 vssd1 vccd1 vccd1 _6175_/Q sky130_fd_sc_hd__dfxtp_1
X_5126_ _6292_/Q _5126_/B vssd1 vssd1 vccd1 vccd1 _5126_/Y sky130_fd_sc_hd__nor2_1
X_5057_ _6386_/Q _6334_/Q _6315_/Q vssd1 vssd1 vccd1 vccd1 _5057_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_79_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4008_ _4007_/X hold280/X _4206_/S vssd1 vssd1 vccd1 vccd1 _6071_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_94_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5959_ _5959_/A _5959_/B vssd1 vssd1 vccd1 vccd1 _5967_/S sky130_fd_sc_hd__or2_4
XFILLER_0_75_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4331__S _4336_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4567__A _5339_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4286__B _5715_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold40 hold40/A vssd1 vssd1 vccd1 vccd1 hold40/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3190__B _3594_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold73 hold73/A vssd1 vssd1 vccd1 vccd1 hold73/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 hold51/A vssd1 vssd1 vccd1 vccd1 hold51/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 hold62/A vssd1 vssd1 vccd1 vccd1 hold62/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4256__A1 _3254_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold95 hold95/A vssd1 vssd1 vccd1 vccd1 hold95/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 hold84/A vssd1 vssd1 vccd1 vccd1 hold84/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4506__S _4509_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_45_wb_clk_i clkbuf_leaf_6_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6444_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_85_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6022__A _6022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_4 _4587_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3365__B _3365_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3310_ _5574_/A _4558_/A _5096_/A vssd1 vssd1 vccd1 vccd1 _4268_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4290_ _6078_/Q _4287_/B _4298_/B vssd1 vssd1 vccd1 vccd1 _4290_/Y sky130_fd_sc_hd__a21oi_1
X_3241_ _4679_/D _3241_/B vssd1 vssd1 vccd1 vccd1 _3242_/B sky130_fd_sc_hd__nor2_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3172_ _5935_/A _5265_/A vssd1 vssd1 vccd1 vccd1 _5941_/A sky130_fd_sc_hd__nor2_2
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5813_ _5813_/A _5813_/B _5811_/X vssd1 vssd1 vccd1 vccd1 _5814_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_8_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5744_ _5745_/B _6371_/Q vssd1 vssd1 vccd1 vccd1 _5757_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_72_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5675_ _6198_/Q _4198_/B _5676_/B1 _6074_/Q _5675_/C1 vssd1 vssd1 vccd1 vccd1 _5677_/A
+ sky130_fd_sc_hd__o221a_1
X_4626_ _3525_/B _4615_/X _4617_/Y _4625_/X vssd1 vssd1 vccd1 vccd1 _6255_/D sky130_fd_sc_hd__o22a_1
XFILLER_0_89_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3275__B _3369_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold510 _6384_/Q vssd1 vssd1 vccd1 vccd1 _5905_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4557_ _4558_/A _5578_/B vssd1 vssd1 vccd1 vccd1 _5574_/B sky130_fd_sc_hd__or2_1
Xhold532 _6248_/Q vssd1 vssd1 vccd1 vccd1 hold532/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold543 _5933_/X vssd1 vssd1 vccd1 vccd1 _6386_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold554 _6443_/Q vssd1 vssd1 vccd1 vccd1 hold554/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold521 _6033_/X vssd1 vssd1 vccd1 vccd1 _6441_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3508_ _3453_/B hold326/X _3507_/X _3449_/X _3471_/B vssd1 vssd1 vccd1 vccd1 _3508_/X
+ sky130_fd_sc_hd__a221o_1
Xhold565 _5934_/X vssd1 vssd1 vccd1 vccd1 hold565/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold587 _6393_/Q vssd1 vssd1 vccd1 vccd1 hold587/X sky130_fd_sc_hd__buf_1
Xhold576 _5885_/X vssd1 vssd1 vccd1 vccd1 _6382_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4488_ hold93/X _4405_/X _4491_/S vssd1 vssd1 vccd1 vccd1 hold94/A sky130_fd_sc_hd__mux2_1
Xhold598 _4630_/X vssd1 vssd1 vccd1 vccd1 _6257_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3439_ _3437_/X _3438_/X _3439_/S vssd1 vssd1 vccd1 vccd1 _5981_/B sky130_fd_sc_hd__mux2_1
XANTENNA__4486__A1 _4392_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6227_ _6271_/CLK _6227_/D fanout170/X vssd1 vssd1 vccd1 vccd1 _6227_/Q sky130_fd_sc_hd__dfstp_1
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6158_ _6354_/CLK _6158_/D vssd1 vssd1 vccd1 vccd1 _6158_/Q sky130_fd_sc_hd__dfxtp_1
X_5109_ _5109_/A _5109_/B vssd1 vssd1 vccd1 vccd1 _5115_/A sky130_fd_sc_hd__xnor2_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6089_ _6204_/CLK _6089_/D fanout174/X vssd1 vssd1 vccd1 vccd1 _6089_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__5710__S _6064_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3997__B1 _3786_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3466__A _6390_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput41 _6261_/Q vssd1 vssd1 vccd1 vccd1 io_out[26] sky130_fd_sc_hd__buf_12
Xoutput30 _6285_/Q vssd1 vssd1 vccd1 vccd1 io_out[16] sky130_fd_sc_hd__buf_12
Xoutput52 _6278_/Q vssd1 vssd1 vccd1 vccd1 io_out[7] sky130_fd_sc_hd__buf_12
XANTENNA__3921__B1 _5597_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5729__A1 _5077_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3790_ _3863_/A _3850_/B _3838_/S vssd1 vssd1 vccd1 vccd1 _4363_/A sky130_fd_sc_hd__or3_4
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5460_ hold601/X _5459_/X _5472_/S vssd1 vssd1 vccd1 vccd1 _5460_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5067__S _5557_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3095__B _3278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4411_ hold87/X hold49/X hold228/X hold141/X _5676_/C1 _5676_/B1 vssd1 vssd1 vccd1
+ vccd1 _4411_/X sky130_fd_sc_hd__mux4_2
XFILLER_0_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5391_ _6417_/Q _5390_/X _5471_/S vssd1 vssd1 vccd1 vccd1 _5391_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_10_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3912__B1 _3781_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4342_ hold77/X _4054_/X _4345_/S vssd1 vssd1 vccd1 vccd1 hold78/A sky130_fd_sc_hd__mux2_1
X_4273_ _4273_/A _4273_/B _4273_/C _4273_/D vssd1 vssd1 vccd1 vccd1 _4274_/B sky130_fd_sc_hd__or4_1
X_3224_ _3369_/B _3566_/B vssd1 vssd1 vccd1 vccd1 _3224_/X sky130_fd_sc_hd__or2_2
X_6012_ _5427_/B _6054_/B _6057_/B _4843_/X vssd1 vssd1 vccd1 vccd1 _6012_/X sky130_fd_sc_hd__o2bb2a_1
.ends

