VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO multiplexer
  CLASS BLOCK ;
  FOREIGN multiplexer ;
  ORIGIN 0.000 0.000 ;
  SIZE 200.000 BY 1000.000 ;
  PIN custom_settings[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 4.000 12.880 ;
    END
  END custom_settings[0]
  PIN custom_settings[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.680 4.000 67.280 ;
    END
  END custom_settings[10]
  PIN custom_settings[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.120 4.000 72.720 ;
    END
  END custom_settings[11]
  PIN custom_settings[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 77.560 4.000 78.160 ;
    END
  END custom_settings[12]
  PIN custom_settings[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 4.000 83.600 ;
    END
  END custom_settings[13]
  PIN custom_settings[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END custom_settings[14]
  PIN custom_settings[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.880 4.000 94.480 ;
    END
  END custom_settings[15]
  PIN custom_settings[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 99.320 4.000 99.920 ;
    END
  END custom_settings[16]
  PIN custom_settings[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.760 4.000 105.360 ;
    END
  END custom_settings[17]
  PIN custom_settings[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.200 4.000 110.800 ;
    END
  END custom_settings[18]
  PIN custom_settings[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END custom_settings[19]
  PIN custom_settings[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.720 4.000 18.320 ;
    END
  END custom_settings[1]
  PIN custom_settings[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.080 4.000 121.680 ;
    END
  END custom_settings[20]
  PIN custom_settings[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.520 4.000 127.120 ;
    END
  END custom_settings[21]
  PIN custom_settings[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.960 4.000 132.560 ;
    END
  END custom_settings[22]
  PIN custom_settings[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.400 4.000 138.000 ;
    END
  END custom_settings[23]
  PIN custom_settings[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END custom_settings[24]
  PIN custom_settings[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.280 4.000 148.880 ;
    END
  END custom_settings[25]
  PIN custom_settings[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.720 4.000 154.320 ;
    END
  END custom_settings[26]
  PIN custom_settings[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.160 4.000 159.760 ;
    END
  END custom_settings[27]
  PIN custom_settings[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 164.600 4.000 165.200 ;
    END
  END custom_settings[28]
  PIN custom_settings[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END custom_settings[29]
  PIN custom_settings[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.160 4.000 23.760 ;
    END
  END custom_settings[2]
  PIN custom_settings[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 175.480 4.000 176.080 ;
    END
  END custom_settings[30]
  PIN custom_settings[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.920 4.000 181.520 ;
    END
  END custom_settings[31]
  PIN custom_settings[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.600 4.000 29.200 ;
    END
  END custom_settings[3]
  PIN custom_settings[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END custom_settings[4]
  PIN custom_settings[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 4.000 40.080 ;
    END
  END custom_settings[5]
  PIN custom_settings[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.920 4.000 45.520 ;
    END
  END custom_settings[6]
  PIN custom_settings[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.360 4.000 50.960 ;
    END
  END custom_settings[7]
  PIN custom_settings[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 4.000 56.400 ;
    END
  END custom_settings[8]
  PIN custom_settings[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END custom_settings[9]
  PIN io_in_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 3.770 996.000 4.050 1000.000 ;
    END
  END io_in_0
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 186.360 4.000 186.960 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.760 4.000 241.360 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 246.200 4.000 246.800 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.640 4.000 252.240 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 257.080 4.000 257.680 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 262.520 4.000 263.120 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 267.960 4.000 268.560 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 273.400 4.000 274.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.840 4.000 279.440 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 284.280 4.000 284.880 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.720 4.000 290.320 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.800 4.000 192.400 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.160 4.000 295.760 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 300.600 4.000 301.200 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.040 4.000 306.640 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 311.480 4.000 312.080 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.920 4.000 317.520 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 322.360 4.000 322.960 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 327.800 4.000 328.400 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.240 4.000 333.840 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 338.680 4.000 339.280 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 344.120 4.000 344.720 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.240 4.000 197.840 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 349.560 4.000 350.160 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 355.000 4.000 355.600 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 360.440 4.000 361.040 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 365.880 4.000 366.480 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 371.320 4.000 371.920 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 376.760 4.000 377.360 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 382.200 4.000 382.800 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 387.640 4.000 388.240 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 202.680 4.000 203.280 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 208.120 4.000 208.720 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 213.560 4.000 214.160 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.000 4.000 219.600 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.440 4.000 225.040 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.880 4.000 230.480 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 235.320 4.000 235.920 ;
    END
  END io_oeb[9]
  PIN io_oeb_scrapcpu[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 795.640 4.000 796.240 ;
    END
  END io_oeb_scrapcpu[0]
  PIN io_oeb_scrapcpu[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 850.040 4.000 850.640 ;
    END
  END io_oeb_scrapcpu[10]
  PIN io_oeb_scrapcpu[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 855.480 4.000 856.080 ;
    END
  END io_oeb_scrapcpu[11]
  PIN io_oeb_scrapcpu[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 860.920 4.000 861.520 ;
    END
  END io_oeb_scrapcpu[12]
  PIN io_oeb_scrapcpu[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 866.360 4.000 866.960 ;
    END
  END io_oeb_scrapcpu[13]
  PIN io_oeb_scrapcpu[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 871.800 4.000 872.400 ;
    END
  END io_oeb_scrapcpu[14]
  PIN io_oeb_scrapcpu[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 877.240 4.000 877.840 ;
    END
  END io_oeb_scrapcpu[15]
  PIN io_oeb_scrapcpu[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 882.680 4.000 883.280 ;
    END
  END io_oeb_scrapcpu[16]
  PIN io_oeb_scrapcpu[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 888.120 4.000 888.720 ;
    END
  END io_oeb_scrapcpu[17]
  PIN io_oeb_scrapcpu[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 893.560 4.000 894.160 ;
    END
  END io_oeb_scrapcpu[18]
  PIN io_oeb_scrapcpu[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 899.000 4.000 899.600 ;
    END
  END io_oeb_scrapcpu[19]
  PIN io_oeb_scrapcpu[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 801.080 4.000 801.680 ;
    END
  END io_oeb_scrapcpu[1]
  PIN io_oeb_scrapcpu[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 904.440 4.000 905.040 ;
    END
  END io_oeb_scrapcpu[20]
  PIN io_oeb_scrapcpu[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 909.880 4.000 910.480 ;
    END
  END io_oeb_scrapcpu[21]
  PIN io_oeb_scrapcpu[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 915.320 4.000 915.920 ;
    END
  END io_oeb_scrapcpu[22]
  PIN io_oeb_scrapcpu[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 920.760 4.000 921.360 ;
    END
  END io_oeb_scrapcpu[23]
  PIN io_oeb_scrapcpu[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 926.200 4.000 926.800 ;
    END
  END io_oeb_scrapcpu[24]
  PIN io_oeb_scrapcpu[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 931.640 4.000 932.240 ;
    END
  END io_oeb_scrapcpu[25]
  PIN io_oeb_scrapcpu[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 937.080 4.000 937.680 ;
    END
  END io_oeb_scrapcpu[26]
  PIN io_oeb_scrapcpu[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 942.520 4.000 943.120 ;
    END
  END io_oeb_scrapcpu[27]
  PIN io_oeb_scrapcpu[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 947.960 4.000 948.560 ;
    END
  END io_oeb_scrapcpu[28]
  PIN io_oeb_scrapcpu[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 953.400 4.000 954.000 ;
    END
  END io_oeb_scrapcpu[29]
  PIN io_oeb_scrapcpu[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 806.520 4.000 807.120 ;
    END
  END io_oeb_scrapcpu[2]
  PIN io_oeb_scrapcpu[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 958.840 4.000 959.440 ;
    END
  END io_oeb_scrapcpu[30]
  PIN io_oeb_scrapcpu[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 964.280 4.000 964.880 ;
    END
  END io_oeb_scrapcpu[31]
  PIN io_oeb_scrapcpu[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 969.720 4.000 970.320 ;
    END
  END io_oeb_scrapcpu[32]
  PIN io_oeb_scrapcpu[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 975.160 4.000 975.760 ;
    END
  END io_oeb_scrapcpu[33]
  PIN io_oeb_scrapcpu[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 980.600 4.000 981.200 ;
    END
  END io_oeb_scrapcpu[34]
  PIN io_oeb_scrapcpu[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 986.040 4.000 986.640 ;
    END
  END io_oeb_scrapcpu[35]
  PIN io_oeb_scrapcpu[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 811.960 4.000 812.560 ;
    END
  END io_oeb_scrapcpu[3]
  PIN io_oeb_scrapcpu[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 817.400 4.000 818.000 ;
    END
  END io_oeb_scrapcpu[4]
  PIN io_oeb_scrapcpu[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 822.840 4.000 823.440 ;
    END
  END io_oeb_scrapcpu[5]
  PIN io_oeb_scrapcpu[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 828.280 4.000 828.880 ;
    END
  END io_oeb_scrapcpu[6]
  PIN io_oeb_scrapcpu[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 833.720 4.000 834.320 ;
    END
  END io_oeb_scrapcpu[7]
  PIN io_oeb_scrapcpu[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 839.160 4.000 839.760 ;
    END
  END io_oeb_scrapcpu[8]
  PIN io_oeb_scrapcpu[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 844.600 4.000 845.200 ;
    END
  END io_oeb_scrapcpu[9]
  PIN io_oeb_vliw[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 599.800 4.000 600.400 ;
    END
  END io_oeb_vliw[0]
  PIN io_oeb_vliw[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 654.200 4.000 654.800 ;
    END
  END io_oeb_vliw[10]
  PIN io_oeb_vliw[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 659.640 4.000 660.240 ;
    END
  END io_oeb_vliw[11]
  PIN io_oeb_vliw[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 665.080 4.000 665.680 ;
    END
  END io_oeb_vliw[12]
  PIN io_oeb_vliw[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 670.520 4.000 671.120 ;
    END
  END io_oeb_vliw[13]
  PIN io_oeb_vliw[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 675.960 4.000 676.560 ;
    END
  END io_oeb_vliw[14]
  PIN io_oeb_vliw[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 681.400 4.000 682.000 ;
    END
  END io_oeb_vliw[15]
  PIN io_oeb_vliw[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 686.840 4.000 687.440 ;
    END
  END io_oeb_vliw[16]
  PIN io_oeb_vliw[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 692.280 4.000 692.880 ;
    END
  END io_oeb_vliw[17]
  PIN io_oeb_vliw[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 697.720 4.000 698.320 ;
    END
  END io_oeb_vliw[18]
  PIN io_oeb_vliw[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 703.160 4.000 703.760 ;
    END
  END io_oeb_vliw[19]
  PIN io_oeb_vliw[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 605.240 4.000 605.840 ;
    END
  END io_oeb_vliw[1]
  PIN io_oeb_vliw[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 708.600 4.000 709.200 ;
    END
  END io_oeb_vliw[20]
  PIN io_oeb_vliw[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 714.040 4.000 714.640 ;
    END
  END io_oeb_vliw[21]
  PIN io_oeb_vliw[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 719.480 4.000 720.080 ;
    END
  END io_oeb_vliw[22]
  PIN io_oeb_vliw[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 724.920 4.000 725.520 ;
    END
  END io_oeb_vliw[23]
  PIN io_oeb_vliw[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 730.360 4.000 730.960 ;
    END
  END io_oeb_vliw[24]
  PIN io_oeb_vliw[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 735.800 4.000 736.400 ;
    END
  END io_oeb_vliw[25]
  PIN io_oeb_vliw[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 741.240 4.000 741.840 ;
    END
  END io_oeb_vliw[26]
  PIN io_oeb_vliw[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 746.680 4.000 747.280 ;
    END
  END io_oeb_vliw[27]
  PIN io_oeb_vliw[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 752.120 4.000 752.720 ;
    END
  END io_oeb_vliw[28]
  PIN io_oeb_vliw[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 757.560 4.000 758.160 ;
    END
  END io_oeb_vliw[29]
  PIN io_oeb_vliw[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 610.680 4.000 611.280 ;
    END
  END io_oeb_vliw[2]
  PIN io_oeb_vliw[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 763.000 4.000 763.600 ;
    END
  END io_oeb_vliw[30]
  PIN io_oeb_vliw[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 768.440 4.000 769.040 ;
    END
  END io_oeb_vliw[31]
  PIN io_oeb_vliw[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 773.880 4.000 774.480 ;
    END
  END io_oeb_vliw[32]
  PIN io_oeb_vliw[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 779.320 4.000 779.920 ;
    END
  END io_oeb_vliw[33]
  PIN io_oeb_vliw[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 784.760 4.000 785.360 ;
    END
  END io_oeb_vliw[34]
  PIN io_oeb_vliw[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 790.200 4.000 790.800 ;
    END
  END io_oeb_vliw[35]
  PIN io_oeb_vliw[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 616.120 4.000 616.720 ;
    END
  END io_oeb_vliw[3]
  PIN io_oeb_vliw[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 621.560 4.000 622.160 ;
    END
  END io_oeb_vliw[4]
  PIN io_oeb_vliw[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 627.000 4.000 627.600 ;
    END
  END io_oeb_vliw[5]
  PIN io_oeb_vliw[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 632.440 4.000 633.040 ;
    END
  END io_oeb_vliw[6]
  PIN io_oeb_vliw[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 637.880 4.000 638.480 ;
    END
  END io_oeb_vliw[7]
  PIN io_oeb_vliw[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 643.320 4.000 643.920 ;
    END
  END io_oeb_vliw[8]
  PIN io_oeb_vliw[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 648.760 4.000 649.360 ;
    END
  END io_oeb_vliw[9]
  PIN io_oeb_z80[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 654.200 200.000 654.800 ;
    END
  END io_oeb_z80[0]
  PIN io_oeb_z80[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 695.000 200.000 695.600 ;
    END
  END io_oeb_z80[10]
  PIN io_oeb_z80[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 699.080 200.000 699.680 ;
    END
  END io_oeb_z80[11]
  PIN io_oeb_z80[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 703.160 200.000 703.760 ;
    END
  END io_oeb_z80[12]
  PIN io_oeb_z80[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 707.240 200.000 707.840 ;
    END
  END io_oeb_z80[13]
  PIN io_oeb_z80[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 711.320 200.000 711.920 ;
    END
  END io_oeb_z80[14]
  PIN io_oeb_z80[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 715.400 200.000 716.000 ;
    END
  END io_oeb_z80[15]
  PIN io_oeb_z80[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 719.480 200.000 720.080 ;
    END
  END io_oeb_z80[16]
  PIN io_oeb_z80[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 723.560 200.000 724.160 ;
    END
  END io_oeb_z80[17]
  PIN io_oeb_z80[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 727.640 200.000 728.240 ;
    END
  END io_oeb_z80[18]
  PIN io_oeb_z80[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 731.720 200.000 732.320 ;
    END
  END io_oeb_z80[19]
  PIN io_oeb_z80[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 658.280 200.000 658.880 ;
    END
  END io_oeb_z80[1]
  PIN io_oeb_z80[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 735.800 200.000 736.400 ;
    END
  END io_oeb_z80[20]
  PIN io_oeb_z80[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 739.880 200.000 740.480 ;
    END
  END io_oeb_z80[21]
  PIN io_oeb_z80[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 743.960 200.000 744.560 ;
    END
  END io_oeb_z80[22]
  PIN io_oeb_z80[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 748.040 200.000 748.640 ;
    END
  END io_oeb_z80[23]
  PIN io_oeb_z80[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 752.120 200.000 752.720 ;
    END
  END io_oeb_z80[24]
  PIN io_oeb_z80[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 756.200 200.000 756.800 ;
    END
  END io_oeb_z80[25]
  PIN io_oeb_z80[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 760.280 200.000 760.880 ;
    END
  END io_oeb_z80[26]
  PIN io_oeb_z80[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 764.360 200.000 764.960 ;
    END
  END io_oeb_z80[27]
  PIN io_oeb_z80[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 768.440 200.000 769.040 ;
    END
  END io_oeb_z80[28]
  PIN io_oeb_z80[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 772.520 200.000 773.120 ;
    END
  END io_oeb_z80[29]
  PIN io_oeb_z80[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 662.360 200.000 662.960 ;
    END
  END io_oeb_z80[2]
  PIN io_oeb_z80[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 776.600 200.000 777.200 ;
    END
  END io_oeb_z80[30]
  PIN io_oeb_z80[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 780.680 200.000 781.280 ;
    END
  END io_oeb_z80[31]
  PIN io_oeb_z80[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 784.760 200.000 785.360 ;
    END
  END io_oeb_z80[32]
  PIN io_oeb_z80[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 788.840 200.000 789.440 ;
    END
  END io_oeb_z80[33]
  PIN io_oeb_z80[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 792.920 200.000 793.520 ;
    END
  END io_oeb_z80[34]
  PIN io_oeb_z80[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 797.000 200.000 797.600 ;
    END
  END io_oeb_z80[35]
  PIN io_oeb_z80[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 666.440 200.000 667.040 ;
    END
  END io_oeb_z80[3]
  PIN io_oeb_z80[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 670.520 200.000 671.120 ;
    END
  END io_oeb_z80[4]
  PIN io_oeb_z80[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 674.600 200.000 675.200 ;
    END
  END io_oeb_z80[5]
  PIN io_oeb_z80[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 678.680 200.000 679.280 ;
    END
  END io_oeb_z80[6]
  PIN io_oeb_z80[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 682.760 200.000 683.360 ;
    END
  END io_oeb_z80[7]
  PIN io_oeb_z80[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 686.840 200.000 687.440 ;
    END
  END io_oeb_z80[8]
  PIN io_oeb_z80[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 690.920 200.000 691.520 ;
    END
  END io_oeb_z80[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 54.440 200.000 55.040 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 95.240 200.000 95.840 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 99.320 200.000 99.920 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 103.400 200.000 104.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 107.480 200.000 108.080 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 111.560 200.000 112.160 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 115.640 200.000 116.240 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 119.720 200.000 120.320 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 123.800 200.000 124.400 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 127.880 200.000 128.480 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 131.960 200.000 132.560 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 58.520 200.000 59.120 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 136.040 200.000 136.640 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 140.120 200.000 140.720 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 144.200 200.000 144.800 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 148.280 200.000 148.880 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 152.360 200.000 152.960 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 156.440 200.000 157.040 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 160.520 200.000 161.120 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 164.600 200.000 165.200 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 168.680 200.000 169.280 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 172.760 200.000 173.360 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 62.600 200.000 63.200 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 176.840 200.000 177.440 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 180.920 200.000 181.520 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 185.000 200.000 185.600 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 189.080 200.000 189.680 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 193.160 200.000 193.760 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 197.240 200.000 197.840 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 201.320 200.000 201.920 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 205.400 200.000 206.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 66.680 200.000 67.280 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 70.760 200.000 71.360 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 74.840 200.000 75.440 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 78.920 200.000 79.520 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 83.000 200.000 83.600 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 87.080 200.000 87.680 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 91.160 200.000 91.760 ;
    END
  END io_out[9]
  PIN io_out_scrapcpu[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 801.080 200.000 801.680 ;
    END
  END io_out_scrapcpu[0]
  PIN io_out_scrapcpu[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 841.880 200.000 842.480 ;
    END
  END io_out_scrapcpu[10]
  PIN io_out_scrapcpu[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 845.960 200.000 846.560 ;
    END
  END io_out_scrapcpu[11]
  PIN io_out_scrapcpu[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 850.040 200.000 850.640 ;
    END
  END io_out_scrapcpu[12]
  PIN io_out_scrapcpu[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 854.120 200.000 854.720 ;
    END
  END io_out_scrapcpu[13]
  PIN io_out_scrapcpu[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 858.200 200.000 858.800 ;
    END
  END io_out_scrapcpu[14]
  PIN io_out_scrapcpu[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 862.280 200.000 862.880 ;
    END
  END io_out_scrapcpu[15]
  PIN io_out_scrapcpu[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 866.360 200.000 866.960 ;
    END
  END io_out_scrapcpu[16]
  PIN io_out_scrapcpu[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 870.440 200.000 871.040 ;
    END
  END io_out_scrapcpu[17]
  PIN io_out_scrapcpu[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 874.520 200.000 875.120 ;
    END
  END io_out_scrapcpu[18]
  PIN io_out_scrapcpu[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 878.600 200.000 879.200 ;
    END
  END io_out_scrapcpu[19]
  PIN io_out_scrapcpu[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 805.160 200.000 805.760 ;
    END
  END io_out_scrapcpu[1]
  PIN io_out_scrapcpu[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 882.680 200.000 883.280 ;
    END
  END io_out_scrapcpu[20]
  PIN io_out_scrapcpu[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 886.760 200.000 887.360 ;
    END
  END io_out_scrapcpu[21]
  PIN io_out_scrapcpu[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 890.840 200.000 891.440 ;
    END
  END io_out_scrapcpu[22]
  PIN io_out_scrapcpu[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 894.920 200.000 895.520 ;
    END
  END io_out_scrapcpu[23]
  PIN io_out_scrapcpu[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 899.000 200.000 899.600 ;
    END
  END io_out_scrapcpu[24]
  PIN io_out_scrapcpu[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 903.080 200.000 903.680 ;
    END
  END io_out_scrapcpu[25]
  PIN io_out_scrapcpu[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 907.160 200.000 907.760 ;
    END
  END io_out_scrapcpu[26]
  PIN io_out_scrapcpu[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 911.240 200.000 911.840 ;
    END
  END io_out_scrapcpu[27]
  PIN io_out_scrapcpu[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 915.320 200.000 915.920 ;
    END
  END io_out_scrapcpu[28]
  PIN io_out_scrapcpu[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 919.400 200.000 920.000 ;
    END
  END io_out_scrapcpu[29]
  PIN io_out_scrapcpu[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 809.240 200.000 809.840 ;
    END
  END io_out_scrapcpu[2]
  PIN io_out_scrapcpu[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 923.480 200.000 924.080 ;
    END
  END io_out_scrapcpu[30]
  PIN io_out_scrapcpu[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 927.560 200.000 928.160 ;
    END
  END io_out_scrapcpu[31]
  PIN io_out_scrapcpu[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 931.640 200.000 932.240 ;
    END
  END io_out_scrapcpu[32]
  PIN io_out_scrapcpu[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 935.720 200.000 936.320 ;
    END
  END io_out_scrapcpu[33]
  PIN io_out_scrapcpu[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 939.800 200.000 940.400 ;
    END
  END io_out_scrapcpu[34]
  PIN io_out_scrapcpu[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 943.880 200.000 944.480 ;
    END
  END io_out_scrapcpu[35]
  PIN io_out_scrapcpu[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 813.320 200.000 813.920 ;
    END
  END io_out_scrapcpu[3]
  PIN io_out_scrapcpu[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 817.400 200.000 818.000 ;
    END
  END io_out_scrapcpu[4]
  PIN io_out_scrapcpu[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 821.480 200.000 822.080 ;
    END
  END io_out_scrapcpu[5]
  PIN io_out_scrapcpu[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 825.560 200.000 826.160 ;
    END
  END io_out_scrapcpu[6]
  PIN io_out_scrapcpu[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 829.640 200.000 830.240 ;
    END
  END io_out_scrapcpu[7]
  PIN io_out_scrapcpu[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 833.720 200.000 834.320 ;
    END
  END io_out_scrapcpu[8]
  PIN io_out_scrapcpu[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 837.800 200.000 838.400 ;
    END
  END io_out_scrapcpu[9]
  PIN io_out_vliw[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 13.890 996.000 14.170 1000.000 ;
    END
  END io_out_vliw[0]
  PIN io_out_vliw[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 64.490 996.000 64.770 1000.000 ;
    END
  END io_out_vliw[10]
  PIN io_out_vliw[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 69.550 996.000 69.830 1000.000 ;
    END
  END io_out_vliw[11]
  PIN io_out_vliw[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 74.610 996.000 74.890 1000.000 ;
    END
  END io_out_vliw[12]
  PIN io_out_vliw[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 79.670 996.000 79.950 1000.000 ;
    END
  END io_out_vliw[13]
  PIN io_out_vliw[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 84.730 996.000 85.010 1000.000 ;
    END
  END io_out_vliw[14]
  PIN io_out_vliw[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 89.790 996.000 90.070 1000.000 ;
    END
  END io_out_vliw[15]
  PIN io_out_vliw[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 94.850 996.000 95.130 1000.000 ;
    END
  END io_out_vliw[16]
  PIN io_out_vliw[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 99.910 996.000 100.190 1000.000 ;
    END
  END io_out_vliw[17]
  PIN io_out_vliw[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 104.970 996.000 105.250 1000.000 ;
    END
  END io_out_vliw[18]
  PIN io_out_vliw[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 110.030 996.000 110.310 1000.000 ;
    END
  END io_out_vliw[19]
  PIN io_out_vliw[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 18.950 996.000 19.230 1000.000 ;
    END
  END io_out_vliw[1]
  PIN io_out_vliw[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 115.090 996.000 115.370 1000.000 ;
    END
  END io_out_vliw[20]
  PIN io_out_vliw[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 120.150 996.000 120.430 1000.000 ;
    END
  END io_out_vliw[21]
  PIN io_out_vliw[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 125.210 996.000 125.490 1000.000 ;
    END
  END io_out_vliw[22]
  PIN io_out_vliw[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 130.270 996.000 130.550 1000.000 ;
    END
  END io_out_vliw[23]
  PIN io_out_vliw[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 135.330 996.000 135.610 1000.000 ;
    END
  END io_out_vliw[24]
  PIN io_out_vliw[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 140.390 996.000 140.670 1000.000 ;
    END
  END io_out_vliw[25]
  PIN io_out_vliw[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 145.450 996.000 145.730 1000.000 ;
    END
  END io_out_vliw[26]
  PIN io_out_vliw[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 150.510 996.000 150.790 1000.000 ;
    END
  END io_out_vliw[27]
  PIN io_out_vliw[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 155.570 996.000 155.850 1000.000 ;
    END
  END io_out_vliw[28]
  PIN io_out_vliw[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 160.630 996.000 160.910 1000.000 ;
    END
  END io_out_vliw[29]
  PIN io_out_vliw[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 24.010 996.000 24.290 1000.000 ;
    END
  END io_out_vliw[2]
  PIN io_out_vliw[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 165.690 996.000 165.970 1000.000 ;
    END
  END io_out_vliw[30]
  PIN io_out_vliw[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 170.750 996.000 171.030 1000.000 ;
    END
  END io_out_vliw[31]
  PIN io_out_vliw[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 175.810 996.000 176.090 1000.000 ;
    END
  END io_out_vliw[32]
  PIN io_out_vliw[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 180.870 996.000 181.150 1000.000 ;
    END
  END io_out_vliw[33]
  PIN io_out_vliw[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 185.930 996.000 186.210 1000.000 ;
    END
  END io_out_vliw[34]
  PIN io_out_vliw[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 190.990 996.000 191.270 1000.000 ;
    END
  END io_out_vliw[35]
  PIN io_out_vliw[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 29.070 996.000 29.350 1000.000 ;
    END
  END io_out_vliw[3]
  PIN io_out_vliw[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 34.130 996.000 34.410 1000.000 ;
    END
  END io_out_vliw[4]
  PIN io_out_vliw[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 39.190 996.000 39.470 1000.000 ;
    END
  END io_out_vliw[5]
  PIN io_out_vliw[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 44.250 996.000 44.530 1000.000 ;
    END
  END io_out_vliw[6]
  PIN io_out_vliw[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 49.310 996.000 49.590 1000.000 ;
    END
  END io_out_vliw[7]
  PIN io_out_vliw[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 54.370 996.000 54.650 1000.000 ;
    END
  END io_out_vliw[8]
  PIN io_out_vliw[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 59.430 996.000 59.710 1000.000 ;
    END
  END io_out_vliw[9]
  PIN io_out_z80[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 503.240 200.000 503.840 ;
    END
  END io_out_z80[0]
  PIN io_out_z80[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 544.040 200.000 544.640 ;
    END
  END io_out_z80[10]
  PIN io_out_z80[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 548.120 200.000 548.720 ;
    END
  END io_out_z80[11]
  PIN io_out_z80[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 552.200 200.000 552.800 ;
    END
  END io_out_z80[12]
  PIN io_out_z80[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 556.280 200.000 556.880 ;
    END
  END io_out_z80[13]
  PIN io_out_z80[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 560.360 200.000 560.960 ;
    END
  END io_out_z80[14]
  PIN io_out_z80[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 564.440 200.000 565.040 ;
    END
  END io_out_z80[15]
  PIN io_out_z80[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 568.520 200.000 569.120 ;
    END
  END io_out_z80[16]
  PIN io_out_z80[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 572.600 200.000 573.200 ;
    END
  END io_out_z80[17]
  PIN io_out_z80[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 576.680 200.000 577.280 ;
    END
  END io_out_z80[18]
  PIN io_out_z80[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 580.760 200.000 581.360 ;
    END
  END io_out_z80[19]
  PIN io_out_z80[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 507.320 200.000 507.920 ;
    END
  END io_out_z80[1]
  PIN io_out_z80[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 584.840 200.000 585.440 ;
    END
  END io_out_z80[20]
  PIN io_out_z80[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 588.920 200.000 589.520 ;
    END
  END io_out_z80[21]
  PIN io_out_z80[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 593.000 200.000 593.600 ;
    END
  END io_out_z80[22]
  PIN io_out_z80[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 597.080 200.000 597.680 ;
    END
  END io_out_z80[23]
  PIN io_out_z80[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 601.160 200.000 601.760 ;
    END
  END io_out_z80[24]
  PIN io_out_z80[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 605.240 200.000 605.840 ;
    END
  END io_out_z80[25]
  PIN io_out_z80[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 609.320 200.000 609.920 ;
    END
  END io_out_z80[26]
  PIN io_out_z80[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 613.400 200.000 614.000 ;
    END
  END io_out_z80[27]
  PIN io_out_z80[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 617.480 200.000 618.080 ;
    END
  END io_out_z80[28]
  PIN io_out_z80[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 621.560 200.000 622.160 ;
    END
  END io_out_z80[29]
  PIN io_out_z80[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 511.400 200.000 512.000 ;
    END
  END io_out_z80[2]
  PIN io_out_z80[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 625.640 200.000 626.240 ;
    END
  END io_out_z80[30]
  PIN io_out_z80[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 629.720 200.000 630.320 ;
    END
  END io_out_z80[31]
  PIN io_out_z80[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 633.800 200.000 634.400 ;
    END
  END io_out_z80[32]
  PIN io_out_z80[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 637.880 200.000 638.480 ;
    END
  END io_out_z80[33]
  PIN io_out_z80[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 641.960 200.000 642.560 ;
    END
  END io_out_z80[34]
  PIN io_out_z80[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 646.040 200.000 646.640 ;
    END
  END io_out_z80[35]
  PIN io_out_z80[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 515.480 200.000 516.080 ;
    END
  END io_out_z80[3]
  PIN io_out_z80[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 519.560 200.000 520.160 ;
    END
  END io_out_z80[4]
  PIN io_out_z80[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 523.640 200.000 524.240 ;
    END
  END io_out_z80[5]
  PIN io_out_z80[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 527.720 200.000 528.320 ;
    END
  END io_out_z80[6]
  PIN io_out_z80[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 531.800 200.000 532.400 ;
    END
  END io_out_z80[7]
  PIN io_out_z80[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 535.880 200.000 536.480 ;
    END
  END io_out_z80[8]
  PIN io_out_z80[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 539.960 200.000 540.560 ;
    END
  END io_out_z80[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 340.040 200.000 340.640 ;
    END
  END la_data_out[0]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 380.840 200.000 381.440 ;
    END
  END la_data_out[10]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 384.920 200.000 385.520 ;
    END
  END la_data_out[11]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 389.000 200.000 389.600 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 393.080 200.000 393.680 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 397.160 200.000 397.760 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 401.240 200.000 401.840 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 405.320 200.000 405.920 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 409.400 200.000 410.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 413.480 200.000 414.080 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 417.560 200.000 418.160 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 344.120 200.000 344.720 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 421.640 200.000 422.240 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 425.720 200.000 426.320 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 429.800 200.000 430.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 433.880 200.000 434.480 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 437.960 200.000 438.560 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 442.040 200.000 442.640 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 446.120 200.000 446.720 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 450.200 200.000 450.800 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 454.280 200.000 454.880 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 458.360 200.000 458.960 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 348.200 200.000 348.800 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 462.440 200.000 463.040 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 466.520 200.000 467.120 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 470.600 200.000 471.200 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 474.680 200.000 475.280 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 478.760 200.000 479.360 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 482.840 200.000 483.440 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 486.920 200.000 487.520 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 491.000 200.000 491.600 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 495.080 200.000 495.680 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 499.160 200.000 499.760 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 352.280 200.000 352.880 ;
    END
  END la_data_out[3]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 356.360 200.000 356.960 ;
    END
  END la_data_out[4]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 360.440 200.000 361.040 ;
    END
  END la_data_out[5]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 364.520 200.000 365.120 ;
    END
  END la_data_out[6]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 368.600 200.000 369.200 ;
    END
  END la_data_out[7]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 372.680 200.000 373.280 ;
    END
  END la_data_out[8]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 376.760 200.000 377.360 ;
    END
  END la_data_out[9]
  PIN rst_scrapcpu
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 196.050 996.000 196.330 1000.000 ;
    END
  END rst_scrapcpu
  PIN rst_vliw
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 8.830 996.000 9.110 1000.000 ;
    END
  END rst_vliw
  PIN rst_z80
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 650.120 200.000 650.720 ;
    END
  END rst_z80
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 987.600 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 987.600 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 393.080 4.000 393.680 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 398.520 4.000 399.120 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 594.360 4.000 594.960 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 0.000 7.270 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.790 0.000 67.070 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.770 0.000 73.050 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.750 0.000 79.030 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.730 0.000 85.010 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.710 0.000 90.990 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.670 0.000 102.950 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.650 0.000 108.930 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.630 0.000 114.910 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.610 0.000 120.890 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 126.590 0.000 126.870 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.570 0.000 132.850 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.530 0.000 144.810 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.510 0.000 150.790 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.490 0.000 156.770 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.470 0.000 162.750 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.450 0.000 168.730 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.430 0.000 174.710 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 18.950 0.000 19.230 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.390 0.000 186.670 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.370 0.000 192.650 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 24.930 0.000 25.210 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 30.910 0.000 31.190 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.890 0.000 37.170 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.870 0.000 43.150 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 0.000 49.130 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.810 0.000 61.090 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 583.480 4.000 584.080 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 403.960 4.000 404.560 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 458.360 4.000 458.960 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 463.800 4.000 464.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 469.240 4.000 469.840 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 474.680 4.000 475.280 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 480.120 4.000 480.720 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 485.560 4.000 486.160 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 491.000 4.000 491.600 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 496.440 4.000 497.040 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 501.880 4.000 502.480 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 507.320 4.000 507.920 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 409.400 4.000 410.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 512.760 4.000 513.360 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 518.200 4.000 518.800 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 523.640 4.000 524.240 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 529.080 4.000 529.680 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 534.520 4.000 535.120 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 539.960 4.000 540.560 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 545.400 4.000 546.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 550.840 4.000 551.440 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 556.280 4.000 556.880 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 561.720 4.000 562.320 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 414.840 4.000 415.440 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 567.160 4.000 567.760 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 572.600 4.000 573.200 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 420.280 4.000 420.880 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 425.720 4.000 426.320 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 431.160 4.000 431.760 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 436.600 4.000 437.200 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 442.040 4.000 442.640 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 447.480 4.000 448.080 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 452.920 4.000 453.520 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 209.480 200.000 210.080 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 250.280 200.000 250.880 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 254.360 200.000 254.960 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 258.440 200.000 259.040 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 262.520 200.000 263.120 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 266.600 200.000 267.200 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 270.680 200.000 271.280 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 274.760 200.000 275.360 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 278.840 200.000 279.440 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 282.920 200.000 283.520 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 287.000 200.000 287.600 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 213.560 200.000 214.160 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 291.080 200.000 291.680 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 295.160 200.000 295.760 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 299.240 200.000 299.840 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 303.320 200.000 303.920 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 307.400 200.000 308.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 311.480 200.000 312.080 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 315.560 200.000 316.160 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 319.640 200.000 320.240 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 323.720 200.000 324.320 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 327.800 200.000 328.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 217.640 200.000 218.240 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 331.880 200.000 332.480 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 335.960 200.000 336.560 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 221.720 200.000 222.320 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 225.800 200.000 226.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 229.880 200.000 230.480 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 233.960 200.000 234.560 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 238.040 200.000 238.640 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 242.120 200.000 242.720 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 246.200 200.000 246.800 ;
    END
  END wbs_dat_o[9]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 588.920 4.000 589.520 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 578.040 4.000 578.640 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 194.120 987.445 ;
      LAYER met1 ;
        RECT 0.070 10.640 199.940 987.600 ;
      LAYER met2 ;
        RECT 0.090 995.720 3.490 996.610 ;
        RECT 4.330 995.720 8.550 996.610 ;
        RECT 9.390 995.720 13.610 996.610 ;
        RECT 14.450 995.720 18.670 996.610 ;
        RECT 19.510 995.720 23.730 996.610 ;
        RECT 24.570 995.720 28.790 996.610 ;
        RECT 29.630 995.720 33.850 996.610 ;
        RECT 34.690 995.720 38.910 996.610 ;
        RECT 39.750 995.720 43.970 996.610 ;
        RECT 44.810 995.720 49.030 996.610 ;
        RECT 49.870 995.720 54.090 996.610 ;
        RECT 54.930 995.720 59.150 996.610 ;
        RECT 59.990 995.720 64.210 996.610 ;
        RECT 65.050 995.720 69.270 996.610 ;
        RECT 70.110 995.720 74.330 996.610 ;
        RECT 75.170 995.720 79.390 996.610 ;
        RECT 80.230 995.720 84.450 996.610 ;
        RECT 85.290 995.720 89.510 996.610 ;
        RECT 90.350 995.720 94.570 996.610 ;
        RECT 95.410 995.720 99.630 996.610 ;
        RECT 100.470 995.720 104.690 996.610 ;
        RECT 105.530 995.720 109.750 996.610 ;
        RECT 110.590 995.720 114.810 996.610 ;
        RECT 115.650 995.720 119.870 996.610 ;
        RECT 120.710 995.720 124.930 996.610 ;
        RECT 125.770 995.720 129.990 996.610 ;
        RECT 130.830 995.720 135.050 996.610 ;
        RECT 135.890 995.720 140.110 996.610 ;
        RECT 140.950 995.720 145.170 996.610 ;
        RECT 146.010 995.720 150.230 996.610 ;
        RECT 151.070 995.720 155.290 996.610 ;
        RECT 156.130 995.720 160.350 996.610 ;
        RECT 161.190 995.720 165.410 996.610 ;
        RECT 166.250 995.720 170.470 996.610 ;
        RECT 171.310 995.720 175.530 996.610 ;
        RECT 176.370 995.720 180.590 996.610 ;
        RECT 181.430 995.720 185.650 996.610 ;
        RECT 186.490 995.720 190.710 996.610 ;
        RECT 191.550 995.720 195.770 996.610 ;
        RECT 196.610 995.720 199.940 996.610 ;
        RECT 0.090 4.280 199.940 995.720 ;
        RECT 0.090 3.670 6.710 4.280 ;
        RECT 7.550 3.670 12.690 4.280 ;
        RECT 13.530 3.670 18.670 4.280 ;
        RECT 19.510 3.670 24.650 4.280 ;
        RECT 25.490 3.670 30.630 4.280 ;
        RECT 31.470 3.670 36.610 4.280 ;
        RECT 37.450 3.670 42.590 4.280 ;
        RECT 43.430 3.670 48.570 4.280 ;
        RECT 49.410 3.670 54.550 4.280 ;
        RECT 55.390 3.670 60.530 4.280 ;
        RECT 61.370 3.670 66.510 4.280 ;
        RECT 67.350 3.670 72.490 4.280 ;
        RECT 73.330 3.670 78.470 4.280 ;
        RECT 79.310 3.670 84.450 4.280 ;
        RECT 85.290 3.670 90.430 4.280 ;
        RECT 91.270 3.670 96.410 4.280 ;
        RECT 97.250 3.670 102.390 4.280 ;
        RECT 103.230 3.670 108.370 4.280 ;
        RECT 109.210 3.670 114.350 4.280 ;
        RECT 115.190 3.670 120.330 4.280 ;
        RECT 121.170 3.670 126.310 4.280 ;
        RECT 127.150 3.670 132.290 4.280 ;
        RECT 133.130 3.670 138.270 4.280 ;
        RECT 139.110 3.670 144.250 4.280 ;
        RECT 145.090 3.670 150.230 4.280 ;
        RECT 151.070 3.670 156.210 4.280 ;
        RECT 157.050 3.670 162.190 4.280 ;
        RECT 163.030 3.670 168.170 4.280 ;
        RECT 169.010 3.670 174.150 4.280 ;
        RECT 174.990 3.670 180.130 4.280 ;
        RECT 180.970 3.670 186.110 4.280 ;
        RECT 186.950 3.670 192.090 4.280 ;
        RECT 192.930 3.670 199.940 4.280 ;
      LAYER met3 ;
        RECT 0.065 987.040 196.000 987.525 ;
        RECT 4.400 985.640 196.000 987.040 ;
        RECT 0.065 981.600 196.000 985.640 ;
        RECT 4.400 980.200 196.000 981.600 ;
        RECT 0.065 976.160 196.000 980.200 ;
        RECT 4.400 974.760 196.000 976.160 ;
        RECT 0.065 970.720 196.000 974.760 ;
        RECT 4.400 969.320 196.000 970.720 ;
        RECT 0.065 965.280 196.000 969.320 ;
        RECT 4.400 963.880 196.000 965.280 ;
        RECT 0.065 959.840 196.000 963.880 ;
        RECT 4.400 958.440 196.000 959.840 ;
        RECT 0.065 954.400 196.000 958.440 ;
        RECT 4.400 953.000 196.000 954.400 ;
        RECT 0.065 948.960 196.000 953.000 ;
        RECT 4.400 947.560 196.000 948.960 ;
        RECT 0.065 944.880 196.000 947.560 ;
        RECT 0.065 943.520 195.600 944.880 ;
        RECT 4.400 943.480 195.600 943.520 ;
        RECT 4.400 942.120 196.000 943.480 ;
        RECT 0.065 940.800 196.000 942.120 ;
        RECT 0.065 939.400 195.600 940.800 ;
        RECT 0.065 938.080 196.000 939.400 ;
        RECT 4.400 936.720 196.000 938.080 ;
        RECT 4.400 936.680 195.600 936.720 ;
        RECT 0.065 935.320 195.600 936.680 ;
        RECT 0.065 932.640 196.000 935.320 ;
        RECT 4.400 931.240 195.600 932.640 ;
        RECT 0.065 928.560 196.000 931.240 ;
        RECT 0.065 927.200 195.600 928.560 ;
        RECT 4.400 927.160 195.600 927.200 ;
        RECT 4.400 925.800 196.000 927.160 ;
        RECT 0.065 924.480 196.000 925.800 ;
        RECT 0.065 923.080 195.600 924.480 ;
        RECT 0.065 921.760 196.000 923.080 ;
        RECT 4.400 920.400 196.000 921.760 ;
        RECT 4.400 920.360 195.600 920.400 ;
        RECT 0.065 919.000 195.600 920.360 ;
        RECT 0.065 916.320 196.000 919.000 ;
        RECT 4.400 914.920 195.600 916.320 ;
        RECT 0.065 912.240 196.000 914.920 ;
        RECT 0.065 910.880 195.600 912.240 ;
        RECT 4.400 910.840 195.600 910.880 ;
        RECT 4.400 909.480 196.000 910.840 ;
        RECT 0.065 908.160 196.000 909.480 ;
        RECT 0.065 906.760 195.600 908.160 ;
        RECT 0.065 905.440 196.000 906.760 ;
        RECT 4.400 904.080 196.000 905.440 ;
        RECT 4.400 904.040 195.600 904.080 ;
        RECT 0.065 902.680 195.600 904.040 ;
        RECT 0.065 900.000 196.000 902.680 ;
        RECT 4.400 898.600 195.600 900.000 ;
        RECT 0.065 895.920 196.000 898.600 ;
        RECT 0.065 894.560 195.600 895.920 ;
        RECT 4.400 894.520 195.600 894.560 ;
        RECT 4.400 893.160 196.000 894.520 ;
        RECT 0.065 891.840 196.000 893.160 ;
        RECT 0.065 890.440 195.600 891.840 ;
        RECT 0.065 889.120 196.000 890.440 ;
        RECT 4.400 887.760 196.000 889.120 ;
        RECT 4.400 887.720 195.600 887.760 ;
        RECT 0.065 886.360 195.600 887.720 ;
        RECT 0.065 883.680 196.000 886.360 ;
        RECT 4.400 882.280 195.600 883.680 ;
        RECT 0.065 879.600 196.000 882.280 ;
        RECT 0.065 878.240 195.600 879.600 ;
        RECT 4.400 878.200 195.600 878.240 ;
        RECT 4.400 876.840 196.000 878.200 ;
        RECT 0.065 875.520 196.000 876.840 ;
        RECT 0.065 874.120 195.600 875.520 ;
        RECT 0.065 872.800 196.000 874.120 ;
        RECT 4.400 871.440 196.000 872.800 ;
        RECT 4.400 871.400 195.600 871.440 ;
        RECT 0.065 870.040 195.600 871.400 ;
        RECT 0.065 867.360 196.000 870.040 ;
        RECT 4.400 865.960 195.600 867.360 ;
        RECT 0.065 863.280 196.000 865.960 ;
        RECT 0.065 861.920 195.600 863.280 ;
        RECT 4.400 861.880 195.600 861.920 ;
        RECT 4.400 860.520 196.000 861.880 ;
        RECT 0.065 859.200 196.000 860.520 ;
        RECT 0.065 857.800 195.600 859.200 ;
        RECT 0.065 856.480 196.000 857.800 ;
        RECT 4.400 855.120 196.000 856.480 ;
        RECT 4.400 855.080 195.600 855.120 ;
        RECT 0.065 853.720 195.600 855.080 ;
        RECT 0.065 851.040 196.000 853.720 ;
        RECT 4.400 849.640 195.600 851.040 ;
        RECT 0.065 846.960 196.000 849.640 ;
        RECT 0.065 845.600 195.600 846.960 ;
        RECT 4.400 845.560 195.600 845.600 ;
        RECT 4.400 844.200 196.000 845.560 ;
        RECT 0.065 842.880 196.000 844.200 ;
        RECT 0.065 841.480 195.600 842.880 ;
        RECT 0.065 840.160 196.000 841.480 ;
        RECT 4.400 838.800 196.000 840.160 ;
        RECT 4.400 838.760 195.600 838.800 ;
        RECT 0.065 837.400 195.600 838.760 ;
        RECT 0.065 834.720 196.000 837.400 ;
        RECT 4.400 833.320 195.600 834.720 ;
        RECT 0.065 830.640 196.000 833.320 ;
        RECT 0.065 829.280 195.600 830.640 ;
        RECT 4.400 829.240 195.600 829.280 ;
        RECT 4.400 827.880 196.000 829.240 ;
        RECT 0.065 826.560 196.000 827.880 ;
        RECT 0.065 825.160 195.600 826.560 ;
        RECT 0.065 823.840 196.000 825.160 ;
        RECT 4.400 822.480 196.000 823.840 ;
        RECT 4.400 822.440 195.600 822.480 ;
        RECT 0.065 821.080 195.600 822.440 ;
        RECT 0.065 818.400 196.000 821.080 ;
        RECT 4.400 817.000 195.600 818.400 ;
        RECT 0.065 814.320 196.000 817.000 ;
        RECT 0.065 812.960 195.600 814.320 ;
        RECT 4.400 812.920 195.600 812.960 ;
        RECT 4.400 811.560 196.000 812.920 ;
        RECT 0.065 810.240 196.000 811.560 ;
        RECT 0.065 808.840 195.600 810.240 ;
        RECT 0.065 807.520 196.000 808.840 ;
        RECT 4.400 806.160 196.000 807.520 ;
        RECT 4.400 806.120 195.600 806.160 ;
        RECT 0.065 804.760 195.600 806.120 ;
        RECT 0.065 802.080 196.000 804.760 ;
        RECT 4.400 800.680 195.600 802.080 ;
        RECT 0.065 798.000 196.000 800.680 ;
        RECT 0.065 796.640 195.600 798.000 ;
        RECT 4.400 796.600 195.600 796.640 ;
        RECT 4.400 795.240 196.000 796.600 ;
        RECT 0.065 793.920 196.000 795.240 ;
        RECT 0.065 792.520 195.600 793.920 ;
        RECT 0.065 791.200 196.000 792.520 ;
        RECT 4.400 789.840 196.000 791.200 ;
        RECT 4.400 789.800 195.600 789.840 ;
        RECT 0.065 788.440 195.600 789.800 ;
        RECT 0.065 785.760 196.000 788.440 ;
        RECT 4.400 784.360 195.600 785.760 ;
        RECT 0.065 781.680 196.000 784.360 ;
        RECT 0.065 780.320 195.600 781.680 ;
        RECT 4.400 780.280 195.600 780.320 ;
        RECT 4.400 778.920 196.000 780.280 ;
        RECT 0.065 777.600 196.000 778.920 ;
        RECT 0.065 776.200 195.600 777.600 ;
        RECT 0.065 774.880 196.000 776.200 ;
        RECT 4.400 773.520 196.000 774.880 ;
        RECT 4.400 773.480 195.600 773.520 ;
        RECT 0.065 772.120 195.600 773.480 ;
        RECT 0.065 769.440 196.000 772.120 ;
        RECT 4.400 768.040 195.600 769.440 ;
        RECT 0.065 765.360 196.000 768.040 ;
        RECT 0.065 764.000 195.600 765.360 ;
        RECT 4.400 763.960 195.600 764.000 ;
        RECT 4.400 762.600 196.000 763.960 ;
        RECT 0.065 761.280 196.000 762.600 ;
        RECT 0.065 759.880 195.600 761.280 ;
        RECT 0.065 758.560 196.000 759.880 ;
        RECT 4.400 757.200 196.000 758.560 ;
        RECT 4.400 757.160 195.600 757.200 ;
        RECT 0.065 755.800 195.600 757.160 ;
        RECT 0.065 753.120 196.000 755.800 ;
        RECT 4.400 751.720 195.600 753.120 ;
        RECT 0.065 749.040 196.000 751.720 ;
        RECT 0.065 747.680 195.600 749.040 ;
        RECT 4.400 747.640 195.600 747.680 ;
        RECT 4.400 746.280 196.000 747.640 ;
        RECT 0.065 744.960 196.000 746.280 ;
        RECT 0.065 743.560 195.600 744.960 ;
        RECT 0.065 742.240 196.000 743.560 ;
        RECT 4.400 740.880 196.000 742.240 ;
        RECT 4.400 740.840 195.600 740.880 ;
        RECT 0.065 739.480 195.600 740.840 ;
        RECT 0.065 736.800 196.000 739.480 ;
        RECT 4.400 735.400 195.600 736.800 ;
        RECT 0.065 732.720 196.000 735.400 ;
        RECT 0.065 731.360 195.600 732.720 ;
        RECT 4.400 731.320 195.600 731.360 ;
        RECT 4.400 729.960 196.000 731.320 ;
        RECT 0.065 728.640 196.000 729.960 ;
        RECT 0.065 727.240 195.600 728.640 ;
        RECT 0.065 725.920 196.000 727.240 ;
        RECT 4.400 724.560 196.000 725.920 ;
        RECT 4.400 724.520 195.600 724.560 ;
        RECT 0.065 723.160 195.600 724.520 ;
        RECT 0.065 720.480 196.000 723.160 ;
        RECT 4.400 719.080 195.600 720.480 ;
        RECT 0.065 716.400 196.000 719.080 ;
        RECT 0.065 715.040 195.600 716.400 ;
        RECT 4.400 715.000 195.600 715.040 ;
        RECT 4.400 713.640 196.000 715.000 ;
        RECT 0.065 712.320 196.000 713.640 ;
        RECT 0.065 710.920 195.600 712.320 ;
        RECT 0.065 709.600 196.000 710.920 ;
        RECT 4.400 708.240 196.000 709.600 ;
        RECT 4.400 708.200 195.600 708.240 ;
        RECT 0.065 706.840 195.600 708.200 ;
        RECT 0.065 704.160 196.000 706.840 ;
        RECT 4.400 702.760 195.600 704.160 ;
        RECT 0.065 700.080 196.000 702.760 ;
        RECT 0.065 698.720 195.600 700.080 ;
        RECT 4.400 698.680 195.600 698.720 ;
        RECT 4.400 697.320 196.000 698.680 ;
        RECT 0.065 696.000 196.000 697.320 ;
        RECT 0.065 694.600 195.600 696.000 ;
        RECT 0.065 693.280 196.000 694.600 ;
        RECT 4.400 691.920 196.000 693.280 ;
        RECT 4.400 691.880 195.600 691.920 ;
        RECT 0.065 690.520 195.600 691.880 ;
        RECT 0.065 687.840 196.000 690.520 ;
        RECT 4.400 686.440 195.600 687.840 ;
        RECT 0.065 683.760 196.000 686.440 ;
        RECT 0.065 682.400 195.600 683.760 ;
        RECT 4.400 682.360 195.600 682.400 ;
        RECT 4.400 681.000 196.000 682.360 ;
        RECT 0.065 679.680 196.000 681.000 ;
        RECT 0.065 678.280 195.600 679.680 ;
        RECT 0.065 676.960 196.000 678.280 ;
        RECT 4.400 675.600 196.000 676.960 ;
        RECT 4.400 675.560 195.600 675.600 ;
        RECT 0.065 674.200 195.600 675.560 ;
        RECT 0.065 671.520 196.000 674.200 ;
        RECT 4.400 670.120 195.600 671.520 ;
        RECT 0.065 667.440 196.000 670.120 ;
        RECT 0.065 666.080 195.600 667.440 ;
        RECT 4.400 666.040 195.600 666.080 ;
        RECT 4.400 664.680 196.000 666.040 ;
        RECT 0.065 663.360 196.000 664.680 ;
        RECT 0.065 661.960 195.600 663.360 ;
        RECT 0.065 660.640 196.000 661.960 ;
        RECT 4.400 659.280 196.000 660.640 ;
        RECT 4.400 659.240 195.600 659.280 ;
        RECT 0.065 657.880 195.600 659.240 ;
        RECT 0.065 655.200 196.000 657.880 ;
        RECT 4.400 653.800 195.600 655.200 ;
        RECT 0.065 651.120 196.000 653.800 ;
        RECT 0.065 649.760 195.600 651.120 ;
        RECT 4.400 649.720 195.600 649.760 ;
        RECT 4.400 648.360 196.000 649.720 ;
        RECT 0.065 647.040 196.000 648.360 ;
        RECT 0.065 645.640 195.600 647.040 ;
        RECT 0.065 644.320 196.000 645.640 ;
        RECT 4.400 642.960 196.000 644.320 ;
        RECT 4.400 642.920 195.600 642.960 ;
        RECT 0.065 641.560 195.600 642.920 ;
        RECT 0.065 638.880 196.000 641.560 ;
        RECT 4.400 637.480 195.600 638.880 ;
        RECT 0.065 634.800 196.000 637.480 ;
        RECT 0.065 633.440 195.600 634.800 ;
        RECT 4.400 633.400 195.600 633.440 ;
        RECT 4.400 632.040 196.000 633.400 ;
        RECT 0.065 630.720 196.000 632.040 ;
        RECT 0.065 629.320 195.600 630.720 ;
        RECT 0.065 628.000 196.000 629.320 ;
        RECT 4.400 626.640 196.000 628.000 ;
        RECT 4.400 626.600 195.600 626.640 ;
        RECT 0.065 625.240 195.600 626.600 ;
        RECT 0.065 622.560 196.000 625.240 ;
        RECT 4.400 621.160 195.600 622.560 ;
        RECT 0.065 618.480 196.000 621.160 ;
        RECT 0.065 617.120 195.600 618.480 ;
        RECT 4.400 617.080 195.600 617.120 ;
        RECT 4.400 615.720 196.000 617.080 ;
        RECT 0.065 614.400 196.000 615.720 ;
        RECT 0.065 613.000 195.600 614.400 ;
        RECT 0.065 611.680 196.000 613.000 ;
        RECT 4.400 610.320 196.000 611.680 ;
        RECT 4.400 610.280 195.600 610.320 ;
        RECT 0.065 608.920 195.600 610.280 ;
        RECT 0.065 606.240 196.000 608.920 ;
        RECT 4.400 604.840 195.600 606.240 ;
        RECT 0.065 602.160 196.000 604.840 ;
        RECT 0.065 600.800 195.600 602.160 ;
        RECT 4.400 600.760 195.600 600.800 ;
        RECT 4.400 599.400 196.000 600.760 ;
        RECT 0.065 598.080 196.000 599.400 ;
        RECT 0.065 596.680 195.600 598.080 ;
        RECT 0.065 595.360 196.000 596.680 ;
        RECT 4.400 594.000 196.000 595.360 ;
        RECT 4.400 593.960 195.600 594.000 ;
        RECT 0.065 592.600 195.600 593.960 ;
        RECT 0.065 589.920 196.000 592.600 ;
        RECT 4.400 588.520 195.600 589.920 ;
        RECT 0.065 585.840 196.000 588.520 ;
        RECT 0.065 584.480 195.600 585.840 ;
        RECT 4.400 584.440 195.600 584.480 ;
        RECT 4.400 583.080 196.000 584.440 ;
        RECT 0.065 581.760 196.000 583.080 ;
        RECT 0.065 580.360 195.600 581.760 ;
        RECT 0.065 579.040 196.000 580.360 ;
        RECT 4.400 577.680 196.000 579.040 ;
        RECT 4.400 577.640 195.600 577.680 ;
        RECT 0.065 576.280 195.600 577.640 ;
        RECT 0.065 573.600 196.000 576.280 ;
        RECT 4.400 572.200 195.600 573.600 ;
        RECT 0.065 569.520 196.000 572.200 ;
        RECT 0.065 568.160 195.600 569.520 ;
        RECT 4.400 568.120 195.600 568.160 ;
        RECT 4.400 566.760 196.000 568.120 ;
        RECT 0.065 565.440 196.000 566.760 ;
        RECT 0.065 564.040 195.600 565.440 ;
        RECT 0.065 562.720 196.000 564.040 ;
        RECT 4.400 561.360 196.000 562.720 ;
        RECT 4.400 561.320 195.600 561.360 ;
        RECT 0.065 559.960 195.600 561.320 ;
        RECT 0.065 557.280 196.000 559.960 ;
        RECT 4.400 555.880 195.600 557.280 ;
        RECT 0.065 553.200 196.000 555.880 ;
        RECT 0.065 551.840 195.600 553.200 ;
        RECT 4.400 551.800 195.600 551.840 ;
        RECT 4.400 550.440 196.000 551.800 ;
        RECT 0.065 549.120 196.000 550.440 ;
        RECT 0.065 547.720 195.600 549.120 ;
        RECT 0.065 546.400 196.000 547.720 ;
        RECT 4.400 545.040 196.000 546.400 ;
        RECT 4.400 545.000 195.600 545.040 ;
        RECT 0.065 543.640 195.600 545.000 ;
        RECT 0.065 540.960 196.000 543.640 ;
        RECT 4.400 539.560 195.600 540.960 ;
        RECT 0.065 536.880 196.000 539.560 ;
        RECT 0.065 535.520 195.600 536.880 ;
        RECT 4.400 535.480 195.600 535.520 ;
        RECT 4.400 534.120 196.000 535.480 ;
        RECT 0.065 532.800 196.000 534.120 ;
        RECT 0.065 531.400 195.600 532.800 ;
        RECT 0.065 530.080 196.000 531.400 ;
        RECT 4.400 528.720 196.000 530.080 ;
        RECT 4.400 528.680 195.600 528.720 ;
        RECT 0.065 527.320 195.600 528.680 ;
        RECT 0.065 524.640 196.000 527.320 ;
        RECT 4.400 523.240 195.600 524.640 ;
        RECT 0.065 520.560 196.000 523.240 ;
        RECT 0.065 519.200 195.600 520.560 ;
        RECT 4.400 519.160 195.600 519.200 ;
        RECT 4.400 517.800 196.000 519.160 ;
        RECT 0.065 516.480 196.000 517.800 ;
        RECT 0.065 515.080 195.600 516.480 ;
        RECT 0.065 513.760 196.000 515.080 ;
        RECT 4.400 512.400 196.000 513.760 ;
        RECT 4.400 512.360 195.600 512.400 ;
        RECT 0.065 511.000 195.600 512.360 ;
        RECT 0.065 508.320 196.000 511.000 ;
        RECT 4.400 506.920 195.600 508.320 ;
        RECT 0.065 504.240 196.000 506.920 ;
        RECT 0.065 502.880 195.600 504.240 ;
        RECT 4.400 502.840 195.600 502.880 ;
        RECT 4.400 501.480 196.000 502.840 ;
        RECT 0.065 500.160 196.000 501.480 ;
        RECT 0.065 498.760 195.600 500.160 ;
        RECT 0.065 497.440 196.000 498.760 ;
        RECT 4.400 496.080 196.000 497.440 ;
        RECT 4.400 496.040 195.600 496.080 ;
        RECT 0.065 494.680 195.600 496.040 ;
        RECT 0.065 492.000 196.000 494.680 ;
        RECT 4.400 490.600 195.600 492.000 ;
        RECT 0.065 487.920 196.000 490.600 ;
        RECT 0.065 486.560 195.600 487.920 ;
        RECT 4.400 486.520 195.600 486.560 ;
        RECT 4.400 485.160 196.000 486.520 ;
        RECT 0.065 483.840 196.000 485.160 ;
        RECT 0.065 482.440 195.600 483.840 ;
        RECT 0.065 481.120 196.000 482.440 ;
        RECT 4.400 479.760 196.000 481.120 ;
        RECT 4.400 479.720 195.600 479.760 ;
        RECT 0.065 478.360 195.600 479.720 ;
        RECT 0.065 475.680 196.000 478.360 ;
        RECT 4.400 474.280 195.600 475.680 ;
        RECT 0.065 471.600 196.000 474.280 ;
        RECT 0.065 470.240 195.600 471.600 ;
        RECT 4.400 470.200 195.600 470.240 ;
        RECT 4.400 468.840 196.000 470.200 ;
        RECT 0.065 467.520 196.000 468.840 ;
        RECT 0.065 466.120 195.600 467.520 ;
        RECT 0.065 464.800 196.000 466.120 ;
        RECT 4.400 463.440 196.000 464.800 ;
        RECT 4.400 463.400 195.600 463.440 ;
        RECT 0.065 462.040 195.600 463.400 ;
        RECT 0.065 459.360 196.000 462.040 ;
        RECT 4.400 457.960 195.600 459.360 ;
        RECT 0.065 455.280 196.000 457.960 ;
        RECT 0.065 453.920 195.600 455.280 ;
        RECT 4.400 453.880 195.600 453.920 ;
        RECT 4.400 452.520 196.000 453.880 ;
        RECT 0.065 451.200 196.000 452.520 ;
        RECT 0.065 449.800 195.600 451.200 ;
        RECT 0.065 448.480 196.000 449.800 ;
        RECT 4.400 447.120 196.000 448.480 ;
        RECT 4.400 447.080 195.600 447.120 ;
        RECT 0.065 445.720 195.600 447.080 ;
        RECT 0.065 443.040 196.000 445.720 ;
        RECT 4.400 441.640 195.600 443.040 ;
        RECT 0.065 438.960 196.000 441.640 ;
        RECT 0.065 437.600 195.600 438.960 ;
        RECT 4.400 437.560 195.600 437.600 ;
        RECT 4.400 436.200 196.000 437.560 ;
        RECT 0.065 434.880 196.000 436.200 ;
        RECT 0.065 433.480 195.600 434.880 ;
        RECT 0.065 432.160 196.000 433.480 ;
        RECT 4.400 430.800 196.000 432.160 ;
        RECT 4.400 430.760 195.600 430.800 ;
        RECT 0.065 429.400 195.600 430.760 ;
        RECT 0.065 426.720 196.000 429.400 ;
        RECT 4.400 425.320 195.600 426.720 ;
        RECT 0.065 422.640 196.000 425.320 ;
        RECT 0.065 421.280 195.600 422.640 ;
        RECT 4.400 421.240 195.600 421.280 ;
        RECT 4.400 419.880 196.000 421.240 ;
        RECT 0.065 418.560 196.000 419.880 ;
        RECT 0.065 417.160 195.600 418.560 ;
        RECT 0.065 415.840 196.000 417.160 ;
        RECT 4.400 414.480 196.000 415.840 ;
        RECT 4.400 414.440 195.600 414.480 ;
        RECT 0.065 413.080 195.600 414.440 ;
        RECT 0.065 410.400 196.000 413.080 ;
        RECT 4.400 409.000 195.600 410.400 ;
        RECT 0.065 406.320 196.000 409.000 ;
        RECT 0.065 404.960 195.600 406.320 ;
        RECT 4.400 404.920 195.600 404.960 ;
        RECT 4.400 403.560 196.000 404.920 ;
        RECT 0.065 402.240 196.000 403.560 ;
        RECT 0.065 400.840 195.600 402.240 ;
        RECT 0.065 399.520 196.000 400.840 ;
        RECT 4.400 398.160 196.000 399.520 ;
        RECT 4.400 398.120 195.600 398.160 ;
        RECT 0.065 396.760 195.600 398.120 ;
        RECT 0.065 394.080 196.000 396.760 ;
        RECT 4.400 392.680 195.600 394.080 ;
        RECT 0.065 390.000 196.000 392.680 ;
        RECT 0.065 388.640 195.600 390.000 ;
        RECT 4.400 388.600 195.600 388.640 ;
        RECT 4.400 387.240 196.000 388.600 ;
        RECT 0.065 385.920 196.000 387.240 ;
        RECT 0.065 384.520 195.600 385.920 ;
        RECT 0.065 383.200 196.000 384.520 ;
        RECT 4.400 381.840 196.000 383.200 ;
        RECT 4.400 381.800 195.600 381.840 ;
        RECT 0.065 380.440 195.600 381.800 ;
        RECT 0.065 377.760 196.000 380.440 ;
        RECT 4.400 376.360 195.600 377.760 ;
        RECT 0.065 373.680 196.000 376.360 ;
        RECT 0.065 372.320 195.600 373.680 ;
        RECT 4.400 372.280 195.600 372.320 ;
        RECT 4.400 370.920 196.000 372.280 ;
        RECT 0.065 369.600 196.000 370.920 ;
        RECT 0.065 368.200 195.600 369.600 ;
        RECT 0.065 366.880 196.000 368.200 ;
        RECT 4.400 365.520 196.000 366.880 ;
        RECT 4.400 365.480 195.600 365.520 ;
        RECT 0.065 364.120 195.600 365.480 ;
        RECT 0.065 361.440 196.000 364.120 ;
        RECT 4.400 360.040 195.600 361.440 ;
        RECT 0.065 357.360 196.000 360.040 ;
        RECT 0.065 356.000 195.600 357.360 ;
        RECT 4.400 355.960 195.600 356.000 ;
        RECT 4.400 354.600 196.000 355.960 ;
        RECT 0.065 353.280 196.000 354.600 ;
        RECT 0.065 351.880 195.600 353.280 ;
        RECT 0.065 350.560 196.000 351.880 ;
        RECT 4.400 349.200 196.000 350.560 ;
        RECT 4.400 349.160 195.600 349.200 ;
        RECT 0.065 347.800 195.600 349.160 ;
        RECT 0.065 345.120 196.000 347.800 ;
        RECT 4.400 343.720 195.600 345.120 ;
        RECT 0.065 341.040 196.000 343.720 ;
        RECT 0.065 339.680 195.600 341.040 ;
        RECT 4.400 339.640 195.600 339.680 ;
        RECT 4.400 338.280 196.000 339.640 ;
        RECT 0.065 336.960 196.000 338.280 ;
        RECT 0.065 335.560 195.600 336.960 ;
        RECT 0.065 334.240 196.000 335.560 ;
        RECT 4.400 332.880 196.000 334.240 ;
        RECT 4.400 332.840 195.600 332.880 ;
        RECT 0.065 331.480 195.600 332.840 ;
        RECT 0.065 328.800 196.000 331.480 ;
        RECT 4.400 327.400 195.600 328.800 ;
        RECT 0.065 324.720 196.000 327.400 ;
        RECT 0.065 323.360 195.600 324.720 ;
        RECT 4.400 323.320 195.600 323.360 ;
        RECT 4.400 321.960 196.000 323.320 ;
        RECT 0.065 320.640 196.000 321.960 ;
        RECT 0.065 319.240 195.600 320.640 ;
        RECT 0.065 317.920 196.000 319.240 ;
        RECT 4.400 316.560 196.000 317.920 ;
        RECT 4.400 316.520 195.600 316.560 ;
        RECT 0.065 315.160 195.600 316.520 ;
        RECT 0.065 312.480 196.000 315.160 ;
        RECT 4.400 311.080 195.600 312.480 ;
        RECT 0.065 308.400 196.000 311.080 ;
        RECT 0.065 307.040 195.600 308.400 ;
        RECT 4.400 307.000 195.600 307.040 ;
        RECT 4.400 305.640 196.000 307.000 ;
        RECT 0.065 304.320 196.000 305.640 ;
        RECT 0.065 302.920 195.600 304.320 ;
        RECT 0.065 301.600 196.000 302.920 ;
        RECT 4.400 300.240 196.000 301.600 ;
        RECT 4.400 300.200 195.600 300.240 ;
        RECT 0.065 298.840 195.600 300.200 ;
        RECT 0.065 296.160 196.000 298.840 ;
        RECT 4.400 294.760 195.600 296.160 ;
        RECT 0.065 292.080 196.000 294.760 ;
        RECT 0.065 290.720 195.600 292.080 ;
        RECT 4.400 290.680 195.600 290.720 ;
        RECT 4.400 289.320 196.000 290.680 ;
        RECT 0.065 288.000 196.000 289.320 ;
        RECT 0.065 286.600 195.600 288.000 ;
        RECT 0.065 285.280 196.000 286.600 ;
        RECT 4.400 283.920 196.000 285.280 ;
        RECT 4.400 283.880 195.600 283.920 ;
        RECT 0.065 282.520 195.600 283.880 ;
        RECT 0.065 279.840 196.000 282.520 ;
        RECT 4.400 278.440 195.600 279.840 ;
        RECT 0.065 275.760 196.000 278.440 ;
        RECT 0.065 274.400 195.600 275.760 ;
        RECT 4.400 274.360 195.600 274.400 ;
        RECT 4.400 273.000 196.000 274.360 ;
        RECT 0.065 271.680 196.000 273.000 ;
        RECT 0.065 270.280 195.600 271.680 ;
        RECT 0.065 268.960 196.000 270.280 ;
        RECT 4.400 267.600 196.000 268.960 ;
        RECT 4.400 267.560 195.600 267.600 ;
        RECT 0.065 266.200 195.600 267.560 ;
        RECT 0.065 263.520 196.000 266.200 ;
        RECT 4.400 262.120 195.600 263.520 ;
        RECT 0.065 259.440 196.000 262.120 ;
        RECT 0.065 258.080 195.600 259.440 ;
        RECT 4.400 258.040 195.600 258.080 ;
        RECT 4.400 256.680 196.000 258.040 ;
        RECT 0.065 255.360 196.000 256.680 ;
        RECT 0.065 253.960 195.600 255.360 ;
        RECT 0.065 252.640 196.000 253.960 ;
        RECT 4.400 251.280 196.000 252.640 ;
        RECT 4.400 251.240 195.600 251.280 ;
        RECT 0.065 249.880 195.600 251.240 ;
        RECT 0.065 247.200 196.000 249.880 ;
        RECT 4.400 245.800 195.600 247.200 ;
        RECT 0.065 243.120 196.000 245.800 ;
        RECT 0.065 241.760 195.600 243.120 ;
        RECT 4.400 241.720 195.600 241.760 ;
        RECT 4.400 240.360 196.000 241.720 ;
        RECT 0.065 239.040 196.000 240.360 ;
        RECT 0.065 237.640 195.600 239.040 ;
        RECT 0.065 236.320 196.000 237.640 ;
        RECT 4.400 234.960 196.000 236.320 ;
        RECT 4.400 234.920 195.600 234.960 ;
        RECT 0.065 233.560 195.600 234.920 ;
        RECT 0.065 230.880 196.000 233.560 ;
        RECT 4.400 229.480 195.600 230.880 ;
        RECT 0.065 226.800 196.000 229.480 ;
        RECT 0.065 225.440 195.600 226.800 ;
        RECT 4.400 225.400 195.600 225.440 ;
        RECT 4.400 224.040 196.000 225.400 ;
        RECT 0.065 222.720 196.000 224.040 ;
        RECT 0.065 221.320 195.600 222.720 ;
        RECT 0.065 220.000 196.000 221.320 ;
        RECT 4.400 218.640 196.000 220.000 ;
        RECT 4.400 218.600 195.600 218.640 ;
        RECT 0.065 217.240 195.600 218.600 ;
        RECT 0.065 214.560 196.000 217.240 ;
        RECT 4.400 213.160 195.600 214.560 ;
        RECT 0.065 210.480 196.000 213.160 ;
        RECT 0.065 209.120 195.600 210.480 ;
        RECT 4.400 209.080 195.600 209.120 ;
        RECT 4.400 207.720 196.000 209.080 ;
        RECT 0.065 206.400 196.000 207.720 ;
        RECT 0.065 205.000 195.600 206.400 ;
        RECT 0.065 203.680 196.000 205.000 ;
        RECT 4.400 202.320 196.000 203.680 ;
        RECT 4.400 202.280 195.600 202.320 ;
        RECT 0.065 200.920 195.600 202.280 ;
        RECT 0.065 198.240 196.000 200.920 ;
        RECT 4.400 196.840 195.600 198.240 ;
        RECT 0.065 194.160 196.000 196.840 ;
        RECT 0.065 192.800 195.600 194.160 ;
        RECT 4.400 192.760 195.600 192.800 ;
        RECT 4.400 191.400 196.000 192.760 ;
        RECT 0.065 190.080 196.000 191.400 ;
        RECT 0.065 188.680 195.600 190.080 ;
        RECT 0.065 187.360 196.000 188.680 ;
        RECT 4.400 186.000 196.000 187.360 ;
        RECT 4.400 185.960 195.600 186.000 ;
        RECT 0.065 184.600 195.600 185.960 ;
        RECT 0.065 181.920 196.000 184.600 ;
        RECT 4.400 180.520 195.600 181.920 ;
        RECT 0.065 177.840 196.000 180.520 ;
        RECT 0.065 176.480 195.600 177.840 ;
        RECT 4.400 176.440 195.600 176.480 ;
        RECT 4.400 175.080 196.000 176.440 ;
        RECT 0.065 173.760 196.000 175.080 ;
        RECT 0.065 172.360 195.600 173.760 ;
        RECT 0.065 171.040 196.000 172.360 ;
        RECT 4.400 169.680 196.000 171.040 ;
        RECT 4.400 169.640 195.600 169.680 ;
        RECT 0.065 168.280 195.600 169.640 ;
        RECT 0.065 165.600 196.000 168.280 ;
        RECT 4.400 164.200 195.600 165.600 ;
        RECT 0.065 161.520 196.000 164.200 ;
        RECT 0.065 160.160 195.600 161.520 ;
        RECT 4.400 160.120 195.600 160.160 ;
        RECT 4.400 158.760 196.000 160.120 ;
        RECT 0.065 157.440 196.000 158.760 ;
        RECT 0.065 156.040 195.600 157.440 ;
        RECT 0.065 154.720 196.000 156.040 ;
        RECT 4.400 153.360 196.000 154.720 ;
        RECT 4.400 153.320 195.600 153.360 ;
        RECT 0.065 151.960 195.600 153.320 ;
        RECT 0.065 149.280 196.000 151.960 ;
        RECT 4.400 147.880 195.600 149.280 ;
        RECT 0.065 145.200 196.000 147.880 ;
        RECT 0.065 143.840 195.600 145.200 ;
        RECT 4.400 143.800 195.600 143.840 ;
        RECT 4.400 142.440 196.000 143.800 ;
        RECT 0.065 141.120 196.000 142.440 ;
        RECT 0.065 139.720 195.600 141.120 ;
        RECT 0.065 138.400 196.000 139.720 ;
        RECT 4.400 137.040 196.000 138.400 ;
        RECT 4.400 137.000 195.600 137.040 ;
        RECT 0.065 135.640 195.600 137.000 ;
        RECT 0.065 132.960 196.000 135.640 ;
        RECT 4.400 131.560 195.600 132.960 ;
        RECT 0.065 128.880 196.000 131.560 ;
        RECT 0.065 127.520 195.600 128.880 ;
        RECT 4.400 127.480 195.600 127.520 ;
        RECT 4.400 126.120 196.000 127.480 ;
        RECT 0.065 124.800 196.000 126.120 ;
        RECT 0.065 123.400 195.600 124.800 ;
        RECT 0.065 122.080 196.000 123.400 ;
        RECT 4.400 120.720 196.000 122.080 ;
        RECT 4.400 120.680 195.600 120.720 ;
        RECT 0.065 119.320 195.600 120.680 ;
        RECT 0.065 116.640 196.000 119.320 ;
        RECT 4.400 115.240 195.600 116.640 ;
        RECT 0.065 112.560 196.000 115.240 ;
        RECT 0.065 111.200 195.600 112.560 ;
        RECT 4.400 111.160 195.600 111.200 ;
        RECT 4.400 109.800 196.000 111.160 ;
        RECT 0.065 108.480 196.000 109.800 ;
        RECT 0.065 107.080 195.600 108.480 ;
        RECT 0.065 105.760 196.000 107.080 ;
        RECT 4.400 104.400 196.000 105.760 ;
        RECT 4.400 104.360 195.600 104.400 ;
        RECT 0.065 103.000 195.600 104.360 ;
        RECT 0.065 100.320 196.000 103.000 ;
        RECT 4.400 98.920 195.600 100.320 ;
        RECT 0.065 96.240 196.000 98.920 ;
        RECT 0.065 94.880 195.600 96.240 ;
        RECT 4.400 94.840 195.600 94.880 ;
        RECT 4.400 93.480 196.000 94.840 ;
        RECT 0.065 92.160 196.000 93.480 ;
        RECT 0.065 90.760 195.600 92.160 ;
        RECT 0.065 89.440 196.000 90.760 ;
        RECT 4.400 88.080 196.000 89.440 ;
        RECT 4.400 88.040 195.600 88.080 ;
        RECT 0.065 86.680 195.600 88.040 ;
        RECT 0.065 84.000 196.000 86.680 ;
        RECT 4.400 82.600 195.600 84.000 ;
        RECT 0.065 79.920 196.000 82.600 ;
        RECT 0.065 78.560 195.600 79.920 ;
        RECT 4.400 78.520 195.600 78.560 ;
        RECT 4.400 77.160 196.000 78.520 ;
        RECT 0.065 75.840 196.000 77.160 ;
        RECT 0.065 74.440 195.600 75.840 ;
        RECT 0.065 73.120 196.000 74.440 ;
        RECT 4.400 71.760 196.000 73.120 ;
        RECT 4.400 71.720 195.600 71.760 ;
        RECT 0.065 70.360 195.600 71.720 ;
        RECT 0.065 67.680 196.000 70.360 ;
        RECT 4.400 66.280 195.600 67.680 ;
        RECT 0.065 63.600 196.000 66.280 ;
        RECT 0.065 62.240 195.600 63.600 ;
        RECT 4.400 62.200 195.600 62.240 ;
        RECT 4.400 60.840 196.000 62.200 ;
        RECT 0.065 59.520 196.000 60.840 ;
        RECT 0.065 58.120 195.600 59.520 ;
        RECT 0.065 56.800 196.000 58.120 ;
        RECT 4.400 55.440 196.000 56.800 ;
        RECT 4.400 55.400 195.600 55.440 ;
        RECT 0.065 54.040 195.600 55.400 ;
        RECT 0.065 51.360 196.000 54.040 ;
        RECT 4.400 49.960 196.000 51.360 ;
        RECT 0.065 45.920 196.000 49.960 ;
        RECT 4.400 44.520 196.000 45.920 ;
        RECT 0.065 40.480 196.000 44.520 ;
        RECT 4.400 39.080 196.000 40.480 ;
        RECT 0.065 35.040 196.000 39.080 ;
        RECT 4.400 33.640 196.000 35.040 ;
        RECT 0.065 29.600 196.000 33.640 ;
        RECT 4.400 28.200 196.000 29.600 ;
        RECT 0.065 24.160 196.000 28.200 ;
        RECT 4.400 22.760 196.000 24.160 ;
        RECT 0.065 18.720 196.000 22.760 ;
        RECT 4.400 17.320 196.000 18.720 ;
        RECT 0.065 13.280 196.000 17.320 ;
        RECT 4.400 11.880 196.000 13.280 ;
        RECT 0.065 10.715 196.000 11.880 ;
      LAYER met4 ;
        RECT 3.055 15.135 20.640 883.825 ;
        RECT 23.040 15.135 97.440 883.825 ;
        RECT 99.840 15.135 174.240 883.825 ;
        RECT 176.640 15.135 185.545 883.825 ;
  END
END multiplexer
END LIBRARY

