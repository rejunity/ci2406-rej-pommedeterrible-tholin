magic
tech sky130A
magscale 1 2
timestamp 1716584809
<< obsli1 >>
rect 1104 2159 78844 97393
<< obsm1 >>
rect 14 2128 79106 97424
<< metal2 >>
rect 1490 99200 1546 100000
rect 3514 99200 3570 100000
rect 5538 99200 5594 100000
rect 7562 99200 7618 100000
rect 9586 99200 9642 100000
rect 11610 99200 11666 100000
rect 13634 99200 13690 100000
rect 15658 99200 15714 100000
rect 17682 99200 17738 100000
rect 19706 99200 19762 100000
rect 21730 99200 21786 100000
rect 23754 99200 23810 100000
rect 25778 99200 25834 100000
rect 27802 99200 27858 100000
rect 29826 99200 29882 100000
rect 31850 99200 31906 100000
rect 33874 99200 33930 100000
rect 35898 99200 35954 100000
rect 37922 99200 37978 100000
rect 39946 99200 40002 100000
rect 41970 99200 42026 100000
rect 43994 99200 44050 100000
rect 46018 99200 46074 100000
rect 48042 99200 48098 100000
rect 50066 99200 50122 100000
rect 52090 99200 52146 100000
rect 54114 99200 54170 100000
rect 56138 99200 56194 100000
rect 58162 99200 58218 100000
rect 60186 99200 60242 100000
rect 62210 99200 62266 100000
rect 64234 99200 64290 100000
rect 66258 99200 66314 100000
rect 68282 99200 68338 100000
rect 70306 99200 70362 100000
rect 72330 99200 72386 100000
rect 74354 99200 74410 100000
rect 76378 99200 76434 100000
rect 78402 99200 78458 100000
rect 1030 0 1086 800
rect 2226 0 2282 800
rect 3422 0 3478 800
rect 4618 0 4674 800
rect 5814 0 5870 800
rect 7010 0 7066 800
rect 8206 0 8262 800
rect 9402 0 9458 800
rect 10598 0 10654 800
rect 11794 0 11850 800
rect 12990 0 13046 800
rect 14186 0 14242 800
rect 15382 0 15438 800
rect 16578 0 16634 800
rect 17774 0 17830 800
rect 18970 0 19026 800
rect 20166 0 20222 800
rect 21362 0 21418 800
rect 22558 0 22614 800
rect 23754 0 23810 800
rect 24950 0 25006 800
rect 26146 0 26202 800
rect 27342 0 27398 800
rect 28538 0 28594 800
rect 29734 0 29790 800
rect 30930 0 30986 800
rect 32126 0 32182 800
rect 33322 0 33378 800
rect 34518 0 34574 800
rect 35714 0 35770 800
rect 36910 0 36966 800
rect 38106 0 38162 800
rect 39302 0 39358 800
rect 40498 0 40554 800
rect 41694 0 41750 800
rect 42890 0 42946 800
rect 44086 0 44142 800
rect 45282 0 45338 800
rect 46478 0 46534 800
rect 47674 0 47730 800
rect 48870 0 48926 800
rect 50066 0 50122 800
rect 51262 0 51318 800
rect 52458 0 52514 800
rect 53654 0 53710 800
rect 54850 0 54906 800
rect 56046 0 56102 800
rect 57242 0 57298 800
rect 58438 0 58494 800
rect 59634 0 59690 800
rect 60830 0 60886 800
rect 62026 0 62082 800
rect 63222 0 63278 800
rect 64418 0 64474 800
rect 65614 0 65670 800
rect 66810 0 66866 800
rect 68006 0 68062 800
rect 69202 0 69258 800
rect 70398 0 70454 800
rect 71594 0 71650 800
rect 72790 0 72846 800
rect 73986 0 74042 800
rect 75182 0 75238 800
rect 76378 0 76434 800
rect 77574 0 77630 800
rect 78770 0 78826 800
<< obsm2 >>
rect 20 99144 1434 99362
rect 1602 99144 3458 99362
rect 3626 99144 5482 99362
rect 5650 99144 7506 99362
rect 7674 99144 9530 99362
rect 9698 99144 11554 99362
rect 11722 99144 13578 99362
rect 13746 99144 15602 99362
rect 15770 99144 17626 99362
rect 17794 99144 19650 99362
rect 19818 99144 21674 99362
rect 21842 99144 23698 99362
rect 23866 99144 25722 99362
rect 25890 99144 27746 99362
rect 27914 99144 29770 99362
rect 29938 99144 31794 99362
rect 31962 99144 33818 99362
rect 33986 99144 35842 99362
rect 36010 99144 37866 99362
rect 38034 99144 39890 99362
rect 40058 99144 41914 99362
rect 42082 99144 43938 99362
rect 44106 99144 45962 99362
rect 46130 99144 47986 99362
rect 48154 99144 50010 99362
rect 50178 99144 52034 99362
rect 52202 99144 54058 99362
rect 54226 99144 56082 99362
rect 56250 99144 58106 99362
rect 58274 99144 60130 99362
rect 60298 99144 62154 99362
rect 62322 99144 64178 99362
rect 64346 99144 66202 99362
rect 66370 99144 68226 99362
rect 68394 99144 70250 99362
rect 70418 99144 72274 99362
rect 72442 99144 74298 99362
rect 74466 99144 76322 99362
rect 76490 99144 78346 99362
rect 78514 99144 79102 99362
rect 20 856 79102 99144
rect 20 734 974 856
rect 1142 734 2170 856
rect 2338 734 3366 856
rect 3534 734 4562 856
rect 4730 734 5758 856
rect 5926 734 6954 856
rect 7122 734 8150 856
rect 8318 734 9346 856
rect 9514 734 10542 856
rect 10710 734 11738 856
rect 11906 734 12934 856
rect 13102 734 14130 856
rect 14298 734 15326 856
rect 15494 734 16522 856
rect 16690 734 17718 856
rect 17886 734 18914 856
rect 19082 734 20110 856
rect 20278 734 21306 856
rect 21474 734 22502 856
rect 22670 734 23698 856
rect 23866 734 24894 856
rect 25062 734 26090 856
rect 26258 734 27286 856
rect 27454 734 28482 856
rect 28650 734 29678 856
rect 29846 734 30874 856
rect 31042 734 32070 856
rect 32238 734 33266 856
rect 33434 734 34462 856
rect 34630 734 35658 856
rect 35826 734 36854 856
rect 37022 734 38050 856
rect 38218 734 39246 856
rect 39414 734 40442 856
rect 40610 734 41638 856
rect 41806 734 42834 856
rect 43002 734 44030 856
rect 44198 734 45226 856
rect 45394 734 46422 856
rect 46590 734 47618 856
rect 47786 734 48814 856
rect 48982 734 50010 856
rect 50178 734 51206 856
rect 51374 734 52402 856
rect 52570 734 53598 856
rect 53766 734 54794 856
rect 54962 734 55990 856
rect 56158 734 57186 856
rect 57354 734 58382 856
rect 58550 734 59578 856
rect 59746 734 60774 856
rect 60942 734 61970 856
rect 62138 734 63166 856
rect 63334 734 64362 856
rect 64530 734 65558 856
rect 65726 734 66754 856
rect 66922 734 67950 856
rect 68118 734 69146 856
rect 69314 734 70342 856
rect 70510 734 71538 856
rect 71706 734 72734 856
rect 72902 734 73930 856
rect 74098 734 75126 856
rect 75294 734 76322 856
rect 76490 734 77518 856
rect 77686 734 78714 856
rect 78882 734 79102 856
<< metal3 >>
rect 0 94664 800 94784
rect 0 93848 800 93968
rect 79200 93576 80000 93696
rect 0 93032 800 93152
rect 79200 92760 80000 92880
rect 0 92216 800 92336
rect 79200 91944 80000 92064
rect 0 91400 800 91520
rect 79200 91128 80000 91248
rect 0 90584 800 90704
rect 79200 90312 80000 90432
rect 0 89768 800 89888
rect 79200 89496 80000 89616
rect 0 88952 800 89072
rect 79200 88680 80000 88800
rect 0 88136 800 88256
rect 79200 87864 80000 87984
rect 0 87320 800 87440
rect 79200 87048 80000 87168
rect 0 86504 800 86624
rect 79200 86232 80000 86352
rect 0 85688 800 85808
rect 79200 85416 80000 85536
rect 0 84872 800 84992
rect 79200 84600 80000 84720
rect 0 84056 800 84176
rect 79200 83784 80000 83904
rect 0 83240 800 83360
rect 79200 82968 80000 83088
rect 0 82424 800 82544
rect 79200 82152 80000 82272
rect 0 81608 800 81728
rect 79200 81336 80000 81456
rect 0 80792 800 80912
rect 79200 80520 80000 80640
rect 0 79976 800 80096
rect 79200 79704 80000 79824
rect 0 79160 800 79280
rect 79200 78888 80000 79008
rect 0 78344 800 78464
rect 79200 78072 80000 78192
rect 0 77528 800 77648
rect 79200 77256 80000 77376
rect 0 76712 800 76832
rect 79200 76440 80000 76560
rect 0 75896 800 76016
rect 79200 75624 80000 75744
rect 0 75080 800 75200
rect 79200 74808 80000 74928
rect 0 74264 800 74384
rect 79200 73992 80000 74112
rect 0 73448 800 73568
rect 79200 73176 80000 73296
rect 0 72632 800 72752
rect 79200 72360 80000 72480
rect 0 71816 800 71936
rect 79200 71544 80000 71664
rect 0 71000 800 71120
rect 79200 70728 80000 70848
rect 0 70184 800 70304
rect 79200 69912 80000 70032
rect 0 69368 800 69488
rect 79200 69096 80000 69216
rect 0 68552 800 68672
rect 79200 68280 80000 68400
rect 0 67736 800 67856
rect 79200 67464 80000 67584
rect 0 66920 800 67040
rect 79200 66648 80000 66768
rect 0 66104 800 66224
rect 79200 65832 80000 65952
rect 0 65288 800 65408
rect 79200 65016 80000 65136
rect 0 64472 800 64592
rect 79200 64200 80000 64320
rect 0 63656 800 63776
rect 79200 63384 80000 63504
rect 0 62840 800 62960
rect 79200 62568 80000 62688
rect 0 62024 800 62144
rect 79200 61752 80000 61872
rect 0 61208 800 61328
rect 79200 60936 80000 61056
rect 0 60392 800 60512
rect 79200 60120 80000 60240
rect 0 59576 800 59696
rect 79200 59304 80000 59424
rect 0 58760 800 58880
rect 79200 58488 80000 58608
rect 0 57944 800 58064
rect 79200 57672 80000 57792
rect 0 57128 800 57248
rect 79200 56856 80000 56976
rect 0 56312 800 56432
rect 79200 56040 80000 56160
rect 0 55496 800 55616
rect 79200 55224 80000 55344
rect 0 54680 800 54800
rect 79200 54408 80000 54528
rect 0 53864 800 53984
rect 79200 53592 80000 53712
rect 0 53048 800 53168
rect 79200 52776 80000 52896
rect 0 52232 800 52352
rect 79200 51960 80000 52080
rect 0 51416 800 51536
rect 79200 51144 80000 51264
rect 0 50600 800 50720
rect 79200 50328 80000 50448
rect 0 49784 800 49904
rect 79200 49512 80000 49632
rect 0 48968 800 49088
rect 79200 48696 80000 48816
rect 0 48152 800 48272
rect 79200 47880 80000 48000
rect 0 47336 800 47456
rect 79200 47064 80000 47184
rect 0 46520 800 46640
rect 79200 46248 80000 46368
rect 0 45704 800 45824
rect 79200 45432 80000 45552
rect 0 44888 800 45008
rect 79200 44616 80000 44736
rect 0 44072 800 44192
rect 79200 43800 80000 43920
rect 0 43256 800 43376
rect 79200 42984 80000 43104
rect 0 42440 800 42560
rect 79200 42168 80000 42288
rect 0 41624 800 41744
rect 79200 41352 80000 41472
rect 0 40808 800 40928
rect 79200 40536 80000 40656
rect 0 39992 800 40112
rect 79200 39720 80000 39840
rect 0 39176 800 39296
rect 79200 38904 80000 39024
rect 0 38360 800 38480
rect 79200 38088 80000 38208
rect 0 37544 800 37664
rect 79200 37272 80000 37392
rect 0 36728 800 36848
rect 79200 36456 80000 36576
rect 0 35912 800 36032
rect 79200 35640 80000 35760
rect 0 35096 800 35216
rect 79200 34824 80000 34944
rect 0 34280 800 34400
rect 79200 34008 80000 34128
rect 0 33464 800 33584
rect 79200 33192 80000 33312
rect 0 32648 800 32768
rect 79200 32376 80000 32496
rect 0 31832 800 31952
rect 79200 31560 80000 31680
rect 0 31016 800 31136
rect 79200 30744 80000 30864
rect 0 30200 800 30320
rect 79200 29928 80000 30048
rect 0 29384 800 29504
rect 79200 29112 80000 29232
rect 0 28568 800 28688
rect 79200 28296 80000 28416
rect 0 27752 800 27872
rect 79200 27480 80000 27600
rect 0 26936 800 27056
rect 79200 26664 80000 26784
rect 0 26120 800 26240
rect 79200 25848 80000 25968
rect 0 25304 800 25424
rect 79200 25032 80000 25152
rect 0 24488 800 24608
rect 79200 24216 80000 24336
rect 0 23672 800 23792
rect 79200 23400 80000 23520
rect 0 22856 800 22976
rect 79200 22584 80000 22704
rect 0 22040 800 22160
rect 79200 21768 80000 21888
rect 0 21224 800 21344
rect 79200 20952 80000 21072
rect 0 20408 800 20528
rect 79200 20136 80000 20256
rect 0 19592 800 19712
rect 79200 19320 80000 19440
rect 0 18776 800 18896
rect 79200 18504 80000 18624
rect 0 17960 800 18080
rect 79200 17688 80000 17808
rect 0 17144 800 17264
rect 79200 16872 80000 16992
rect 0 16328 800 16448
rect 79200 16056 80000 16176
rect 0 15512 800 15632
rect 79200 15240 80000 15360
rect 0 14696 800 14816
rect 79200 14424 80000 14544
rect 0 13880 800 14000
rect 79200 13608 80000 13728
rect 0 13064 800 13184
rect 79200 12792 80000 12912
rect 0 12248 800 12368
rect 79200 11976 80000 12096
rect 0 11432 800 11552
rect 79200 11160 80000 11280
rect 0 10616 800 10736
rect 79200 10344 80000 10464
rect 0 9800 800 9920
rect 79200 9528 80000 9648
rect 0 8984 800 9104
rect 79200 8712 80000 8832
rect 0 8168 800 8288
rect 79200 7896 80000 8016
rect 0 7352 800 7472
rect 79200 7080 80000 7200
rect 0 6536 800 6656
rect 79200 6264 80000 6384
rect 0 5720 800 5840
rect 0 4904 800 5024
<< obsm3 >>
rect 798 94864 79200 97409
rect 880 94584 79200 94864
rect 798 94048 79200 94584
rect 880 93776 79200 94048
rect 880 93768 79120 93776
rect 798 93496 79120 93768
rect 798 93232 79200 93496
rect 880 92960 79200 93232
rect 880 92952 79120 92960
rect 798 92680 79120 92952
rect 798 92416 79200 92680
rect 880 92144 79200 92416
rect 880 92136 79120 92144
rect 798 91864 79120 92136
rect 798 91600 79200 91864
rect 880 91328 79200 91600
rect 880 91320 79120 91328
rect 798 91048 79120 91320
rect 798 90784 79200 91048
rect 880 90512 79200 90784
rect 880 90504 79120 90512
rect 798 90232 79120 90504
rect 798 89968 79200 90232
rect 880 89696 79200 89968
rect 880 89688 79120 89696
rect 798 89416 79120 89688
rect 798 89152 79200 89416
rect 880 88880 79200 89152
rect 880 88872 79120 88880
rect 798 88600 79120 88872
rect 798 88336 79200 88600
rect 880 88064 79200 88336
rect 880 88056 79120 88064
rect 798 87784 79120 88056
rect 798 87520 79200 87784
rect 880 87248 79200 87520
rect 880 87240 79120 87248
rect 798 86968 79120 87240
rect 798 86704 79200 86968
rect 880 86432 79200 86704
rect 880 86424 79120 86432
rect 798 86152 79120 86424
rect 798 85888 79200 86152
rect 880 85616 79200 85888
rect 880 85608 79120 85616
rect 798 85336 79120 85608
rect 798 85072 79200 85336
rect 880 84800 79200 85072
rect 880 84792 79120 84800
rect 798 84520 79120 84792
rect 798 84256 79200 84520
rect 880 83984 79200 84256
rect 880 83976 79120 83984
rect 798 83704 79120 83976
rect 798 83440 79200 83704
rect 880 83168 79200 83440
rect 880 83160 79120 83168
rect 798 82888 79120 83160
rect 798 82624 79200 82888
rect 880 82352 79200 82624
rect 880 82344 79120 82352
rect 798 82072 79120 82344
rect 798 81808 79200 82072
rect 880 81536 79200 81808
rect 880 81528 79120 81536
rect 798 81256 79120 81528
rect 798 80992 79200 81256
rect 880 80720 79200 80992
rect 880 80712 79120 80720
rect 798 80440 79120 80712
rect 798 80176 79200 80440
rect 880 79904 79200 80176
rect 880 79896 79120 79904
rect 798 79624 79120 79896
rect 798 79360 79200 79624
rect 880 79088 79200 79360
rect 880 79080 79120 79088
rect 798 78808 79120 79080
rect 798 78544 79200 78808
rect 880 78272 79200 78544
rect 880 78264 79120 78272
rect 798 77992 79120 78264
rect 798 77728 79200 77992
rect 880 77456 79200 77728
rect 880 77448 79120 77456
rect 798 77176 79120 77448
rect 798 76912 79200 77176
rect 880 76640 79200 76912
rect 880 76632 79120 76640
rect 798 76360 79120 76632
rect 798 76096 79200 76360
rect 880 75824 79200 76096
rect 880 75816 79120 75824
rect 798 75544 79120 75816
rect 798 75280 79200 75544
rect 880 75008 79200 75280
rect 880 75000 79120 75008
rect 798 74728 79120 75000
rect 798 74464 79200 74728
rect 880 74192 79200 74464
rect 880 74184 79120 74192
rect 798 73912 79120 74184
rect 798 73648 79200 73912
rect 880 73376 79200 73648
rect 880 73368 79120 73376
rect 798 73096 79120 73368
rect 798 72832 79200 73096
rect 880 72560 79200 72832
rect 880 72552 79120 72560
rect 798 72280 79120 72552
rect 798 72016 79200 72280
rect 880 71744 79200 72016
rect 880 71736 79120 71744
rect 798 71464 79120 71736
rect 798 71200 79200 71464
rect 880 70928 79200 71200
rect 880 70920 79120 70928
rect 798 70648 79120 70920
rect 798 70384 79200 70648
rect 880 70112 79200 70384
rect 880 70104 79120 70112
rect 798 69832 79120 70104
rect 798 69568 79200 69832
rect 880 69296 79200 69568
rect 880 69288 79120 69296
rect 798 69016 79120 69288
rect 798 68752 79200 69016
rect 880 68480 79200 68752
rect 880 68472 79120 68480
rect 798 68200 79120 68472
rect 798 67936 79200 68200
rect 880 67664 79200 67936
rect 880 67656 79120 67664
rect 798 67384 79120 67656
rect 798 67120 79200 67384
rect 880 66848 79200 67120
rect 880 66840 79120 66848
rect 798 66568 79120 66840
rect 798 66304 79200 66568
rect 880 66032 79200 66304
rect 880 66024 79120 66032
rect 798 65752 79120 66024
rect 798 65488 79200 65752
rect 880 65216 79200 65488
rect 880 65208 79120 65216
rect 798 64936 79120 65208
rect 798 64672 79200 64936
rect 880 64400 79200 64672
rect 880 64392 79120 64400
rect 798 64120 79120 64392
rect 798 63856 79200 64120
rect 880 63584 79200 63856
rect 880 63576 79120 63584
rect 798 63304 79120 63576
rect 798 63040 79200 63304
rect 880 62768 79200 63040
rect 880 62760 79120 62768
rect 798 62488 79120 62760
rect 798 62224 79200 62488
rect 880 61952 79200 62224
rect 880 61944 79120 61952
rect 798 61672 79120 61944
rect 798 61408 79200 61672
rect 880 61136 79200 61408
rect 880 61128 79120 61136
rect 798 60856 79120 61128
rect 798 60592 79200 60856
rect 880 60320 79200 60592
rect 880 60312 79120 60320
rect 798 60040 79120 60312
rect 798 59776 79200 60040
rect 880 59504 79200 59776
rect 880 59496 79120 59504
rect 798 59224 79120 59496
rect 798 58960 79200 59224
rect 880 58688 79200 58960
rect 880 58680 79120 58688
rect 798 58408 79120 58680
rect 798 58144 79200 58408
rect 880 57872 79200 58144
rect 880 57864 79120 57872
rect 798 57592 79120 57864
rect 798 57328 79200 57592
rect 880 57056 79200 57328
rect 880 57048 79120 57056
rect 798 56776 79120 57048
rect 798 56512 79200 56776
rect 880 56240 79200 56512
rect 880 56232 79120 56240
rect 798 55960 79120 56232
rect 798 55696 79200 55960
rect 880 55424 79200 55696
rect 880 55416 79120 55424
rect 798 55144 79120 55416
rect 798 54880 79200 55144
rect 880 54608 79200 54880
rect 880 54600 79120 54608
rect 798 54328 79120 54600
rect 798 54064 79200 54328
rect 880 53792 79200 54064
rect 880 53784 79120 53792
rect 798 53512 79120 53784
rect 798 53248 79200 53512
rect 880 52976 79200 53248
rect 880 52968 79120 52976
rect 798 52696 79120 52968
rect 798 52432 79200 52696
rect 880 52160 79200 52432
rect 880 52152 79120 52160
rect 798 51880 79120 52152
rect 798 51616 79200 51880
rect 880 51344 79200 51616
rect 880 51336 79120 51344
rect 798 51064 79120 51336
rect 798 50800 79200 51064
rect 880 50528 79200 50800
rect 880 50520 79120 50528
rect 798 50248 79120 50520
rect 798 49984 79200 50248
rect 880 49712 79200 49984
rect 880 49704 79120 49712
rect 798 49432 79120 49704
rect 798 49168 79200 49432
rect 880 48896 79200 49168
rect 880 48888 79120 48896
rect 798 48616 79120 48888
rect 798 48352 79200 48616
rect 880 48080 79200 48352
rect 880 48072 79120 48080
rect 798 47800 79120 48072
rect 798 47536 79200 47800
rect 880 47264 79200 47536
rect 880 47256 79120 47264
rect 798 46984 79120 47256
rect 798 46720 79200 46984
rect 880 46448 79200 46720
rect 880 46440 79120 46448
rect 798 46168 79120 46440
rect 798 45904 79200 46168
rect 880 45632 79200 45904
rect 880 45624 79120 45632
rect 798 45352 79120 45624
rect 798 45088 79200 45352
rect 880 44816 79200 45088
rect 880 44808 79120 44816
rect 798 44536 79120 44808
rect 798 44272 79200 44536
rect 880 44000 79200 44272
rect 880 43992 79120 44000
rect 798 43720 79120 43992
rect 798 43456 79200 43720
rect 880 43184 79200 43456
rect 880 43176 79120 43184
rect 798 42904 79120 43176
rect 798 42640 79200 42904
rect 880 42368 79200 42640
rect 880 42360 79120 42368
rect 798 42088 79120 42360
rect 798 41824 79200 42088
rect 880 41552 79200 41824
rect 880 41544 79120 41552
rect 798 41272 79120 41544
rect 798 41008 79200 41272
rect 880 40736 79200 41008
rect 880 40728 79120 40736
rect 798 40456 79120 40728
rect 798 40192 79200 40456
rect 880 39920 79200 40192
rect 880 39912 79120 39920
rect 798 39640 79120 39912
rect 798 39376 79200 39640
rect 880 39104 79200 39376
rect 880 39096 79120 39104
rect 798 38824 79120 39096
rect 798 38560 79200 38824
rect 880 38288 79200 38560
rect 880 38280 79120 38288
rect 798 38008 79120 38280
rect 798 37744 79200 38008
rect 880 37472 79200 37744
rect 880 37464 79120 37472
rect 798 37192 79120 37464
rect 798 36928 79200 37192
rect 880 36656 79200 36928
rect 880 36648 79120 36656
rect 798 36376 79120 36648
rect 798 36112 79200 36376
rect 880 35840 79200 36112
rect 880 35832 79120 35840
rect 798 35560 79120 35832
rect 798 35296 79200 35560
rect 880 35024 79200 35296
rect 880 35016 79120 35024
rect 798 34744 79120 35016
rect 798 34480 79200 34744
rect 880 34208 79200 34480
rect 880 34200 79120 34208
rect 798 33928 79120 34200
rect 798 33664 79200 33928
rect 880 33392 79200 33664
rect 880 33384 79120 33392
rect 798 33112 79120 33384
rect 798 32848 79200 33112
rect 880 32576 79200 32848
rect 880 32568 79120 32576
rect 798 32296 79120 32568
rect 798 32032 79200 32296
rect 880 31760 79200 32032
rect 880 31752 79120 31760
rect 798 31480 79120 31752
rect 798 31216 79200 31480
rect 880 30944 79200 31216
rect 880 30936 79120 30944
rect 798 30664 79120 30936
rect 798 30400 79200 30664
rect 880 30128 79200 30400
rect 880 30120 79120 30128
rect 798 29848 79120 30120
rect 798 29584 79200 29848
rect 880 29312 79200 29584
rect 880 29304 79120 29312
rect 798 29032 79120 29304
rect 798 28768 79200 29032
rect 880 28496 79200 28768
rect 880 28488 79120 28496
rect 798 28216 79120 28488
rect 798 27952 79200 28216
rect 880 27680 79200 27952
rect 880 27672 79120 27680
rect 798 27400 79120 27672
rect 798 27136 79200 27400
rect 880 26864 79200 27136
rect 880 26856 79120 26864
rect 798 26584 79120 26856
rect 798 26320 79200 26584
rect 880 26048 79200 26320
rect 880 26040 79120 26048
rect 798 25768 79120 26040
rect 798 25504 79200 25768
rect 880 25232 79200 25504
rect 880 25224 79120 25232
rect 798 24952 79120 25224
rect 798 24688 79200 24952
rect 880 24416 79200 24688
rect 880 24408 79120 24416
rect 798 24136 79120 24408
rect 798 23872 79200 24136
rect 880 23600 79200 23872
rect 880 23592 79120 23600
rect 798 23320 79120 23592
rect 798 23056 79200 23320
rect 880 22784 79200 23056
rect 880 22776 79120 22784
rect 798 22504 79120 22776
rect 798 22240 79200 22504
rect 880 21968 79200 22240
rect 880 21960 79120 21968
rect 798 21688 79120 21960
rect 798 21424 79200 21688
rect 880 21152 79200 21424
rect 880 21144 79120 21152
rect 798 20872 79120 21144
rect 798 20608 79200 20872
rect 880 20336 79200 20608
rect 880 20328 79120 20336
rect 798 20056 79120 20328
rect 798 19792 79200 20056
rect 880 19520 79200 19792
rect 880 19512 79120 19520
rect 798 19240 79120 19512
rect 798 18976 79200 19240
rect 880 18704 79200 18976
rect 880 18696 79120 18704
rect 798 18424 79120 18696
rect 798 18160 79200 18424
rect 880 17888 79200 18160
rect 880 17880 79120 17888
rect 798 17608 79120 17880
rect 798 17344 79200 17608
rect 880 17072 79200 17344
rect 880 17064 79120 17072
rect 798 16792 79120 17064
rect 798 16528 79200 16792
rect 880 16256 79200 16528
rect 880 16248 79120 16256
rect 798 15976 79120 16248
rect 798 15712 79200 15976
rect 880 15440 79200 15712
rect 880 15432 79120 15440
rect 798 15160 79120 15432
rect 798 14896 79200 15160
rect 880 14624 79200 14896
rect 880 14616 79120 14624
rect 798 14344 79120 14616
rect 798 14080 79200 14344
rect 880 13808 79200 14080
rect 880 13800 79120 13808
rect 798 13528 79120 13800
rect 798 13264 79200 13528
rect 880 12992 79200 13264
rect 880 12984 79120 12992
rect 798 12712 79120 12984
rect 798 12448 79200 12712
rect 880 12176 79200 12448
rect 880 12168 79120 12176
rect 798 11896 79120 12168
rect 798 11632 79200 11896
rect 880 11360 79200 11632
rect 880 11352 79120 11360
rect 798 11080 79120 11352
rect 798 10816 79200 11080
rect 880 10544 79200 10816
rect 880 10536 79120 10544
rect 798 10264 79120 10536
rect 798 10000 79200 10264
rect 880 9728 79200 10000
rect 880 9720 79120 9728
rect 798 9448 79120 9720
rect 798 9184 79200 9448
rect 880 8912 79200 9184
rect 880 8904 79120 8912
rect 798 8632 79120 8904
rect 798 8368 79200 8632
rect 880 8096 79200 8368
rect 880 8088 79120 8096
rect 798 7816 79120 8088
rect 798 7552 79200 7816
rect 880 7280 79200 7552
rect 880 7272 79120 7280
rect 798 7000 79120 7272
rect 798 6736 79200 7000
rect 880 6464 79200 6736
rect 880 6456 79120 6464
rect 798 6184 79120 6456
rect 798 5920 79200 6184
rect 880 5640 79200 5920
rect 798 5104 79200 5640
rect 880 4824 79200 5104
rect 798 2143 79200 4824
<< metal4 >>
rect 4208 2128 4528 97424
rect 19568 2128 19888 97424
rect 34928 2128 35248 97424
rect 50288 2128 50608 97424
rect 65648 2128 65968 97424
<< obsm4 >>
rect 1163 5203 4128 80205
rect 4608 5203 19488 80205
rect 19968 5203 34848 80205
rect 35328 5203 50208 80205
rect 50688 5203 65568 80205
rect 66048 5203 76669 80205
<< labels >>
rlabel metal2 s 3422 0 3478 800 6 custom_settings[0]
port 1 nsew signal output
rlabel metal2 s 15382 0 15438 800 6 custom_settings[10]
port 2 nsew signal output
rlabel metal2 s 16578 0 16634 800 6 custom_settings[11]
port 3 nsew signal output
rlabel metal2 s 17774 0 17830 800 6 custom_settings[12]
port 4 nsew signal output
rlabel metal2 s 18970 0 19026 800 6 custom_settings[13]
port 5 nsew signal output
rlabel metal2 s 20166 0 20222 800 6 custom_settings[14]
port 6 nsew signal output
rlabel metal2 s 21362 0 21418 800 6 custom_settings[15]
port 7 nsew signal output
rlabel metal2 s 22558 0 22614 800 6 custom_settings[16]
port 8 nsew signal output
rlabel metal2 s 23754 0 23810 800 6 custom_settings[17]
port 9 nsew signal output
rlabel metal2 s 24950 0 25006 800 6 custom_settings[18]
port 10 nsew signal output
rlabel metal2 s 26146 0 26202 800 6 custom_settings[19]
port 11 nsew signal output
rlabel metal2 s 4618 0 4674 800 6 custom_settings[1]
port 12 nsew signal output
rlabel metal2 s 27342 0 27398 800 6 custom_settings[20]
port 13 nsew signal output
rlabel metal2 s 28538 0 28594 800 6 custom_settings[21]
port 14 nsew signal output
rlabel metal2 s 29734 0 29790 800 6 custom_settings[22]
port 15 nsew signal output
rlabel metal2 s 30930 0 30986 800 6 custom_settings[23]
port 16 nsew signal output
rlabel metal2 s 32126 0 32182 800 6 custom_settings[24]
port 17 nsew signal output
rlabel metal2 s 33322 0 33378 800 6 custom_settings[25]
port 18 nsew signal output
rlabel metal2 s 34518 0 34574 800 6 custom_settings[26]
port 19 nsew signal output
rlabel metal2 s 35714 0 35770 800 6 custom_settings[27]
port 20 nsew signal output
rlabel metal2 s 36910 0 36966 800 6 custom_settings[28]
port 21 nsew signal output
rlabel metal2 s 38106 0 38162 800 6 custom_settings[29]
port 22 nsew signal output
rlabel metal2 s 5814 0 5870 800 6 custom_settings[2]
port 23 nsew signal output
rlabel metal2 s 39302 0 39358 800 6 custom_settings[30]
port 24 nsew signal output
rlabel metal2 s 40498 0 40554 800 6 custom_settings[31]
port 25 nsew signal output
rlabel metal2 s 7010 0 7066 800 6 custom_settings[3]
port 26 nsew signal output
rlabel metal2 s 8206 0 8262 800 6 custom_settings[4]
port 27 nsew signal output
rlabel metal2 s 9402 0 9458 800 6 custom_settings[5]
port 28 nsew signal output
rlabel metal2 s 10598 0 10654 800 6 custom_settings[6]
port 29 nsew signal output
rlabel metal2 s 11794 0 11850 800 6 custom_settings[7]
port 30 nsew signal output
rlabel metal2 s 12990 0 13046 800 6 custom_settings[8]
port 31 nsew signal output
rlabel metal2 s 14186 0 14242 800 6 custom_settings[9]
port 32 nsew signal output
rlabel metal2 s 1490 99200 1546 100000 6 io_in_0
port 33 nsew signal input
rlabel metal3 s 0 4904 800 5024 6 io_oeb[0]
port 34 nsew signal output
rlabel metal3 s 0 13064 800 13184 6 io_oeb[10]
port 35 nsew signal output
rlabel metal3 s 0 13880 800 14000 6 io_oeb[11]
port 36 nsew signal output
rlabel metal3 s 0 14696 800 14816 6 io_oeb[12]
port 37 nsew signal output
rlabel metal3 s 0 15512 800 15632 6 io_oeb[13]
port 38 nsew signal output
rlabel metal3 s 0 16328 800 16448 6 io_oeb[14]
port 39 nsew signal output
rlabel metal3 s 0 17144 800 17264 6 io_oeb[15]
port 40 nsew signal output
rlabel metal3 s 0 17960 800 18080 6 io_oeb[16]
port 41 nsew signal output
rlabel metal3 s 0 18776 800 18896 6 io_oeb[17]
port 42 nsew signal output
rlabel metal3 s 0 19592 800 19712 6 io_oeb[18]
port 43 nsew signal output
rlabel metal3 s 0 20408 800 20528 6 io_oeb[19]
port 44 nsew signal output
rlabel metal3 s 0 5720 800 5840 6 io_oeb[1]
port 45 nsew signal output
rlabel metal3 s 0 21224 800 21344 6 io_oeb[20]
port 46 nsew signal output
rlabel metal3 s 0 22040 800 22160 6 io_oeb[21]
port 47 nsew signal output
rlabel metal3 s 0 22856 800 22976 6 io_oeb[22]
port 48 nsew signal output
rlabel metal3 s 0 23672 800 23792 6 io_oeb[23]
port 49 nsew signal output
rlabel metal3 s 0 24488 800 24608 6 io_oeb[24]
port 50 nsew signal output
rlabel metal3 s 0 25304 800 25424 6 io_oeb[25]
port 51 nsew signal output
rlabel metal3 s 0 26120 800 26240 6 io_oeb[26]
port 52 nsew signal output
rlabel metal3 s 0 26936 800 27056 6 io_oeb[27]
port 53 nsew signal output
rlabel metal3 s 0 27752 800 27872 6 io_oeb[28]
port 54 nsew signal output
rlabel metal3 s 0 28568 800 28688 6 io_oeb[29]
port 55 nsew signal output
rlabel metal3 s 0 6536 800 6656 6 io_oeb[2]
port 56 nsew signal output
rlabel metal3 s 0 29384 800 29504 6 io_oeb[30]
port 57 nsew signal output
rlabel metal3 s 0 30200 800 30320 6 io_oeb[31]
port 58 nsew signal output
rlabel metal3 s 0 31016 800 31136 6 io_oeb[32]
port 59 nsew signal output
rlabel metal3 s 0 31832 800 31952 6 io_oeb[33]
port 60 nsew signal output
rlabel metal3 s 0 32648 800 32768 6 io_oeb[34]
port 61 nsew signal output
rlabel metal3 s 0 33464 800 33584 6 io_oeb[35]
port 62 nsew signal output
rlabel metal3 s 0 34280 800 34400 6 io_oeb[36]
port 63 nsew signal output
rlabel metal3 s 0 35096 800 35216 6 io_oeb[37]
port 64 nsew signal output
rlabel metal3 s 0 7352 800 7472 6 io_oeb[3]
port 65 nsew signal output
rlabel metal3 s 0 8168 800 8288 6 io_oeb[4]
port 66 nsew signal output
rlabel metal3 s 0 8984 800 9104 6 io_oeb[5]
port 67 nsew signal output
rlabel metal3 s 0 9800 800 9920 6 io_oeb[6]
port 68 nsew signal output
rlabel metal3 s 0 10616 800 10736 6 io_oeb[7]
port 69 nsew signal output
rlabel metal3 s 0 11432 800 11552 6 io_oeb[8]
port 70 nsew signal output
rlabel metal3 s 0 12248 800 12368 6 io_oeb[9]
port 71 nsew signal output
rlabel metal3 s 0 66104 800 66224 6 io_oeb_scrapcpu[0]
port 72 nsew signal input
rlabel metal3 s 0 74264 800 74384 6 io_oeb_scrapcpu[10]
port 73 nsew signal input
rlabel metal3 s 0 75080 800 75200 6 io_oeb_scrapcpu[11]
port 74 nsew signal input
rlabel metal3 s 0 75896 800 76016 6 io_oeb_scrapcpu[12]
port 75 nsew signal input
rlabel metal3 s 0 76712 800 76832 6 io_oeb_scrapcpu[13]
port 76 nsew signal input
rlabel metal3 s 0 77528 800 77648 6 io_oeb_scrapcpu[14]
port 77 nsew signal input
rlabel metal3 s 0 78344 800 78464 6 io_oeb_scrapcpu[15]
port 78 nsew signal input
rlabel metal3 s 0 79160 800 79280 6 io_oeb_scrapcpu[16]
port 79 nsew signal input
rlabel metal3 s 0 79976 800 80096 6 io_oeb_scrapcpu[17]
port 80 nsew signal input
rlabel metal3 s 0 80792 800 80912 6 io_oeb_scrapcpu[18]
port 81 nsew signal input
rlabel metal3 s 0 81608 800 81728 6 io_oeb_scrapcpu[19]
port 82 nsew signal input
rlabel metal3 s 0 66920 800 67040 6 io_oeb_scrapcpu[1]
port 83 nsew signal input
rlabel metal3 s 0 82424 800 82544 6 io_oeb_scrapcpu[20]
port 84 nsew signal input
rlabel metal3 s 0 83240 800 83360 6 io_oeb_scrapcpu[21]
port 85 nsew signal input
rlabel metal3 s 0 84056 800 84176 6 io_oeb_scrapcpu[22]
port 86 nsew signal input
rlabel metal3 s 0 84872 800 84992 6 io_oeb_scrapcpu[23]
port 87 nsew signal input
rlabel metal3 s 0 85688 800 85808 6 io_oeb_scrapcpu[24]
port 88 nsew signal input
rlabel metal3 s 0 86504 800 86624 6 io_oeb_scrapcpu[25]
port 89 nsew signal input
rlabel metal3 s 0 87320 800 87440 6 io_oeb_scrapcpu[26]
port 90 nsew signal input
rlabel metal3 s 0 88136 800 88256 6 io_oeb_scrapcpu[27]
port 91 nsew signal input
rlabel metal3 s 0 88952 800 89072 6 io_oeb_scrapcpu[28]
port 92 nsew signal input
rlabel metal3 s 0 89768 800 89888 6 io_oeb_scrapcpu[29]
port 93 nsew signal input
rlabel metal3 s 0 67736 800 67856 6 io_oeb_scrapcpu[2]
port 94 nsew signal input
rlabel metal3 s 0 90584 800 90704 6 io_oeb_scrapcpu[30]
port 95 nsew signal input
rlabel metal3 s 0 91400 800 91520 6 io_oeb_scrapcpu[31]
port 96 nsew signal input
rlabel metal3 s 0 92216 800 92336 6 io_oeb_scrapcpu[32]
port 97 nsew signal input
rlabel metal3 s 0 93032 800 93152 6 io_oeb_scrapcpu[33]
port 98 nsew signal input
rlabel metal3 s 0 93848 800 93968 6 io_oeb_scrapcpu[34]
port 99 nsew signal input
rlabel metal3 s 0 94664 800 94784 6 io_oeb_scrapcpu[35]
port 100 nsew signal input
rlabel metal3 s 0 68552 800 68672 6 io_oeb_scrapcpu[3]
port 101 nsew signal input
rlabel metal3 s 0 69368 800 69488 6 io_oeb_scrapcpu[4]
port 102 nsew signal input
rlabel metal3 s 0 70184 800 70304 6 io_oeb_scrapcpu[5]
port 103 nsew signal input
rlabel metal3 s 0 71000 800 71120 6 io_oeb_scrapcpu[6]
port 104 nsew signal input
rlabel metal3 s 0 71816 800 71936 6 io_oeb_scrapcpu[7]
port 105 nsew signal input
rlabel metal3 s 0 72632 800 72752 6 io_oeb_scrapcpu[8]
port 106 nsew signal input
rlabel metal3 s 0 73448 800 73568 6 io_oeb_scrapcpu[9]
port 107 nsew signal input
rlabel metal2 s 3514 99200 3570 100000 6 io_out[0]
port 108 nsew signal output
rlabel metal2 s 23754 99200 23810 100000 6 io_out[10]
port 109 nsew signal output
rlabel metal2 s 25778 99200 25834 100000 6 io_out[11]
port 110 nsew signal output
rlabel metal2 s 27802 99200 27858 100000 6 io_out[12]
port 111 nsew signal output
rlabel metal2 s 29826 99200 29882 100000 6 io_out[13]
port 112 nsew signal output
rlabel metal2 s 31850 99200 31906 100000 6 io_out[14]
port 113 nsew signal output
rlabel metal2 s 33874 99200 33930 100000 6 io_out[15]
port 114 nsew signal output
rlabel metal2 s 35898 99200 35954 100000 6 io_out[16]
port 115 nsew signal output
rlabel metal2 s 37922 99200 37978 100000 6 io_out[17]
port 116 nsew signal output
rlabel metal2 s 39946 99200 40002 100000 6 io_out[18]
port 117 nsew signal output
rlabel metal2 s 41970 99200 42026 100000 6 io_out[19]
port 118 nsew signal output
rlabel metal2 s 5538 99200 5594 100000 6 io_out[1]
port 119 nsew signal output
rlabel metal2 s 43994 99200 44050 100000 6 io_out[20]
port 120 nsew signal output
rlabel metal2 s 46018 99200 46074 100000 6 io_out[21]
port 121 nsew signal output
rlabel metal2 s 48042 99200 48098 100000 6 io_out[22]
port 122 nsew signal output
rlabel metal2 s 50066 99200 50122 100000 6 io_out[23]
port 123 nsew signal output
rlabel metal2 s 52090 99200 52146 100000 6 io_out[24]
port 124 nsew signal output
rlabel metal2 s 54114 99200 54170 100000 6 io_out[25]
port 125 nsew signal output
rlabel metal2 s 56138 99200 56194 100000 6 io_out[26]
port 126 nsew signal output
rlabel metal2 s 58162 99200 58218 100000 6 io_out[27]
port 127 nsew signal output
rlabel metal2 s 60186 99200 60242 100000 6 io_out[28]
port 128 nsew signal output
rlabel metal2 s 62210 99200 62266 100000 6 io_out[29]
port 129 nsew signal output
rlabel metal2 s 7562 99200 7618 100000 6 io_out[2]
port 130 nsew signal output
rlabel metal2 s 64234 99200 64290 100000 6 io_out[30]
port 131 nsew signal output
rlabel metal2 s 66258 99200 66314 100000 6 io_out[31]
port 132 nsew signal output
rlabel metal2 s 68282 99200 68338 100000 6 io_out[32]
port 133 nsew signal output
rlabel metal2 s 70306 99200 70362 100000 6 io_out[33]
port 134 nsew signal output
rlabel metal2 s 72330 99200 72386 100000 6 io_out[34]
port 135 nsew signal output
rlabel metal2 s 74354 99200 74410 100000 6 io_out[35]
port 136 nsew signal output
rlabel metal2 s 76378 99200 76434 100000 6 io_out[36]
port 137 nsew signal output
rlabel metal2 s 78402 99200 78458 100000 6 io_out[37]
port 138 nsew signal output
rlabel metal2 s 9586 99200 9642 100000 6 io_out[3]
port 139 nsew signal output
rlabel metal2 s 11610 99200 11666 100000 6 io_out[4]
port 140 nsew signal output
rlabel metal2 s 13634 99200 13690 100000 6 io_out[5]
port 141 nsew signal output
rlabel metal2 s 15658 99200 15714 100000 6 io_out[6]
port 142 nsew signal output
rlabel metal2 s 17682 99200 17738 100000 6 io_out[7]
port 143 nsew signal output
rlabel metal2 s 19706 99200 19762 100000 6 io_out[8]
port 144 nsew signal output
rlabel metal2 s 21730 99200 21786 100000 6 io_out[9]
port 145 nsew signal output
rlabel metal3 s 0 36728 800 36848 6 io_out_scrapcpu[0]
port 146 nsew signal input
rlabel metal3 s 0 44888 800 45008 6 io_out_scrapcpu[10]
port 147 nsew signal input
rlabel metal3 s 0 45704 800 45824 6 io_out_scrapcpu[11]
port 148 nsew signal input
rlabel metal3 s 0 46520 800 46640 6 io_out_scrapcpu[12]
port 149 nsew signal input
rlabel metal3 s 0 47336 800 47456 6 io_out_scrapcpu[13]
port 150 nsew signal input
rlabel metal3 s 0 48152 800 48272 6 io_out_scrapcpu[14]
port 151 nsew signal input
rlabel metal3 s 0 48968 800 49088 6 io_out_scrapcpu[15]
port 152 nsew signal input
rlabel metal3 s 0 49784 800 49904 6 io_out_scrapcpu[16]
port 153 nsew signal input
rlabel metal3 s 0 50600 800 50720 6 io_out_scrapcpu[17]
port 154 nsew signal input
rlabel metal3 s 0 51416 800 51536 6 io_out_scrapcpu[18]
port 155 nsew signal input
rlabel metal3 s 0 52232 800 52352 6 io_out_scrapcpu[19]
port 156 nsew signal input
rlabel metal3 s 0 37544 800 37664 6 io_out_scrapcpu[1]
port 157 nsew signal input
rlabel metal3 s 0 53048 800 53168 6 io_out_scrapcpu[20]
port 158 nsew signal input
rlabel metal3 s 0 53864 800 53984 6 io_out_scrapcpu[21]
port 159 nsew signal input
rlabel metal3 s 0 54680 800 54800 6 io_out_scrapcpu[22]
port 160 nsew signal input
rlabel metal3 s 0 55496 800 55616 6 io_out_scrapcpu[23]
port 161 nsew signal input
rlabel metal3 s 0 56312 800 56432 6 io_out_scrapcpu[24]
port 162 nsew signal input
rlabel metal3 s 0 57128 800 57248 6 io_out_scrapcpu[25]
port 163 nsew signal input
rlabel metal3 s 0 57944 800 58064 6 io_out_scrapcpu[26]
port 164 nsew signal input
rlabel metal3 s 0 58760 800 58880 6 io_out_scrapcpu[27]
port 165 nsew signal input
rlabel metal3 s 0 59576 800 59696 6 io_out_scrapcpu[28]
port 166 nsew signal input
rlabel metal3 s 0 60392 800 60512 6 io_out_scrapcpu[29]
port 167 nsew signal input
rlabel metal3 s 0 38360 800 38480 6 io_out_scrapcpu[2]
port 168 nsew signal input
rlabel metal3 s 0 61208 800 61328 6 io_out_scrapcpu[30]
port 169 nsew signal input
rlabel metal3 s 0 62024 800 62144 6 io_out_scrapcpu[31]
port 170 nsew signal input
rlabel metal3 s 0 62840 800 62960 6 io_out_scrapcpu[32]
port 171 nsew signal input
rlabel metal3 s 0 63656 800 63776 6 io_out_scrapcpu[33]
port 172 nsew signal input
rlabel metal3 s 0 64472 800 64592 6 io_out_scrapcpu[34]
port 173 nsew signal input
rlabel metal3 s 0 65288 800 65408 6 io_out_scrapcpu[35]
port 174 nsew signal input
rlabel metal3 s 0 39176 800 39296 6 io_out_scrapcpu[3]
port 175 nsew signal input
rlabel metal3 s 0 39992 800 40112 6 io_out_scrapcpu[4]
port 176 nsew signal input
rlabel metal3 s 0 40808 800 40928 6 io_out_scrapcpu[5]
port 177 nsew signal input
rlabel metal3 s 0 41624 800 41744 6 io_out_scrapcpu[6]
port 178 nsew signal input
rlabel metal3 s 0 42440 800 42560 6 io_out_scrapcpu[7]
port 179 nsew signal input
rlabel metal3 s 0 43256 800 43376 6 io_out_scrapcpu[8]
port 180 nsew signal input
rlabel metal3 s 0 44072 800 44192 6 io_out_scrapcpu[9]
port 181 nsew signal input
rlabel metal3 s 79200 35640 80000 35760 6 la_data_out[0]
port 182 nsew signal output
rlabel metal3 s 79200 43800 80000 43920 6 la_data_out[10]
port 183 nsew signal output
rlabel metal3 s 79200 44616 80000 44736 6 la_data_out[11]
port 184 nsew signal output
rlabel metal3 s 79200 45432 80000 45552 6 la_data_out[12]
port 185 nsew signal output
rlabel metal3 s 79200 46248 80000 46368 6 la_data_out[13]
port 186 nsew signal output
rlabel metal3 s 79200 47064 80000 47184 6 la_data_out[14]
port 187 nsew signal output
rlabel metal3 s 79200 47880 80000 48000 6 la_data_out[15]
port 188 nsew signal output
rlabel metal3 s 79200 48696 80000 48816 6 la_data_out[16]
port 189 nsew signal output
rlabel metal3 s 79200 49512 80000 49632 6 la_data_out[17]
port 190 nsew signal output
rlabel metal3 s 79200 50328 80000 50448 6 la_data_out[18]
port 191 nsew signal output
rlabel metal3 s 79200 51144 80000 51264 6 la_data_out[19]
port 192 nsew signal output
rlabel metal3 s 79200 36456 80000 36576 6 la_data_out[1]
port 193 nsew signal output
rlabel metal3 s 79200 51960 80000 52080 6 la_data_out[20]
port 194 nsew signal output
rlabel metal3 s 79200 52776 80000 52896 6 la_data_out[21]
port 195 nsew signal output
rlabel metal3 s 79200 53592 80000 53712 6 la_data_out[22]
port 196 nsew signal output
rlabel metal3 s 79200 54408 80000 54528 6 la_data_out[23]
port 197 nsew signal output
rlabel metal3 s 79200 55224 80000 55344 6 la_data_out[24]
port 198 nsew signal output
rlabel metal3 s 79200 56040 80000 56160 6 la_data_out[25]
port 199 nsew signal output
rlabel metal3 s 79200 56856 80000 56976 6 la_data_out[26]
port 200 nsew signal output
rlabel metal3 s 79200 57672 80000 57792 6 la_data_out[27]
port 201 nsew signal output
rlabel metal3 s 79200 58488 80000 58608 6 la_data_out[28]
port 202 nsew signal output
rlabel metal3 s 79200 59304 80000 59424 6 la_data_out[29]
port 203 nsew signal output
rlabel metal3 s 79200 37272 80000 37392 6 la_data_out[2]
port 204 nsew signal output
rlabel metal3 s 79200 60120 80000 60240 6 la_data_out[30]
port 205 nsew signal output
rlabel metal3 s 79200 60936 80000 61056 6 la_data_out[31]
port 206 nsew signal output
rlabel metal3 s 79200 61752 80000 61872 6 la_data_out[32]
port 207 nsew signal output
rlabel metal3 s 79200 62568 80000 62688 6 la_data_out[33]
port 208 nsew signal output
rlabel metal3 s 79200 63384 80000 63504 6 la_data_out[34]
port 209 nsew signal output
rlabel metal3 s 79200 64200 80000 64320 6 la_data_out[35]
port 210 nsew signal output
rlabel metal3 s 79200 65016 80000 65136 6 la_data_out[36]
port 211 nsew signal output
rlabel metal3 s 79200 65832 80000 65952 6 la_data_out[37]
port 212 nsew signal output
rlabel metal3 s 79200 66648 80000 66768 6 la_data_out[38]
port 213 nsew signal output
rlabel metal3 s 79200 67464 80000 67584 6 la_data_out[39]
port 214 nsew signal output
rlabel metal3 s 79200 38088 80000 38208 6 la_data_out[3]
port 215 nsew signal output
rlabel metal3 s 79200 38904 80000 39024 6 la_data_out[4]
port 216 nsew signal output
rlabel metal3 s 79200 39720 80000 39840 6 la_data_out[5]
port 217 nsew signal output
rlabel metal3 s 79200 40536 80000 40656 6 la_data_out[6]
port 218 nsew signal output
rlabel metal3 s 79200 41352 80000 41472 6 la_data_out[7]
port 219 nsew signal output
rlabel metal3 s 79200 42168 80000 42288 6 la_data_out[8]
port 220 nsew signal output
rlabel metal3 s 79200 42984 80000 43104 6 la_data_out[9]
port 221 nsew signal output
rlabel metal3 s 0 35912 800 36032 6 rst_scrapcpu
port 222 nsew signal output
rlabel metal4 s 4208 2128 4528 97424 6 vccd1
port 223 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 97424 6 vccd1
port 223 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 97424 6 vccd1
port 223 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 97424 6 vssd1
port 224 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 97424 6 vssd1
port 224 nsew ground bidirectional
rlabel metal2 s 1030 0 1086 800 6 wb_clk_i
port 225 nsew signal input
rlabel metal2 s 2226 0 2282 800 6 wb_rst_i
port 226 nsew signal input
rlabel metal3 s 79200 34824 80000 34944 6 wbs_ack_o
port 227 nsew signal output
rlabel metal2 s 41694 0 41750 800 6 wbs_adr_i[0]
port 228 nsew signal input
rlabel metal2 s 53654 0 53710 800 6 wbs_adr_i[10]
port 229 nsew signal input
rlabel metal2 s 54850 0 54906 800 6 wbs_adr_i[11]
port 230 nsew signal input
rlabel metal2 s 56046 0 56102 800 6 wbs_adr_i[12]
port 231 nsew signal input
rlabel metal2 s 57242 0 57298 800 6 wbs_adr_i[13]
port 232 nsew signal input
rlabel metal2 s 58438 0 58494 800 6 wbs_adr_i[14]
port 233 nsew signal input
rlabel metal2 s 59634 0 59690 800 6 wbs_adr_i[15]
port 234 nsew signal input
rlabel metal2 s 60830 0 60886 800 6 wbs_adr_i[16]
port 235 nsew signal input
rlabel metal2 s 62026 0 62082 800 6 wbs_adr_i[17]
port 236 nsew signal input
rlabel metal2 s 63222 0 63278 800 6 wbs_adr_i[18]
port 237 nsew signal input
rlabel metal2 s 64418 0 64474 800 6 wbs_adr_i[19]
port 238 nsew signal input
rlabel metal2 s 42890 0 42946 800 6 wbs_adr_i[1]
port 239 nsew signal input
rlabel metal2 s 65614 0 65670 800 6 wbs_adr_i[20]
port 240 nsew signal input
rlabel metal2 s 66810 0 66866 800 6 wbs_adr_i[21]
port 241 nsew signal input
rlabel metal2 s 68006 0 68062 800 6 wbs_adr_i[22]
port 242 nsew signal input
rlabel metal2 s 69202 0 69258 800 6 wbs_adr_i[23]
port 243 nsew signal input
rlabel metal2 s 70398 0 70454 800 6 wbs_adr_i[24]
port 244 nsew signal input
rlabel metal2 s 71594 0 71650 800 6 wbs_adr_i[25]
port 245 nsew signal input
rlabel metal2 s 72790 0 72846 800 6 wbs_adr_i[26]
port 246 nsew signal input
rlabel metal2 s 73986 0 74042 800 6 wbs_adr_i[27]
port 247 nsew signal input
rlabel metal2 s 75182 0 75238 800 6 wbs_adr_i[28]
port 248 nsew signal input
rlabel metal2 s 76378 0 76434 800 6 wbs_adr_i[29]
port 249 nsew signal input
rlabel metal2 s 44086 0 44142 800 6 wbs_adr_i[2]
port 250 nsew signal input
rlabel metal2 s 77574 0 77630 800 6 wbs_adr_i[30]
port 251 nsew signal input
rlabel metal2 s 78770 0 78826 800 6 wbs_adr_i[31]
port 252 nsew signal input
rlabel metal2 s 45282 0 45338 800 6 wbs_adr_i[3]
port 253 nsew signal input
rlabel metal2 s 46478 0 46534 800 6 wbs_adr_i[4]
port 254 nsew signal input
rlabel metal2 s 47674 0 47730 800 6 wbs_adr_i[5]
port 255 nsew signal input
rlabel metal2 s 48870 0 48926 800 6 wbs_adr_i[6]
port 256 nsew signal input
rlabel metal2 s 50066 0 50122 800 6 wbs_adr_i[7]
port 257 nsew signal input
rlabel metal2 s 51262 0 51318 800 6 wbs_adr_i[8]
port 258 nsew signal input
rlabel metal2 s 52458 0 52514 800 6 wbs_adr_i[9]
port 259 nsew signal input
rlabel metal3 s 79200 33192 80000 33312 6 wbs_cyc_i
port 260 nsew signal input
rlabel metal3 s 79200 68280 80000 68400 6 wbs_dat_i[0]
port 261 nsew signal input
rlabel metal3 s 79200 76440 80000 76560 6 wbs_dat_i[10]
port 262 nsew signal input
rlabel metal3 s 79200 77256 80000 77376 6 wbs_dat_i[11]
port 263 nsew signal input
rlabel metal3 s 79200 78072 80000 78192 6 wbs_dat_i[12]
port 264 nsew signal input
rlabel metal3 s 79200 78888 80000 79008 6 wbs_dat_i[13]
port 265 nsew signal input
rlabel metal3 s 79200 79704 80000 79824 6 wbs_dat_i[14]
port 266 nsew signal input
rlabel metal3 s 79200 80520 80000 80640 6 wbs_dat_i[15]
port 267 nsew signal input
rlabel metal3 s 79200 81336 80000 81456 6 wbs_dat_i[16]
port 268 nsew signal input
rlabel metal3 s 79200 82152 80000 82272 6 wbs_dat_i[17]
port 269 nsew signal input
rlabel metal3 s 79200 82968 80000 83088 6 wbs_dat_i[18]
port 270 nsew signal input
rlabel metal3 s 79200 83784 80000 83904 6 wbs_dat_i[19]
port 271 nsew signal input
rlabel metal3 s 79200 69096 80000 69216 6 wbs_dat_i[1]
port 272 nsew signal input
rlabel metal3 s 79200 84600 80000 84720 6 wbs_dat_i[20]
port 273 nsew signal input
rlabel metal3 s 79200 85416 80000 85536 6 wbs_dat_i[21]
port 274 nsew signal input
rlabel metal3 s 79200 86232 80000 86352 6 wbs_dat_i[22]
port 275 nsew signal input
rlabel metal3 s 79200 87048 80000 87168 6 wbs_dat_i[23]
port 276 nsew signal input
rlabel metal3 s 79200 87864 80000 87984 6 wbs_dat_i[24]
port 277 nsew signal input
rlabel metal3 s 79200 88680 80000 88800 6 wbs_dat_i[25]
port 278 nsew signal input
rlabel metal3 s 79200 89496 80000 89616 6 wbs_dat_i[26]
port 279 nsew signal input
rlabel metal3 s 79200 90312 80000 90432 6 wbs_dat_i[27]
port 280 nsew signal input
rlabel metal3 s 79200 91128 80000 91248 6 wbs_dat_i[28]
port 281 nsew signal input
rlabel metal3 s 79200 91944 80000 92064 6 wbs_dat_i[29]
port 282 nsew signal input
rlabel metal3 s 79200 69912 80000 70032 6 wbs_dat_i[2]
port 283 nsew signal input
rlabel metal3 s 79200 92760 80000 92880 6 wbs_dat_i[30]
port 284 nsew signal input
rlabel metal3 s 79200 93576 80000 93696 6 wbs_dat_i[31]
port 285 nsew signal input
rlabel metal3 s 79200 70728 80000 70848 6 wbs_dat_i[3]
port 286 nsew signal input
rlabel metal3 s 79200 71544 80000 71664 6 wbs_dat_i[4]
port 287 nsew signal input
rlabel metal3 s 79200 72360 80000 72480 6 wbs_dat_i[5]
port 288 nsew signal input
rlabel metal3 s 79200 73176 80000 73296 6 wbs_dat_i[6]
port 289 nsew signal input
rlabel metal3 s 79200 73992 80000 74112 6 wbs_dat_i[7]
port 290 nsew signal input
rlabel metal3 s 79200 74808 80000 74928 6 wbs_dat_i[8]
port 291 nsew signal input
rlabel metal3 s 79200 75624 80000 75744 6 wbs_dat_i[9]
port 292 nsew signal input
rlabel metal3 s 79200 6264 80000 6384 6 wbs_dat_o[0]
port 293 nsew signal output
rlabel metal3 s 79200 14424 80000 14544 6 wbs_dat_o[10]
port 294 nsew signal output
rlabel metal3 s 79200 15240 80000 15360 6 wbs_dat_o[11]
port 295 nsew signal output
rlabel metal3 s 79200 16056 80000 16176 6 wbs_dat_o[12]
port 296 nsew signal output
rlabel metal3 s 79200 16872 80000 16992 6 wbs_dat_o[13]
port 297 nsew signal output
rlabel metal3 s 79200 17688 80000 17808 6 wbs_dat_o[14]
port 298 nsew signal output
rlabel metal3 s 79200 18504 80000 18624 6 wbs_dat_o[15]
port 299 nsew signal output
rlabel metal3 s 79200 19320 80000 19440 6 wbs_dat_o[16]
port 300 nsew signal output
rlabel metal3 s 79200 20136 80000 20256 6 wbs_dat_o[17]
port 301 nsew signal output
rlabel metal3 s 79200 20952 80000 21072 6 wbs_dat_o[18]
port 302 nsew signal output
rlabel metal3 s 79200 21768 80000 21888 6 wbs_dat_o[19]
port 303 nsew signal output
rlabel metal3 s 79200 7080 80000 7200 6 wbs_dat_o[1]
port 304 nsew signal output
rlabel metal3 s 79200 22584 80000 22704 6 wbs_dat_o[20]
port 305 nsew signal output
rlabel metal3 s 79200 23400 80000 23520 6 wbs_dat_o[21]
port 306 nsew signal output
rlabel metal3 s 79200 24216 80000 24336 6 wbs_dat_o[22]
port 307 nsew signal output
rlabel metal3 s 79200 25032 80000 25152 6 wbs_dat_o[23]
port 308 nsew signal output
rlabel metal3 s 79200 25848 80000 25968 6 wbs_dat_o[24]
port 309 nsew signal output
rlabel metal3 s 79200 26664 80000 26784 6 wbs_dat_o[25]
port 310 nsew signal output
rlabel metal3 s 79200 27480 80000 27600 6 wbs_dat_o[26]
port 311 nsew signal output
rlabel metal3 s 79200 28296 80000 28416 6 wbs_dat_o[27]
port 312 nsew signal output
rlabel metal3 s 79200 29112 80000 29232 6 wbs_dat_o[28]
port 313 nsew signal output
rlabel metal3 s 79200 29928 80000 30048 6 wbs_dat_o[29]
port 314 nsew signal output
rlabel metal3 s 79200 7896 80000 8016 6 wbs_dat_o[2]
port 315 nsew signal output
rlabel metal3 s 79200 30744 80000 30864 6 wbs_dat_o[30]
port 316 nsew signal output
rlabel metal3 s 79200 31560 80000 31680 6 wbs_dat_o[31]
port 317 nsew signal output
rlabel metal3 s 79200 8712 80000 8832 6 wbs_dat_o[3]
port 318 nsew signal output
rlabel metal3 s 79200 9528 80000 9648 6 wbs_dat_o[4]
port 319 nsew signal output
rlabel metal3 s 79200 10344 80000 10464 6 wbs_dat_o[5]
port 320 nsew signal output
rlabel metal3 s 79200 11160 80000 11280 6 wbs_dat_o[6]
port 321 nsew signal output
rlabel metal3 s 79200 11976 80000 12096 6 wbs_dat_o[7]
port 322 nsew signal output
rlabel metal3 s 79200 12792 80000 12912 6 wbs_dat_o[8]
port 323 nsew signal output
rlabel metal3 s 79200 13608 80000 13728 6 wbs_dat_o[9]
port 324 nsew signal output
rlabel metal3 s 79200 34008 80000 34128 6 wbs_stb_i
port 325 nsew signal input
rlabel metal3 s 79200 32376 80000 32496 6 wbs_we_i
port 326 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 80000 100000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 4780526
string GDS_FILE /run/media/tholin/8a6b8802-051e-45a8-8492-771202e4c08a/caravel_user_project/openlane/Multiplexer/runs/24_05_24_23_02/results/signoff/multiplexer.magic.gds
string GDS_START 367830
<< end >>

