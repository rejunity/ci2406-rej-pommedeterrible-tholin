magic
tech sky130B
magscale 1 2
timestamp 1717184365
<< obsli1 >>
rect 1104 2159 38824 197489
<< obsm1 >>
rect 14 2128 39914 197520
<< metal2 >>
rect 754 199200 810 200000
rect 1766 199200 1822 200000
rect 2778 199200 2834 200000
rect 3790 199200 3846 200000
rect 4802 199200 4858 200000
rect 5814 199200 5870 200000
rect 6826 199200 6882 200000
rect 7838 199200 7894 200000
rect 8850 199200 8906 200000
rect 9862 199200 9918 200000
rect 10874 199200 10930 200000
rect 11886 199200 11942 200000
rect 12898 199200 12954 200000
rect 13910 199200 13966 200000
rect 14922 199200 14978 200000
rect 15934 199200 15990 200000
rect 16946 199200 17002 200000
rect 17958 199200 18014 200000
rect 18970 199200 19026 200000
rect 19982 199200 20038 200000
rect 20994 199200 21050 200000
rect 22006 199200 22062 200000
rect 23018 199200 23074 200000
rect 24030 199200 24086 200000
rect 25042 199200 25098 200000
rect 26054 199200 26110 200000
rect 27066 199200 27122 200000
rect 28078 199200 28134 200000
rect 29090 199200 29146 200000
rect 30102 199200 30158 200000
rect 31114 199200 31170 200000
rect 32126 199200 32182 200000
rect 33138 199200 33194 200000
rect 34150 199200 34206 200000
rect 35162 199200 35218 200000
rect 36174 199200 36230 200000
rect 37186 199200 37242 200000
rect 38198 199200 38254 200000
rect 39210 199200 39266 200000
rect 1398 0 1454 800
rect 2594 0 2650 800
rect 3790 0 3846 800
rect 4986 0 5042 800
rect 6182 0 6238 800
rect 7378 0 7434 800
rect 8574 0 8630 800
rect 9770 0 9826 800
rect 10966 0 11022 800
rect 12162 0 12218 800
rect 13358 0 13414 800
rect 14554 0 14610 800
rect 15750 0 15806 800
rect 16946 0 17002 800
rect 18142 0 18198 800
rect 19338 0 19394 800
rect 20534 0 20590 800
rect 21730 0 21786 800
rect 22926 0 22982 800
rect 24122 0 24178 800
rect 25318 0 25374 800
rect 26514 0 26570 800
rect 27710 0 27766 800
rect 28906 0 28962 800
rect 30102 0 30158 800
rect 31298 0 31354 800
rect 32494 0 32550 800
rect 33690 0 33746 800
rect 34886 0 34942 800
rect 36082 0 36138 800
rect 37278 0 37334 800
rect 38474 0 38530 800
<< obsm2 >>
rect 20 199144 698 199322
rect 866 199144 1710 199322
rect 1878 199144 2722 199322
rect 2890 199144 3734 199322
rect 3902 199144 4746 199322
rect 4914 199144 5758 199322
rect 5926 199144 6770 199322
rect 6938 199144 7782 199322
rect 7950 199144 8794 199322
rect 8962 199144 9806 199322
rect 9974 199144 10818 199322
rect 10986 199144 11830 199322
rect 11998 199144 12842 199322
rect 13010 199144 13854 199322
rect 14022 199144 14866 199322
rect 15034 199144 15878 199322
rect 16046 199144 16890 199322
rect 17058 199144 17902 199322
rect 18070 199144 18914 199322
rect 19082 199144 19926 199322
rect 20094 199144 20938 199322
rect 21106 199144 21950 199322
rect 22118 199144 22962 199322
rect 23130 199144 23974 199322
rect 24142 199144 24986 199322
rect 25154 199144 25998 199322
rect 26166 199144 27010 199322
rect 27178 199144 28022 199322
rect 28190 199144 29034 199322
rect 29202 199144 30046 199322
rect 30214 199144 31058 199322
rect 31226 199144 32070 199322
rect 32238 199144 33082 199322
rect 33250 199144 34094 199322
rect 34262 199144 35106 199322
rect 35274 199144 36118 199322
rect 36286 199144 37130 199322
rect 37298 199144 38142 199322
rect 38310 199144 39154 199322
rect 39322 199144 39988 199322
rect 20 856 39988 199144
rect 20 734 1342 856
rect 1510 734 2538 856
rect 2706 734 3734 856
rect 3902 734 4930 856
rect 5098 734 6126 856
rect 6294 734 7322 856
rect 7490 734 8518 856
rect 8686 734 9714 856
rect 9882 734 10910 856
rect 11078 734 12106 856
rect 12274 734 13302 856
rect 13470 734 14498 856
rect 14666 734 15694 856
rect 15862 734 16890 856
rect 17058 734 18086 856
rect 18254 734 19282 856
rect 19450 734 20478 856
rect 20646 734 21674 856
rect 21842 734 22870 856
rect 23038 734 24066 856
rect 24234 734 25262 856
rect 25430 734 26458 856
rect 26626 734 27654 856
rect 27822 734 28850 856
rect 29018 734 30046 856
rect 30214 734 31242 856
rect 31410 734 32438 856
rect 32606 734 33634 856
rect 33802 734 34830 856
rect 34998 734 36026 856
rect 36194 734 37222 856
rect 37390 734 38418 856
rect 38586 734 39988 856
<< metal3 >>
rect 0 197208 800 197328
rect 0 196120 800 196240
rect 0 195032 800 195152
rect 0 193944 800 194064
rect 0 192856 800 192976
rect 0 191768 800 191888
rect 0 190680 800 190800
rect 0 189592 800 189712
rect 39200 188776 40000 188896
rect 0 188504 800 188624
rect 39200 187960 40000 188080
rect 0 187416 800 187536
rect 39200 187144 40000 187264
rect 0 186328 800 186448
rect 39200 186328 40000 186448
rect 39200 185512 40000 185632
rect 0 185240 800 185360
rect 39200 184696 40000 184816
rect 0 184152 800 184272
rect 39200 183880 40000 184000
rect 0 183064 800 183184
rect 39200 183064 40000 183184
rect 39200 182248 40000 182368
rect 0 181976 800 182096
rect 39200 181432 40000 181552
rect 0 180888 800 181008
rect 39200 180616 40000 180736
rect 0 179800 800 179920
rect 39200 179800 40000 179920
rect 39200 178984 40000 179104
rect 0 178712 800 178832
rect 39200 178168 40000 178288
rect 0 177624 800 177744
rect 39200 177352 40000 177472
rect 0 176536 800 176656
rect 39200 176536 40000 176656
rect 39200 175720 40000 175840
rect 0 175448 800 175568
rect 39200 174904 40000 175024
rect 0 174360 800 174480
rect 39200 174088 40000 174208
rect 0 173272 800 173392
rect 39200 173272 40000 173392
rect 39200 172456 40000 172576
rect 0 172184 800 172304
rect 39200 171640 40000 171760
rect 0 171096 800 171216
rect 39200 170824 40000 170944
rect 0 170008 800 170128
rect 39200 170008 40000 170128
rect 39200 169192 40000 169312
rect 0 168920 800 169040
rect 39200 168376 40000 168496
rect 0 167832 800 167952
rect 39200 167560 40000 167680
rect 0 166744 800 166864
rect 39200 166744 40000 166864
rect 39200 165928 40000 166048
rect 0 165656 800 165776
rect 39200 165112 40000 165232
rect 0 164568 800 164688
rect 39200 164296 40000 164416
rect 0 163480 800 163600
rect 39200 163480 40000 163600
rect 39200 162664 40000 162784
rect 0 162392 800 162512
rect 39200 161848 40000 161968
rect 0 161304 800 161424
rect 39200 161032 40000 161152
rect 0 160216 800 160336
rect 39200 160216 40000 160336
rect 39200 159400 40000 159520
rect 0 159128 800 159248
rect 39200 158584 40000 158704
rect 0 158040 800 158160
rect 39200 157768 40000 157888
rect 0 156952 800 157072
rect 39200 156952 40000 157072
rect 39200 156136 40000 156256
rect 0 155864 800 155984
rect 39200 155320 40000 155440
rect 0 154776 800 154896
rect 39200 154504 40000 154624
rect 0 153688 800 153808
rect 39200 153688 40000 153808
rect 39200 152872 40000 152992
rect 0 152600 800 152720
rect 39200 152056 40000 152176
rect 0 151512 800 151632
rect 39200 151240 40000 151360
rect 0 150424 800 150544
rect 39200 150424 40000 150544
rect 39200 149608 40000 149728
rect 0 149336 800 149456
rect 39200 148792 40000 148912
rect 0 148248 800 148368
rect 39200 147976 40000 148096
rect 0 147160 800 147280
rect 39200 147160 40000 147280
rect 39200 146344 40000 146464
rect 0 146072 800 146192
rect 39200 145528 40000 145648
rect 0 144984 800 145104
rect 39200 144712 40000 144832
rect 0 143896 800 144016
rect 39200 143896 40000 144016
rect 39200 143080 40000 143200
rect 0 142808 800 142928
rect 39200 142264 40000 142384
rect 0 141720 800 141840
rect 39200 141448 40000 141568
rect 0 140632 800 140752
rect 39200 140632 40000 140752
rect 39200 139816 40000 139936
rect 0 139544 800 139664
rect 39200 139000 40000 139120
rect 0 138456 800 138576
rect 39200 138184 40000 138304
rect 0 137368 800 137488
rect 39200 137368 40000 137488
rect 39200 136552 40000 136672
rect 0 136280 800 136400
rect 39200 135736 40000 135856
rect 0 135192 800 135312
rect 39200 134920 40000 135040
rect 0 134104 800 134224
rect 39200 134104 40000 134224
rect 39200 133288 40000 133408
rect 0 133016 800 133136
rect 39200 132472 40000 132592
rect 0 131928 800 132048
rect 39200 131656 40000 131776
rect 0 130840 800 130960
rect 39200 130840 40000 130960
rect 39200 130024 40000 130144
rect 0 129752 800 129872
rect 39200 129208 40000 129328
rect 0 128664 800 128784
rect 39200 128392 40000 128512
rect 0 127576 800 127696
rect 39200 127576 40000 127696
rect 39200 126760 40000 126880
rect 0 126488 800 126608
rect 39200 125944 40000 126064
rect 0 125400 800 125520
rect 39200 125128 40000 125248
rect 0 124312 800 124432
rect 39200 124312 40000 124432
rect 39200 123496 40000 123616
rect 0 123224 800 123344
rect 39200 122680 40000 122800
rect 0 122136 800 122256
rect 39200 121864 40000 121984
rect 0 121048 800 121168
rect 39200 121048 40000 121168
rect 39200 120232 40000 120352
rect 0 119960 800 120080
rect 39200 119416 40000 119536
rect 0 118872 800 118992
rect 39200 118600 40000 118720
rect 0 117784 800 117904
rect 39200 117784 40000 117904
rect 39200 116968 40000 117088
rect 0 116696 800 116816
rect 39200 116152 40000 116272
rect 0 115608 800 115728
rect 39200 115336 40000 115456
rect 0 114520 800 114640
rect 39200 114520 40000 114640
rect 39200 113704 40000 113824
rect 0 113432 800 113552
rect 39200 112888 40000 113008
rect 0 112344 800 112464
rect 39200 112072 40000 112192
rect 0 111256 800 111376
rect 39200 111256 40000 111376
rect 39200 110440 40000 110560
rect 0 110168 800 110288
rect 39200 109624 40000 109744
rect 0 109080 800 109200
rect 39200 108808 40000 108928
rect 0 107992 800 108112
rect 39200 107992 40000 108112
rect 39200 107176 40000 107296
rect 0 106904 800 107024
rect 39200 106360 40000 106480
rect 0 105816 800 105936
rect 39200 105544 40000 105664
rect 0 104728 800 104848
rect 39200 104728 40000 104848
rect 39200 103912 40000 104032
rect 0 103640 800 103760
rect 39200 103096 40000 103216
rect 0 102552 800 102672
rect 39200 102280 40000 102400
rect 0 101464 800 101584
rect 39200 101464 40000 101584
rect 39200 100648 40000 100768
rect 0 100376 800 100496
rect 39200 99832 40000 99952
rect 0 99288 800 99408
rect 39200 99016 40000 99136
rect 0 98200 800 98320
rect 39200 98200 40000 98320
rect 39200 97384 40000 97504
rect 0 97112 800 97232
rect 39200 96568 40000 96688
rect 0 96024 800 96144
rect 39200 95752 40000 95872
rect 0 94936 800 95056
rect 39200 94936 40000 95056
rect 39200 94120 40000 94240
rect 0 93848 800 93968
rect 39200 93304 40000 93424
rect 0 92760 800 92880
rect 39200 92488 40000 92608
rect 0 91672 800 91792
rect 39200 91672 40000 91792
rect 39200 90856 40000 90976
rect 0 90584 800 90704
rect 39200 90040 40000 90160
rect 0 89496 800 89616
rect 39200 89224 40000 89344
rect 0 88408 800 88528
rect 39200 88408 40000 88528
rect 39200 87592 40000 87712
rect 0 87320 800 87440
rect 39200 86776 40000 86896
rect 0 86232 800 86352
rect 39200 85960 40000 86080
rect 0 85144 800 85264
rect 39200 85144 40000 85264
rect 39200 84328 40000 84448
rect 0 84056 800 84176
rect 39200 83512 40000 83632
rect 0 82968 800 83088
rect 39200 82696 40000 82816
rect 0 81880 800 82000
rect 39200 81880 40000 82000
rect 39200 81064 40000 81184
rect 0 80792 800 80912
rect 39200 80248 40000 80368
rect 0 79704 800 79824
rect 39200 79432 40000 79552
rect 0 78616 800 78736
rect 39200 78616 40000 78736
rect 39200 77800 40000 77920
rect 0 77528 800 77648
rect 39200 76984 40000 77104
rect 0 76440 800 76560
rect 39200 76168 40000 76288
rect 0 75352 800 75472
rect 39200 75352 40000 75472
rect 39200 74536 40000 74656
rect 0 74264 800 74384
rect 39200 73720 40000 73840
rect 0 73176 800 73296
rect 39200 72904 40000 73024
rect 0 72088 800 72208
rect 39200 72088 40000 72208
rect 39200 71272 40000 71392
rect 0 71000 800 71120
rect 39200 70456 40000 70576
rect 0 69912 800 70032
rect 39200 69640 40000 69760
rect 0 68824 800 68944
rect 39200 68824 40000 68944
rect 39200 68008 40000 68128
rect 0 67736 800 67856
rect 39200 67192 40000 67312
rect 0 66648 800 66768
rect 39200 66376 40000 66496
rect 0 65560 800 65680
rect 39200 65560 40000 65680
rect 39200 64744 40000 64864
rect 0 64472 800 64592
rect 39200 63928 40000 64048
rect 0 63384 800 63504
rect 39200 63112 40000 63232
rect 0 62296 800 62416
rect 39200 62296 40000 62416
rect 39200 61480 40000 61600
rect 0 61208 800 61328
rect 39200 60664 40000 60784
rect 0 60120 800 60240
rect 39200 59848 40000 59968
rect 0 59032 800 59152
rect 39200 59032 40000 59152
rect 39200 58216 40000 58336
rect 0 57944 800 58064
rect 39200 57400 40000 57520
rect 0 56856 800 56976
rect 39200 56584 40000 56704
rect 0 55768 800 55888
rect 39200 55768 40000 55888
rect 39200 54952 40000 55072
rect 0 54680 800 54800
rect 39200 54136 40000 54256
rect 0 53592 800 53712
rect 39200 53320 40000 53440
rect 0 52504 800 52624
rect 39200 52504 40000 52624
rect 39200 51688 40000 51808
rect 0 51416 800 51536
rect 39200 50872 40000 50992
rect 0 50328 800 50448
rect 39200 50056 40000 50176
rect 0 49240 800 49360
rect 39200 49240 40000 49360
rect 39200 48424 40000 48544
rect 0 48152 800 48272
rect 39200 47608 40000 47728
rect 0 47064 800 47184
rect 39200 46792 40000 46912
rect 0 45976 800 46096
rect 39200 45976 40000 46096
rect 39200 45160 40000 45280
rect 0 44888 800 45008
rect 39200 44344 40000 44464
rect 0 43800 800 43920
rect 39200 43528 40000 43648
rect 0 42712 800 42832
rect 39200 42712 40000 42832
rect 39200 41896 40000 42016
rect 0 41624 800 41744
rect 39200 41080 40000 41200
rect 0 40536 800 40656
rect 39200 40264 40000 40384
rect 0 39448 800 39568
rect 39200 39448 40000 39568
rect 39200 38632 40000 38752
rect 0 38360 800 38480
rect 39200 37816 40000 37936
rect 0 37272 800 37392
rect 39200 37000 40000 37120
rect 0 36184 800 36304
rect 39200 36184 40000 36304
rect 39200 35368 40000 35488
rect 0 35096 800 35216
rect 39200 34552 40000 34672
rect 0 34008 800 34128
rect 39200 33736 40000 33856
rect 0 32920 800 33040
rect 39200 32920 40000 33040
rect 39200 32104 40000 32224
rect 0 31832 800 31952
rect 39200 31288 40000 31408
rect 0 30744 800 30864
rect 39200 30472 40000 30592
rect 0 29656 800 29776
rect 39200 29656 40000 29776
rect 39200 28840 40000 28960
rect 0 28568 800 28688
rect 39200 28024 40000 28144
rect 0 27480 800 27600
rect 39200 27208 40000 27328
rect 0 26392 800 26512
rect 39200 26392 40000 26512
rect 39200 25576 40000 25696
rect 0 25304 800 25424
rect 39200 24760 40000 24880
rect 0 24216 800 24336
rect 39200 23944 40000 24064
rect 0 23128 800 23248
rect 39200 23128 40000 23248
rect 39200 22312 40000 22432
rect 0 22040 800 22160
rect 39200 21496 40000 21616
rect 0 20952 800 21072
rect 39200 20680 40000 20800
rect 0 19864 800 19984
rect 39200 19864 40000 19984
rect 39200 19048 40000 19168
rect 0 18776 800 18896
rect 39200 18232 40000 18352
rect 0 17688 800 17808
rect 39200 17416 40000 17536
rect 0 16600 800 16720
rect 39200 16600 40000 16720
rect 39200 15784 40000 15904
rect 0 15512 800 15632
rect 39200 14968 40000 15088
rect 0 14424 800 14544
rect 39200 14152 40000 14272
rect 0 13336 800 13456
rect 39200 13336 40000 13456
rect 39200 12520 40000 12640
rect 0 12248 800 12368
rect 39200 11704 40000 11824
rect 0 11160 800 11280
rect 39200 10888 40000 11008
rect 0 10072 800 10192
rect 0 8984 800 9104
rect 0 7896 800 8016
rect 0 6808 800 6928
rect 0 5720 800 5840
rect 0 4632 800 4752
rect 0 3544 800 3664
rect 0 2456 800 2576
<< obsm3 >>
rect 289 197408 39200 197505
rect 880 197128 39200 197408
rect 289 196320 39200 197128
rect 880 196040 39200 196320
rect 289 195232 39200 196040
rect 880 194952 39200 195232
rect 289 194144 39200 194952
rect 880 193864 39200 194144
rect 289 193056 39200 193864
rect 880 192776 39200 193056
rect 289 191968 39200 192776
rect 880 191688 39200 191968
rect 289 190880 39200 191688
rect 880 190600 39200 190880
rect 289 189792 39200 190600
rect 880 189512 39200 189792
rect 289 188976 39200 189512
rect 289 188704 39120 188976
rect 880 188696 39120 188704
rect 880 188424 39200 188696
rect 289 188160 39200 188424
rect 289 187880 39120 188160
rect 289 187616 39200 187880
rect 880 187344 39200 187616
rect 880 187336 39120 187344
rect 289 187064 39120 187336
rect 289 186528 39200 187064
rect 880 186248 39120 186528
rect 289 185712 39200 186248
rect 289 185440 39120 185712
rect 880 185432 39120 185440
rect 880 185160 39200 185432
rect 289 184896 39200 185160
rect 289 184616 39120 184896
rect 289 184352 39200 184616
rect 880 184080 39200 184352
rect 880 184072 39120 184080
rect 289 183800 39120 184072
rect 289 183264 39200 183800
rect 880 182984 39120 183264
rect 289 182448 39200 182984
rect 289 182176 39120 182448
rect 880 182168 39120 182176
rect 880 181896 39200 182168
rect 289 181632 39200 181896
rect 289 181352 39120 181632
rect 289 181088 39200 181352
rect 880 180816 39200 181088
rect 880 180808 39120 180816
rect 289 180536 39120 180808
rect 289 180000 39200 180536
rect 880 179720 39120 180000
rect 289 179184 39200 179720
rect 289 178912 39120 179184
rect 880 178904 39120 178912
rect 880 178632 39200 178904
rect 289 178368 39200 178632
rect 289 178088 39120 178368
rect 289 177824 39200 178088
rect 880 177552 39200 177824
rect 880 177544 39120 177552
rect 289 177272 39120 177544
rect 289 176736 39200 177272
rect 880 176456 39120 176736
rect 289 175920 39200 176456
rect 289 175648 39120 175920
rect 880 175640 39120 175648
rect 880 175368 39200 175640
rect 289 175104 39200 175368
rect 289 174824 39120 175104
rect 289 174560 39200 174824
rect 880 174288 39200 174560
rect 880 174280 39120 174288
rect 289 174008 39120 174280
rect 289 173472 39200 174008
rect 880 173192 39120 173472
rect 289 172656 39200 173192
rect 289 172384 39120 172656
rect 880 172376 39120 172384
rect 880 172104 39200 172376
rect 289 171840 39200 172104
rect 289 171560 39120 171840
rect 289 171296 39200 171560
rect 880 171024 39200 171296
rect 880 171016 39120 171024
rect 289 170744 39120 171016
rect 289 170208 39200 170744
rect 880 169928 39120 170208
rect 289 169392 39200 169928
rect 289 169120 39120 169392
rect 880 169112 39120 169120
rect 880 168840 39200 169112
rect 289 168576 39200 168840
rect 289 168296 39120 168576
rect 289 168032 39200 168296
rect 880 167760 39200 168032
rect 880 167752 39120 167760
rect 289 167480 39120 167752
rect 289 166944 39200 167480
rect 880 166664 39120 166944
rect 289 166128 39200 166664
rect 289 165856 39120 166128
rect 880 165848 39120 165856
rect 880 165576 39200 165848
rect 289 165312 39200 165576
rect 289 165032 39120 165312
rect 289 164768 39200 165032
rect 880 164496 39200 164768
rect 880 164488 39120 164496
rect 289 164216 39120 164488
rect 289 163680 39200 164216
rect 880 163400 39120 163680
rect 289 162864 39200 163400
rect 289 162592 39120 162864
rect 880 162584 39120 162592
rect 880 162312 39200 162584
rect 289 162048 39200 162312
rect 289 161768 39120 162048
rect 289 161504 39200 161768
rect 880 161232 39200 161504
rect 880 161224 39120 161232
rect 289 160952 39120 161224
rect 289 160416 39200 160952
rect 880 160136 39120 160416
rect 289 159600 39200 160136
rect 289 159328 39120 159600
rect 880 159320 39120 159328
rect 880 159048 39200 159320
rect 289 158784 39200 159048
rect 289 158504 39120 158784
rect 289 158240 39200 158504
rect 880 157968 39200 158240
rect 880 157960 39120 157968
rect 289 157688 39120 157960
rect 289 157152 39200 157688
rect 880 156872 39120 157152
rect 289 156336 39200 156872
rect 289 156064 39120 156336
rect 880 156056 39120 156064
rect 880 155784 39200 156056
rect 289 155520 39200 155784
rect 289 155240 39120 155520
rect 289 154976 39200 155240
rect 880 154704 39200 154976
rect 880 154696 39120 154704
rect 289 154424 39120 154696
rect 289 153888 39200 154424
rect 880 153608 39120 153888
rect 289 153072 39200 153608
rect 289 152800 39120 153072
rect 880 152792 39120 152800
rect 880 152520 39200 152792
rect 289 152256 39200 152520
rect 289 151976 39120 152256
rect 289 151712 39200 151976
rect 880 151440 39200 151712
rect 880 151432 39120 151440
rect 289 151160 39120 151432
rect 289 150624 39200 151160
rect 880 150344 39120 150624
rect 289 149808 39200 150344
rect 289 149536 39120 149808
rect 880 149528 39120 149536
rect 880 149256 39200 149528
rect 289 148992 39200 149256
rect 289 148712 39120 148992
rect 289 148448 39200 148712
rect 880 148176 39200 148448
rect 880 148168 39120 148176
rect 289 147896 39120 148168
rect 289 147360 39200 147896
rect 880 147080 39120 147360
rect 289 146544 39200 147080
rect 289 146272 39120 146544
rect 880 146264 39120 146272
rect 880 145992 39200 146264
rect 289 145728 39200 145992
rect 289 145448 39120 145728
rect 289 145184 39200 145448
rect 880 144912 39200 145184
rect 880 144904 39120 144912
rect 289 144632 39120 144904
rect 289 144096 39200 144632
rect 880 143816 39120 144096
rect 289 143280 39200 143816
rect 289 143008 39120 143280
rect 880 143000 39120 143008
rect 880 142728 39200 143000
rect 289 142464 39200 142728
rect 289 142184 39120 142464
rect 289 141920 39200 142184
rect 880 141648 39200 141920
rect 880 141640 39120 141648
rect 289 141368 39120 141640
rect 289 140832 39200 141368
rect 880 140552 39120 140832
rect 289 140016 39200 140552
rect 289 139744 39120 140016
rect 880 139736 39120 139744
rect 880 139464 39200 139736
rect 289 139200 39200 139464
rect 289 138920 39120 139200
rect 289 138656 39200 138920
rect 880 138384 39200 138656
rect 880 138376 39120 138384
rect 289 138104 39120 138376
rect 289 137568 39200 138104
rect 880 137288 39120 137568
rect 289 136752 39200 137288
rect 289 136480 39120 136752
rect 880 136472 39120 136480
rect 880 136200 39200 136472
rect 289 135936 39200 136200
rect 289 135656 39120 135936
rect 289 135392 39200 135656
rect 880 135120 39200 135392
rect 880 135112 39120 135120
rect 289 134840 39120 135112
rect 289 134304 39200 134840
rect 880 134024 39120 134304
rect 289 133488 39200 134024
rect 289 133216 39120 133488
rect 880 133208 39120 133216
rect 880 132936 39200 133208
rect 289 132672 39200 132936
rect 289 132392 39120 132672
rect 289 132128 39200 132392
rect 880 131856 39200 132128
rect 880 131848 39120 131856
rect 289 131576 39120 131848
rect 289 131040 39200 131576
rect 880 130760 39120 131040
rect 289 130224 39200 130760
rect 289 129952 39120 130224
rect 880 129944 39120 129952
rect 880 129672 39200 129944
rect 289 129408 39200 129672
rect 289 129128 39120 129408
rect 289 128864 39200 129128
rect 880 128592 39200 128864
rect 880 128584 39120 128592
rect 289 128312 39120 128584
rect 289 127776 39200 128312
rect 880 127496 39120 127776
rect 289 126960 39200 127496
rect 289 126688 39120 126960
rect 880 126680 39120 126688
rect 880 126408 39200 126680
rect 289 126144 39200 126408
rect 289 125864 39120 126144
rect 289 125600 39200 125864
rect 880 125328 39200 125600
rect 880 125320 39120 125328
rect 289 125048 39120 125320
rect 289 124512 39200 125048
rect 880 124232 39120 124512
rect 289 123696 39200 124232
rect 289 123424 39120 123696
rect 880 123416 39120 123424
rect 880 123144 39200 123416
rect 289 122880 39200 123144
rect 289 122600 39120 122880
rect 289 122336 39200 122600
rect 880 122064 39200 122336
rect 880 122056 39120 122064
rect 289 121784 39120 122056
rect 289 121248 39200 121784
rect 880 120968 39120 121248
rect 289 120432 39200 120968
rect 289 120160 39120 120432
rect 880 120152 39120 120160
rect 880 119880 39200 120152
rect 289 119616 39200 119880
rect 289 119336 39120 119616
rect 289 119072 39200 119336
rect 880 118800 39200 119072
rect 880 118792 39120 118800
rect 289 118520 39120 118792
rect 289 117984 39200 118520
rect 880 117704 39120 117984
rect 289 117168 39200 117704
rect 289 116896 39120 117168
rect 880 116888 39120 116896
rect 880 116616 39200 116888
rect 289 116352 39200 116616
rect 289 116072 39120 116352
rect 289 115808 39200 116072
rect 880 115536 39200 115808
rect 880 115528 39120 115536
rect 289 115256 39120 115528
rect 289 114720 39200 115256
rect 880 114440 39120 114720
rect 289 113904 39200 114440
rect 289 113632 39120 113904
rect 880 113624 39120 113632
rect 880 113352 39200 113624
rect 289 113088 39200 113352
rect 289 112808 39120 113088
rect 289 112544 39200 112808
rect 880 112272 39200 112544
rect 880 112264 39120 112272
rect 289 111992 39120 112264
rect 289 111456 39200 111992
rect 880 111176 39120 111456
rect 289 110640 39200 111176
rect 289 110368 39120 110640
rect 880 110360 39120 110368
rect 880 110088 39200 110360
rect 289 109824 39200 110088
rect 289 109544 39120 109824
rect 289 109280 39200 109544
rect 880 109008 39200 109280
rect 880 109000 39120 109008
rect 289 108728 39120 109000
rect 289 108192 39200 108728
rect 880 107912 39120 108192
rect 289 107376 39200 107912
rect 289 107104 39120 107376
rect 880 107096 39120 107104
rect 880 106824 39200 107096
rect 289 106560 39200 106824
rect 289 106280 39120 106560
rect 289 106016 39200 106280
rect 880 105744 39200 106016
rect 880 105736 39120 105744
rect 289 105464 39120 105736
rect 289 104928 39200 105464
rect 880 104648 39120 104928
rect 289 104112 39200 104648
rect 289 103840 39120 104112
rect 880 103832 39120 103840
rect 880 103560 39200 103832
rect 289 103296 39200 103560
rect 289 103016 39120 103296
rect 289 102752 39200 103016
rect 880 102480 39200 102752
rect 880 102472 39120 102480
rect 289 102200 39120 102472
rect 289 101664 39200 102200
rect 880 101384 39120 101664
rect 289 100848 39200 101384
rect 289 100576 39120 100848
rect 880 100568 39120 100576
rect 880 100296 39200 100568
rect 289 100032 39200 100296
rect 289 99752 39120 100032
rect 289 99488 39200 99752
rect 880 99216 39200 99488
rect 880 99208 39120 99216
rect 289 98936 39120 99208
rect 289 98400 39200 98936
rect 880 98120 39120 98400
rect 289 97584 39200 98120
rect 289 97312 39120 97584
rect 880 97304 39120 97312
rect 880 97032 39200 97304
rect 289 96768 39200 97032
rect 289 96488 39120 96768
rect 289 96224 39200 96488
rect 880 95952 39200 96224
rect 880 95944 39120 95952
rect 289 95672 39120 95944
rect 289 95136 39200 95672
rect 880 94856 39120 95136
rect 289 94320 39200 94856
rect 289 94048 39120 94320
rect 880 94040 39120 94048
rect 880 93768 39200 94040
rect 289 93504 39200 93768
rect 289 93224 39120 93504
rect 289 92960 39200 93224
rect 880 92688 39200 92960
rect 880 92680 39120 92688
rect 289 92408 39120 92680
rect 289 91872 39200 92408
rect 880 91592 39120 91872
rect 289 91056 39200 91592
rect 289 90784 39120 91056
rect 880 90776 39120 90784
rect 880 90504 39200 90776
rect 289 90240 39200 90504
rect 289 89960 39120 90240
rect 289 89696 39200 89960
rect 880 89424 39200 89696
rect 880 89416 39120 89424
rect 289 89144 39120 89416
rect 289 88608 39200 89144
rect 880 88328 39120 88608
rect 289 87792 39200 88328
rect 289 87520 39120 87792
rect 880 87512 39120 87520
rect 880 87240 39200 87512
rect 289 86976 39200 87240
rect 289 86696 39120 86976
rect 289 86432 39200 86696
rect 880 86160 39200 86432
rect 880 86152 39120 86160
rect 289 85880 39120 86152
rect 289 85344 39200 85880
rect 880 85064 39120 85344
rect 289 84528 39200 85064
rect 289 84256 39120 84528
rect 880 84248 39120 84256
rect 880 83976 39200 84248
rect 289 83712 39200 83976
rect 289 83432 39120 83712
rect 289 83168 39200 83432
rect 880 82896 39200 83168
rect 880 82888 39120 82896
rect 289 82616 39120 82888
rect 289 82080 39200 82616
rect 880 81800 39120 82080
rect 289 81264 39200 81800
rect 289 80992 39120 81264
rect 880 80984 39120 80992
rect 880 80712 39200 80984
rect 289 80448 39200 80712
rect 289 80168 39120 80448
rect 289 79904 39200 80168
rect 880 79632 39200 79904
rect 880 79624 39120 79632
rect 289 79352 39120 79624
rect 289 78816 39200 79352
rect 880 78536 39120 78816
rect 289 78000 39200 78536
rect 289 77728 39120 78000
rect 880 77720 39120 77728
rect 880 77448 39200 77720
rect 289 77184 39200 77448
rect 289 76904 39120 77184
rect 289 76640 39200 76904
rect 880 76368 39200 76640
rect 880 76360 39120 76368
rect 289 76088 39120 76360
rect 289 75552 39200 76088
rect 880 75272 39120 75552
rect 289 74736 39200 75272
rect 289 74464 39120 74736
rect 880 74456 39120 74464
rect 880 74184 39200 74456
rect 289 73920 39200 74184
rect 289 73640 39120 73920
rect 289 73376 39200 73640
rect 880 73104 39200 73376
rect 880 73096 39120 73104
rect 289 72824 39120 73096
rect 289 72288 39200 72824
rect 880 72008 39120 72288
rect 289 71472 39200 72008
rect 289 71200 39120 71472
rect 880 71192 39120 71200
rect 880 70920 39200 71192
rect 289 70656 39200 70920
rect 289 70376 39120 70656
rect 289 70112 39200 70376
rect 880 69840 39200 70112
rect 880 69832 39120 69840
rect 289 69560 39120 69832
rect 289 69024 39200 69560
rect 880 68744 39120 69024
rect 289 68208 39200 68744
rect 289 67936 39120 68208
rect 880 67928 39120 67936
rect 880 67656 39200 67928
rect 289 67392 39200 67656
rect 289 67112 39120 67392
rect 289 66848 39200 67112
rect 880 66576 39200 66848
rect 880 66568 39120 66576
rect 289 66296 39120 66568
rect 289 65760 39200 66296
rect 880 65480 39120 65760
rect 289 64944 39200 65480
rect 289 64672 39120 64944
rect 880 64664 39120 64672
rect 880 64392 39200 64664
rect 289 64128 39200 64392
rect 289 63848 39120 64128
rect 289 63584 39200 63848
rect 880 63312 39200 63584
rect 880 63304 39120 63312
rect 289 63032 39120 63304
rect 289 62496 39200 63032
rect 880 62216 39120 62496
rect 289 61680 39200 62216
rect 289 61408 39120 61680
rect 880 61400 39120 61408
rect 880 61128 39200 61400
rect 289 60864 39200 61128
rect 289 60584 39120 60864
rect 289 60320 39200 60584
rect 880 60048 39200 60320
rect 880 60040 39120 60048
rect 289 59768 39120 60040
rect 289 59232 39200 59768
rect 880 58952 39120 59232
rect 289 58416 39200 58952
rect 289 58144 39120 58416
rect 880 58136 39120 58144
rect 880 57864 39200 58136
rect 289 57600 39200 57864
rect 289 57320 39120 57600
rect 289 57056 39200 57320
rect 880 56784 39200 57056
rect 880 56776 39120 56784
rect 289 56504 39120 56776
rect 289 55968 39200 56504
rect 880 55688 39120 55968
rect 289 55152 39200 55688
rect 289 54880 39120 55152
rect 880 54872 39120 54880
rect 880 54600 39200 54872
rect 289 54336 39200 54600
rect 289 54056 39120 54336
rect 289 53792 39200 54056
rect 880 53520 39200 53792
rect 880 53512 39120 53520
rect 289 53240 39120 53512
rect 289 52704 39200 53240
rect 880 52424 39120 52704
rect 289 51888 39200 52424
rect 289 51616 39120 51888
rect 880 51608 39120 51616
rect 880 51336 39200 51608
rect 289 51072 39200 51336
rect 289 50792 39120 51072
rect 289 50528 39200 50792
rect 880 50256 39200 50528
rect 880 50248 39120 50256
rect 289 49976 39120 50248
rect 289 49440 39200 49976
rect 880 49160 39120 49440
rect 289 48624 39200 49160
rect 289 48352 39120 48624
rect 880 48344 39120 48352
rect 880 48072 39200 48344
rect 289 47808 39200 48072
rect 289 47528 39120 47808
rect 289 47264 39200 47528
rect 880 46992 39200 47264
rect 880 46984 39120 46992
rect 289 46712 39120 46984
rect 289 46176 39200 46712
rect 880 45896 39120 46176
rect 289 45360 39200 45896
rect 289 45088 39120 45360
rect 880 45080 39120 45088
rect 880 44808 39200 45080
rect 289 44544 39200 44808
rect 289 44264 39120 44544
rect 289 44000 39200 44264
rect 880 43728 39200 44000
rect 880 43720 39120 43728
rect 289 43448 39120 43720
rect 289 42912 39200 43448
rect 880 42632 39120 42912
rect 289 42096 39200 42632
rect 289 41824 39120 42096
rect 880 41816 39120 41824
rect 880 41544 39200 41816
rect 289 41280 39200 41544
rect 289 41000 39120 41280
rect 289 40736 39200 41000
rect 880 40464 39200 40736
rect 880 40456 39120 40464
rect 289 40184 39120 40456
rect 289 39648 39200 40184
rect 880 39368 39120 39648
rect 289 38832 39200 39368
rect 289 38560 39120 38832
rect 880 38552 39120 38560
rect 880 38280 39200 38552
rect 289 38016 39200 38280
rect 289 37736 39120 38016
rect 289 37472 39200 37736
rect 880 37200 39200 37472
rect 880 37192 39120 37200
rect 289 36920 39120 37192
rect 289 36384 39200 36920
rect 880 36104 39120 36384
rect 289 35568 39200 36104
rect 289 35296 39120 35568
rect 880 35288 39120 35296
rect 880 35016 39200 35288
rect 289 34752 39200 35016
rect 289 34472 39120 34752
rect 289 34208 39200 34472
rect 880 33936 39200 34208
rect 880 33928 39120 33936
rect 289 33656 39120 33928
rect 289 33120 39200 33656
rect 880 32840 39120 33120
rect 289 32304 39200 32840
rect 289 32032 39120 32304
rect 880 32024 39120 32032
rect 880 31752 39200 32024
rect 289 31488 39200 31752
rect 289 31208 39120 31488
rect 289 30944 39200 31208
rect 880 30672 39200 30944
rect 880 30664 39120 30672
rect 289 30392 39120 30664
rect 289 29856 39200 30392
rect 880 29576 39120 29856
rect 289 29040 39200 29576
rect 289 28768 39120 29040
rect 880 28760 39120 28768
rect 880 28488 39200 28760
rect 289 28224 39200 28488
rect 289 27944 39120 28224
rect 289 27680 39200 27944
rect 880 27408 39200 27680
rect 880 27400 39120 27408
rect 289 27128 39120 27400
rect 289 26592 39200 27128
rect 880 26312 39120 26592
rect 289 25776 39200 26312
rect 289 25504 39120 25776
rect 880 25496 39120 25504
rect 880 25224 39200 25496
rect 289 24960 39200 25224
rect 289 24680 39120 24960
rect 289 24416 39200 24680
rect 880 24144 39200 24416
rect 880 24136 39120 24144
rect 289 23864 39120 24136
rect 289 23328 39200 23864
rect 880 23048 39120 23328
rect 289 22512 39200 23048
rect 289 22240 39120 22512
rect 880 22232 39120 22240
rect 880 21960 39200 22232
rect 289 21696 39200 21960
rect 289 21416 39120 21696
rect 289 21152 39200 21416
rect 880 20880 39200 21152
rect 880 20872 39120 20880
rect 289 20600 39120 20872
rect 289 20064 39200 20600
rect 880 19784 39120 20064
rect 289 19248 39200 19784
rect 289 18976 39120 19248
rect 880 18968 39120 18976
rect 880 18696 39200 18968
rect 289 18432 39200 18696
rect 289 18152 39120 18432
rect 289 17888 39200 18152
rect 880 17616 39200 17888
rect 880 17608 39120 17616
rect 289 17336 39120 17608
rect 289 16800 39200 17336
rect 880 16520 39120 16800
rect 289 15984 39200 16520
rect 289 15712 39120 15984
rect 880 15704 39120 15712
rect 880 15432 39200 15704
rect 289 15168 39200 15432
rect 289 14888 39120 15168
rect 289 14624 39200 14888
rect 880 14352 39200 14624
rect 880 14344 39120 14352
rect 289 14072 39120 14344
rect 289 13536 39200 14072
rect 880 13256 39120 13536
rect 289 12720 39200 13256
rect 289 12448 39120 12720
rect 880 12440 39120 12448
rect 880 12168 39200 12440
rect 289 11904 39200 12168
rect 289 11624 39120 11904
rect 289 11360 39200 11624
rect 880 11088 39200 11360
rect 880 11080 39120 11088
rect 289 10808 39120 11080
rect 289 10272 39200 10808
rect 880 9992 39200 10272
rect 289 9184 39200 9992
rect 880 8904 39200 9184
rect 289 8096 39200 8904
rect 880 7816 39200 8096
rect 289 7008 39200 7816
rect 880 6728 39200 7008
rect 289 5920 39200 6728
rect 880 5640 39200 5920
rect 289 4832 39200 5640
rect 880 4552 39200 4832
rect 289 3744 39200 4552
rect 880 3464 39200 3744
rect 289 2656 39200 3464
rect 880 2376 39200 2656
rect 289 2143 39200 2376
<< metal4 >>
rect 4208 2128 4528 197520
rect 19568 2128 19888 197520
rect 34928 2128 35248 197520
<< obsm4 >>
rect 611 3979 4128 181389
rect 4608 3979 19488 181389
rect 19968 3979 34848 181389
rect 35328 3979 37109 181389
<< labels >>
rlabel metal3 s 0 2456 800 2576 6 custom_settings[0]
port 1 nsew signal output
rlabel metal3 s 0 13336 800 13456 6 custom_settings[10]
port 2 nsew signal output
rlabel metal3 s 0 14424 800 14544 6 custom_settings[11]
port 3 nsew signal output
rlabel metal3 s 0 15512 800 15632 6 custom_settings[12]
port 4 nsew signal output
rlabel metal3 s 0 16600 800 16720 6 custom_settings[13]
port 5 nsew signal output
rlabel metal3 s 0 17688 800 17808 6 custom_settings[14]
port 6 nsew signal output
rlabel metal3 s 0 18776 800 18896 6 custom_settings[15]
port 7 nsew signal output
rlabel metal3 s 0 19864 800 19984 6 custom_settings[16]
port 8 nsew signal output
rlabel metal3 s 0 20952 800 21072 6 custom_settings[17]
port 9 nsew signal output
rlabel metal3 s 0 22040 800 22160 6 custom_settings[18]
port 10 nsew signal output
rlabel metal3 s 0 23128 800 23248 6 custom_settings[19]
port 11 nsew signal output
rlabel metal3 s 0 3544 800 3664 6 custom_settings[1]
port 12 nsew signal output
rlabel metal3 s 0 24216 800 24336 6 custom_settings[20]
port 13 nsew signal output
rlabel metal3 s 0 25304 800 25424 6 custom_settings[21]
port 14 nsew signal output
rlabel metal3 s 0 26392 800 26512 6 custom_settings[22]
port 15 nsew signal output
rlabel metal3 s 0 27480 800 27600 6 custom_settings[23]
port 16 nsew signal output
rlabel metal3 s 0 28568 800 28688 6 custom_settings[24]
port 17 nsew signal output
rlabel metal3 s 0 29656 800 29776 6 custom_settings[25]
port 18 nsew signal output
rlabel metal3 s 0 30744 800 30864 6 custom_settings[26]
port 19 nsew signal output
rlabel metal3 s 0 31832 800 31952 6 custom_settings[27]
port 20 nsew signal output
rlabel metal3 s 0 32920 800 33040 6 custom_settings[28]
port 21 nsew signal output
rlabel metal3 s 0 34008 800 34128 6 custom_settings[29]
port 22 nsew signal output
rlabel metal3 s 0 4632 800 4752 6 custom_settings[2]
port 23 nsew signal output
rlabel metal3 s 0 35096 800 35216 6 custom_settings[30]
port 24 nsew signal output
rlabel metal3 s 0 36184 800 36304 6 custom_settings[31]
port 25 nsew signal output
rlabel metal3 s 0 5720 800 5840 6 custom_settings[3]
port 26 nsew signal output
rlabel metal3 s 0 6808 800 6928 6 custom_settings[4]
port 27 nsew signal output
rlabel metal3 s 0 7896 800 8016 6 custom_settings[5]
port 28 nsew signal output
rlabel metal3 s 0 8984 800 9104 6 custom_settings[6]
port 29 nsew signal output
rlabel metal3 s 0 10072 800 10192 6 custom_settings[7]
port 30 nsew signal output
rlabel metal3 s 0 11160 800 11280 6 custom_settings[8]
port 31 nsew signal output
rlabel metal3 s 0 12248 800 12368 6 custom_settings[9]
port 32 nsew signal output
rlabel metal2 s 754 199200 810 200000 6 io_in_0
port 33 nsew signal input
rlabel metal3 s 0 37272 800 37392 6 io_oeb[0]
port 34 nsew signal output
rlabel metal3 s 0 48152 800 48272 6 io_oeb[10]
port 35 nsew signal output
rlabel metal3 s 0 49240 800 49360 6 io_oeb[11]
port 36 nsew signal output
rlabel metal3 s 0 50328 800 50448 6 io_oeb[12]
port 37 nsew signal output
rlabel metal3 s 0 51416 800 51536 6 io_oeb[13]
port 38 nsew signal output
rlabel metal3 s 0 52504 800 52624 6 io_oeb[14]
port 39 nsew signal output
rlabel metal3 s 0 53592 800 53712 6 io_oeb[15]
port 40 nsew signal output
rlabel metal3 s 0 54680 800 54800 6 io_oeb[16]
port 41 nsew signal output
rlabel metal3 s 0 55768 800 55888 6 io_oeb[17]
port 42 nsew signal output
rlabel metal3 s 0 56856 800 56976 6 io_oeb[18]
port 43 nsew signal output
rlabel metal3 s 0 57944 800 58064 6 io_oeb[19]
port 44 nsew signal output
rlabel metal3 s 0 38360 800 38480 6 io_oeb[1]
port 45 nsew signal output
rlabel metal3 s 0 59032 800 59152 6 io_oeb[20]
port 46 nsew signal output
rlabel metal3 s 0 60120 800 60240 6 io_oeb[21]
port 47 nsew signal output
rlabel metal3 s 0 61208 800 61328 6 io_oeb[22]
port 48 nsew signal output
rlabel metal3 s 0 62296 800 62416 6 io_oeb[23]
port 49 nsew signal output
rlabel metal3 s 0 63384 800 63504 6 io_oeb[24]
port 50 nsew signal output
rlabel metal3 s 0 64472 800 64592 6 io_oeb[25]
port 51 nsew signal output
rlabel metal3 s 0 65560 800 65680 6 io_oeb[26]
port 52 nsew signal output
rlabel metal3 s 0 66648 800 66768 6 io_oeb[27]
port 53 nsew signal output
rlabel metal3 s 0 67736 800 67856 6 io_oeb[28]
port 54 nsew signal output
rlabel metal3 s 0 68824 800 68944 6 io_oeb[29]
port 55 nsew signal output
rlabel metal3 s 0 39448 800 39568 6 io_oeb[2]
port 56 nsew signal output
rlabel metal3 s 0 69912 800 70032 6 io_oeb[30]
port 57 nsew signal output
rlabel metal3 s 0 71000 800 71120 6 io_oeb[31]
port 58 nsew signal output
rlabel metal3 s 0 72088 800 72208 6 io_oeb[32]
port 59 nsew signal output
rlabel metal3 s 0 73176 800 73296 6 io_oeb[33]
port 60 nsew signal output
rlabel metal3 s 0 74264 800 74384 6 io_oeb[34]
port 61 nsew signal output
rlabel metal3 s 0 75352 800 75472 6 io_oeb[35]
port 62 nsew signal output
rlabel metal3 s 0 76440 800 76560 6 io_oeb[36]
port 63 nsew signal output
rlabel metal3 s 0 77528 800 77648 6 io_oeb[37]
port 64 nsew signal output
rlabel metal3 s 0 40536 800 40656 6 io_oeb[3]
port 65 nsew signal output
rlabel metal3 s 0 41624 800 41744 6 io_oeb[4]
port 66 nsew signal output
rlabel metal3 s 0 42712 800 42832 6 io_oeb[5]
port 67 nsew signal output
rlabel metal3 s 0 43800 800 43920 6 io_oeb[6]
port 68 nsew signal output
rlabel metal3 s 0 44888 800 45008 6 io_oeb[7]
port 69 nsew signal output
rlabel metal3 s 0 45976 800 46096 6 io_oeb[8]
port 70 nsew signal output
rlabel metal3 s 0 47064 800 47184 6 io_oeb[9]
port 71 nsew signal output
rlabel metal3 s 0 159128 800 159248 6 io_oeb_scrapcpu[0]
port 72 nsew signal input
rlabel metal3 s 0 170008 800 170128 6 io_oeb_scrapcpu[10]
port 73 nsew signal input
rlabel metal3 s 0 171096 800 171216 6 io_oeb_scrapcpu[11]
port 74 nsew signal input
rlabel metal3 s 0 172184 800 172304 6 io_oeb_scrapcpu[12]
port 75 nsew signal input
rlabel metal3 s 0 173272 800 173392 6 io_oeb_scrapcpu[13]
port 76 nsew signal input
rlabel metal3 s 0 174360 800 174480 6 io_oeb_scrapcpu[14]
port 77 nsew signal input
rlabel metal3 s 0 175448 800 175568 6 io_oeb_scrapcpu[15]
port 78 nsew signal input
rlabel metal3 s 0 176536 800 176656 6 io_oeb_scrapcpu[16]
port 79 nsew signal input
rlabel metal3 s 0 177624 800 177744 6 io_oeb_scrapcpu[17]
port 80 nsew signal input
rlabel metal3 s 0 178712 800 178832 6 io_oeb_scrapcpu[18]
port 81 nsew signal input
rlabel metal3 s 0 179800 800 179920 6 io_oeb_scrapcpu[19]
port 82 nsew signal input
rlabel metal3 s 0 160216 800 160336 6 io_oeb_scrapcpu[1]
port 83 nsew signal input
rlabel metal3 s 0 180888 800 181008 6 io_oeb_scrapcpu[20]
port 84 nsew signal input
rlabel metal3 s 0 181976 800 182096 6 io_oeb_scrapcpu[21]
port 85 nsew signal input
rlabel metal3 s 0 183064 800 183184 6 io_oeb_scrapcpu[22]
port 86 nsew signal input
rlabel metal3 s 0 184152 800 184272 6 io_oeb_scrapcpu[23]
port 87 nsew signal input
rlabel metal3 s 0 185240 800 185360 6 io_oeb_scrapcpu[24]
port 88 nsew signal input
rlabel metal3 s 0 186328 800 186448 6 io_oeb_scrapcpu[25]
port 89 nsew signal input
rlabel metal3 s 0 187416 800 187536 6 io_oeb_scrapcpu[26]
port 90 nsew signal input
rlabel metal3 s 0 188504 800 188624 6 io_oeb_scrapcpu[27]
port 91 nsew signal input
rlabel metal3 s 0 189592 800 189712 6 io_oeb_scrapcpu[28]
port 92 nsew signal input
rlabel metal3 s 0 190680 800 190800 6 io_oeb_scrapcpu[29]
port 93 nsew signal input
rlabel metal3 s 0 161304 800 161424 6 io_oeb_scrapcpu[2]
port 94 nsew signal input
rlabel metal3 s 0 191768 800 191888 6 io_oeb_scrapcpu[30]
port 95 nsew signal input
rlabel metal3 s 0 192856 800 192976 6 io_oeb_scrapcpu[31]
port 96 nsew signal input
rlabel metal3 s 0 193944 800 194064 6 io_oeb_scrapcpu[32]
port 97 nsew signal input
rlabel metal3 s 0 195032 800 195152 6 io_oeb_scrapcpu[33]
port 98 nsew signal input
rlabel metal3 s 0 196120 800 196240 6 io_oeb_scrapcpu[34]
port 99 nsew signal input
rlabel metal3 s 0 197208 800 197328 6 io_oeb_scrapcpu[35]
port 100 nsew signal input
rlabel metal3 s 0 162392 800 162512 6 io_oeb_scrapcpu[3]
port 101 nsew signal input
rlabel metal3 s 0 163480 800 163600 6 io_oeb_scrapcpu[4]
port 102 nsew signal input
rlabel metal3 s 0 164568 800 164688 6 io_oeb_scrapcpu[5]
port 103 nsew signal input
rlabel metal3 s 0 165656 800 165776 6 io_oeb_scrapcpu[6]
port 104 nsew signal input
rlabel metal3 s 0 166744 800 166864 6 io_oeb_scrapcpu[7]
port 105 nsew signal input
rlabel metal3 s 0 167832 800 167952 6 io_oeb_scrapcpu[8]
port 106 nsew signal input
rlabel metal3 s 0 168920 800 169040 6 io_oeb_scrapcpu[9]
port 107 nsew signal input
rlabel metal3 s 0 119960 800 120080 6 io_oeb_vliw[0]
port 108 nsew signal input
rlabel metal3 s 0 130840 800 130960 6 io_oeb_vliw[10]
port 109 nsew signal input
rlabel metal3 s 0 131928 800 132048 6 io_oeb_vliw[11]
port 110 nsew signal input
rlabel metal3 s 0 133016 800 133136 6 io_oeb_vliw[12]
port 111 nsew signal input
rlabel metal3 s 0 134104 800 134224 6 io_oeb_vliw[13]
port 112 nsew signal input
rlabel metal3 s 0 135192 800 135312 6 io_oeb_vliw[14]
port 113 nsew signal input
rlabel metal3 s 0 136280 800 136400 6 io_oeb_vliw[15]
port 114 nsew signal input
rlabel metal3 s 0 137368 800 137488 6 io_oeb_vliw[16]
port 115 nsew signal input
rlabel metal3 s 0 138456 800 138576 6 io_oeb_vliw[17]
port 116 nsew signal input
rlabel metal3 s 0 139544 800 139664 6 io_oeb_vliw[18]
port 117 nsew signal input
rlabel metal3 s 0 140632 800 140752 6 io_oeb_vliw[19]
port 118 nsew signal input
rlabel metal3 s 0 121048 800 121168 6 io_oeb_vliw[1]
port 119 nsew signal input
rlabel metal3 s 0 141720 800 141840 6 io_oeb_vliw[20]
port 120 nsew signal input
rlabel metal3 s 0 142808 800 142928 6 io_oeb_vliw[21]
port 121 nsew signal input
rlabel metal3 s 0 143896 800 144016 6 io_oeb_vliw[22]
port 122 nsew signal input
rlabel metal3 s 0 144984 800 145104 6 io_oeb_vliw[23]
port 123 nsew signal input
rlabel metal3 s 0 146072 800 146192 6 io_oeb_vliw[24]
port 124 nsew signal input
rlabel metal3 s 0 147160 800 147280 6 io_oeb_vliw[25]
port 125 nsew signal input
rlabel metal3 s 0 148248 800 148368 6 io_oeb_vliw[26]
port 126 nsew signal input
rlabel metal3 s 0 149336 800 149456 6 io_oeb_vliw[27]
port 127 nsew signal input
rlabel metal3 s 0 150424 800 150544 6 io_oeb_vliw[28]
port 128 nsew signal input
rlabel metal3 s 0 151512 800 151632 6 io_oeb_vliw[29]
port 129 nsew signal input
rlabel metal3 s 0 122136 800 122256 6 io_oeb_vliw[2]
port 130 nsew signal input
rlabel metal3 s 0 152600 800 152720 6 io_oeb_vliw[30]
port 131 nsew signal input
rlabel metal3 s 0 153688 800 153808 6 io_oeb_vliw[31]
port 132 nsew signal input
rlabel metal3 s 0 154776 800 154896 6 io_oeb_vliw[32]
port 133 nsew signal input
rlabel metal3 s 0 155864 800 155984 6 io_oeb_vliw[33]
port 134 nsew signal input
rlabel metal3 s 0 156952 800 157072 6 io_oeb_vliw[34]
port 135 nsew signal input
rlabel metal3 s 0 158040 800 158160 6 io_oeb_vliw[35]
port 136 nsew signal input
rlabel metal3 s 0 123224 800 123344 6 io_oeb_vliw[3]
port 137 nsew signal input
rlabel metal3 s 0 124312 800 124432 6 io_oeb_vliw[4]
port 138 nsew signal input
rlabel metal3 s 0 125400 800 125520 6 io_oeb_vliw[5]
port 139 nsew signal input
rlabel metal3 s 0 126488 800 126608 6 io_oeb_vliw[6]
port 140 nsew signal input
rlabel metal3 s 0 127576 800 127696 6 io_oeb_vliw[7]
port 141 nsew signal input
rlabel metal3 s 0 128664 800 128784 6 io_oeb_vliw[8]
port 142 nsew signal input
rlabel metal3 s 0 129752 800 129872 6 io_oeb_vliw[9]
port 143 nsew signal input
rlabel metal3 s 39200 130840 40000 130960 6 io_oeb_z80[0]
port 144 nsew signal input
rlabel metal3 s 39200 139000 40000 139120 6 io_oeb_z80[10]
port 145 nsew signal input
rlabel metal3 s 39200 139816 40000 139936 6 io_oeb_z80[11]
port 146 nsew signal input
rlabel metal3 s 39200 140632 40000 140752 6 io_oeb_z80[12]
port 147 nsew signal input
rlabel metal3 s 39200 141448 40000 141568 6 io_oeb_z80[13]
port 148 nsew signal input
rlabel metal3 s 39200 142264 40000 142384 6 io_oeb_z80[14]
port 149 nsew signal input
rlabel metal3 s 39200 143080 40000 143200 6 io_oeb_z80[15]
port 150 nsew signal input
rlabel metal3 s 39200 143896 40000 144016 6 io_oeb_z80[16]
port 151 nsew signal input
rlabel metal3 s 39200 144712 40000 144832 6 io_oeb_z80[17]
port 152 nsew signal input
rlabel metal3 s 39200 145528 40000 145648 6 io_oeb_z80[18]
port 153 nsew signal input
rlabel metal3 s 39200 146344 40000 146464 6 io_oeb_z80[19]
port 154 nsew signal input
rlabel metal3 s 39200 131656 40000 131776 6 io_oeb_z80[1]
port 155 nsew signal input
rlabel metal3 s 39200 147160 40000 147280 6 io_oeb_z80[20]
port 156 nsew signal input
rlabel metal3 s 39200 147976 40000 148096 6 io_oeb_z80[21]
port 157 nsew signal input
rlabel metal3 s 39200 148792 40000 148912 6 io_oeb_z80[22]
port 158 nsew signal input
rlabel metal3 s 39200 149608 40000 149728 6 io_oeb_z80[23]
port 159 nsew signal input
rlabel metal3 s 39200 150424 40000 150544 6 io_oeb_z80[24]
port 160 nsew signal input
rlabel metal3 s 39200 151240 40000 151360 6 io_oeb_z80[25]
port 161 nsew signal input
rlabel metal3 s 39200 152056 40000 152176 6 io_oeb_z80[26]
port 162 nsew signal input
rlabel metal3 s 39200 152872 40000 152992 6 io_oeb_z80[27]
port 163 nsew signal input
rlabel metal3 s 39200 153688 40000 153808 6 io_oeb_z80[28]
port 164 nsew signal input
rlabel metal3 s 39200 154504 40000 154624 6 io_oeb_z80[29]
port 165 nsew signal input
rlabel metal3 s 39200 132472 40000 132592 6 io_oeb_z80[2]
port 166 nsew signal input
rlabel metal3 s 39200 155320 40000 155440 6 io_oeb_z80[30]
port 167 nsew signal input
rlabel metal3 s 39200 156136 40000 156256 6 io_oeb_z80[31]
port 168 nsew signal input
rlabel metal3 s 39200 156952 40000 157072 6 io_oeb_z80[32]
port 169 nsew signal input
rlabel metal3 s 39200 157768 40000 157888 6 io_oeb_z80[33]
port 170 nsew signal input
rlabel metal3 s 39200 158584 40000 158704 6 io_oeb_z80[34]
port 171 nsew signal input
rlabel metal3 s 39200 159400 40000 159520 6 io_oeb_z80[35]
port 172 nsew signal input
rlabel metal3 s 39200 133288 40000 133408 6 io_oeb_z80[3]
port 173 nsew signal input
rlabel metal3 s 39200 134104 40000 134224 6 io_oeb_z80[4]
port 174 nsew signal input
rlabel metal3 s 39200 134920 40000 135040 6 io_oeb_z80[5]
port 175 nsew signal input
rlabel metal3 s 39200 135736 40000 135856 6 io_oeb_z80[6]
port 176 nsew signal input
rlabel metal3 s 39200 136552 40000 136672 6 io_oeb_z80[7]
port 177 nsew signal input
rlabel metal3 s 39200 137368 40000 137488 6 io_oeb_z80[8]
port 178 nsew signal input
rlabel metal3 s 39200 138184 40000 138304 6 io_oeb_z80[9]
port 179 nsew signal input
rlabel metal3 s 39200 10888 40000 11008 6 io_out[0]
port 180 nsew signal output
rlabel metal3 s 39200 19048 40000 19168 6 io_out[10]
port 181 nsew signal output
rlabel metal3 s 39200 19864 40000 19984 6 io_out[11]
port 182 nsew signal output
rlabel metal3 s 39200 20680 40000 20800 6 io_out[12]
port 183 nsew signal output
rlabel metal3 s 39200 21496 40000 21616 6 io_out[13]
port 184 nsew signal output
rlabel metal3 s 39200 22312 40000 22432 6 io_out[14]
port 185 nsew signal output
rlabel metal3 s 39200 23128 40000 23248 6 io_out[15]
port 186 nsew signal output
rlabel metal3 s 39200 23944 40000 24064 6 io_out[16]
port 187 nsew signal output
rlabel metal3 s 39200 24760 40000 24880 6 io_out[17]
port 188 nsew signal output
rlabel metal3 s 39200 25576 40000 25696 6 io_out[18]
port 189 nsew signal output
rlabel metal3 s 39200 26392 40000 26512 6 io_out[19]
port 190 nsew signal output
rlabel metal3 s 39200 11704 40000 11824 6 io_out[1]
port 191 nsew signal output
rlabel metal3 s 39200 27208 40000 27328 6 io_out[20]
port 192 nsew signal output
rlabel metal3 s 39200 28024 40000 28144 6 io_out[21]
port 193 nsew signal output
rlabel metal3 s 39200 28840 40000 28960 6 io_out[22]
port 194 nsew signal output
rlabel metal3 s 39200 29656 40000 29776 6 io_out[23]
port 195 nsew signal output
rlabel metal3 s 39200 30472 40000 30592 6 io_out[24]
port 196 nsew signal output
rlabel metal3 s 39200 31288 40000 31408 6 io_out[25]
port 197 nsew signal output
rlabel metal3 s 39200 32104 40000 32224 6 io_out[26]
port 198 nsew signal output
rlabel metal3 s 39200 32920 40000 33040 6 io_out[27]
port 199 nsew signal output
rlabel metal3 s 39200 33736 40000 33856 6 io_out[28]
port 200 nsew signal output
rlabel metal3 s 39200 34552 40000 34672 6 io_out[29]
port 201 nsew signal output
rlabel metal3 s 39200 12520 40000 12640 6 io_out[2]
port 202 nsew signal output
rlabel metal3 s 39200 35368 40000 35488 6 io_out[30]
port 203 nsew signal output
rlabel metal3 s 39200 36184 40000 36304 6 io_out[31]
port 204 nsew signal output
rlabel metal3 s 39200 37000 40000 37120 6 io_out[32]
port 205 nsew signal output
rlabel metal3 s 39200 37816 40000 37936 6 io_out[33]
port 206 nsew signal output
rlabel metal3 s 39200 38632 40000 38752 6 io_out[34]
port 207 nsew signal output
rlabel metal3 s 39200 39448 40000 39568 6 io_out[35]
port 208 nsew signal output
rlabel metal3 s 39200 40264 40000 40384 6 io_out[36]
port 209 nsew signal output
rlabel metal3 s 39200 41080 40000 41200 6 io_out[37]
port 210 nsew signal output
rlabel metal3 s 39200 13336 40000 13456 6 io_out[3]
port 211 nsew signal output
rlabel metal3 s 39200 14152 40000 14272 6 io_out[4]
port 212 nsew signal output
rlabel metal3 s 39200 14968 40000 15088 6 io_out[5]
port 213 nsew signal output
rlabel metal3 s 39200 15784 40000 15904 6 io_out[6]
port 214 nsew signal output
rlabel metal3 s 39200 16600 40000 16720 6 io_out[7]
port 215 nsew signal output
rlabel metal3 s 39200 17416 40000 17536 6 io_out[8]
port 216 nsew signal output
rlabel metal3 s 39200 18232 40000 18352 6 io_out[9]
port 217 nsew signal output
rlabel metal3 s 39200 160216 40000 160336 6 io_out_scrapcpu[0]
port 218 nsew signal input
rlabel metal3 s 39200 168376 40000 168496 6 io_out_scrapcpu[10]
port 219 nsew signal input
rlabel metal3 s 39200 169192 40000 169312 6 io_out_scrapcpu[11]
port 220 nsew signal input
rlabel metal3 s 39200 170008 40000 170128 6 io_out_scrapcpu[12]
port 221 nsew signal input
rlabel metal3 s 39200 170824 40000 170944 6 io_out_scrapcpu[13]
port 222 nsew signal input
rlabel metal3 s 39200 171640 40000 171760 6 io_out_scrapcpu[14]
port 223 nsew signal input
rlabel metal3 s 39200 172456 40000 172576 6 io_out_scrapcpu[15]
port 224 nsew signal input
rlabel metal3 s 39200 173272 40000 173392 6 io_out_scrapcpu[16]
port 225 nsew signal input
rlabel metal3 s 39200 174088 40000 174208 6 io_out_scrapcpu[17]
port 226 nsew signal input
rlabel metal3 s 39200 174904 40000 175024 6 io_out_scrapcpu[18]
port 227 nsew signal input
rlabel metal3 s 39200 175720 40000 175840 6 io_out_scrapcpu[19]
port 228 nsew signal input
rlabel metal3 s 39200 161032 40000 161152 6 io_out_scrapcpu[1]
port 229 nsew signal input
rlabel metal3 s 39200 176536 40000 176656 6 io_out_scrapcpu[20]
port 230 nsew signal input
rlabel metal3 s 39200 177352 40000 177472 6 io_out_scrapcpu[21]
port 231 nsew signal input
rlabel metal3 s 39200 178168 40000 178288 6 io_out_scrapcpu[22]
port 232 nsew signal input
rlabel metal3 s 39200 178984 40000 179104 6 io_out_scrapcpu[23]
port 233 nsew signal input
rlabel metal3 s 39200 179800 40000 179920 6 io_out_scrapcpu[24]
port 234 nsew signal input
rlabel metal3 s 39200 180616 40000 180736 6 io_out_scrapcpu[25]
port 235 nsew signal input
rlabel metal3 s 39200 181432 40000 181552 6 io_out_scrapcpu[26]
port 236 nsew signal input
rlabel metal3 s 39200 182248 40000 182368 6 io_out_scrapcpu[27]
port 237 nsew signal input
rlabel metal3 s 39200 183064 40000 183184 6 io_out_scrapcpu[28]
port 238 nsew signal input
rlabel metal3 s 39200 183880 40000 184000 6 io_out_scrapcpu[29]
port 239 nsew signal input
rlabel metal3 s 39200 161848 40000 161968 6 io_out_scrapcpu[2]
port 240 nsew signal input
rlabel metal3 s 39200 184696 40000 184816 6 io_out_scrapcpu[30]
port 241 nsew signal input
rlabel metal3 s 39200 185512 40000 185632 6 io_out_scrapcpu[31]
port 242 nsew signal input
rlabel metal3 s 39200 186328 40000 186448 6 io_out_scrapcpu[32]
port 243 nsew signal input
rlabel metal3 s 39200 187144 40000 187264 6 io_out_scrapcpu[33]
port 244 nsew signal input
rlabel metal3 s 39200 187960 40000 188080 6 io_out_scrapcpu[34]
port 245 nsew signal input
rlabel metal3 s 39200 188776 40000 188896 6 io_out_scrapcpu[35]
port 246 nsew signal input
rlabel metal3 s 39200 162664 40000 162784 6 io_out_scrapcpu[3]
port 247 nsew signal input
rlabel metal3 s 39200 163480 40000 163600 6 io_out_scrapcpu[4]
port 248 nsew signal input
rlabel metal3 s 39200 164296 40000 164416 6 io_out_scrapcpu[5]
port 249 nsew signal input
rlabel metal3 s 39200 165112 40000 165232 6 io_out_scrapcpu[6]
port 250 nsew signal input
rlabel metal3 s 39200 165928 40000 166048 6 io_out_scrapcpu[7]
port 251 nsew signal input
rlabel metal3 s 39200 166744 40000 166864 6 io_out_scrapcpu[8]
port 252 nsew signal input
rlabel metal3 s 39200 167560 40000 167680 6 io_out_scrapcpu[9]
port 253 nsew signal input
rlabel metal2 s 2778 199200 2834 200000 6 io_out_vliw[0]
port 254 nsew signal input
rlabel metal2 s 12898 199200 12954 200000 6 io_out_vliw[10]
port 255 nsew signal input
rlabel metal2 s 13910 199200 13966 200000 6 io_out_vliw[11]
port 256 nsew signal input
rlabel metal2 s 14922 199200 14978 200000 6 io_out_vliw[12]
port 257 nsew signal input
rlabel metal2 s 15934 199200 15990 200000 6 io_out_vliw[13]
port 258 nsew signal input
rlabel metal2 s 16946 199200 17002 200000 6 io_out_vliw[14]
port 259 nsew signal input
rlabel metal2 s 17958 199200 18014 200000 6 io_out_vliw[15]
port 260 nsew signal input
rlabel metal2 s 18970 199200 19026 200000 6 io_out_vliw[16]
port 261 nsew signal input
rlabel metal2 s 19982 199200 20038 200000 6 io_out_vliw[17]
port 262 nsew signal input
rlabel metal2 s 20994 199200 21050 200000 6 io_out_vliw[18]
port 263 nsew signal input
rlabel metal2 s 22006 199200 22062 200000 6 io_out_vliw[19]
port 264 nsew signal input
rlabel metal2 s 3790 199200 3846 200000 6 io_out_vliw[1]
port 265 nsew signal input
rlabel metal2 s 23018 199200 23074 200000 6 io_out_vliw[20]
port 266 nsew signal input
rlabel metal2 s 24030 199200 24086 200000 6 io_out_vliw[21]
port 267 nsew signal input
rlabel metal2 s 25042 199200 25098 200000 6 io_out_vliw[22]
port 268 nsew signal input
rlabel metal2 s 26054 199200 26110 200000 6 io_out_vliw[23]
port 269 nsew signal input
rlabel metal2 s 27066 199200 27122 200000 6 io_out_vliw[24]
port 270 nsew signal input
rlabel metal2 s 28078 199200 28134 200000 6 io_out_vliw[25]
port 271 nsew signal input
rlabel metal2 s 29090 199200 29146 200000 6 io_out_vliw[26]
port 272 nsew signal input
rlabel metal2 s 30102 199200 30158 200000 6 io_out_vliw[27]
port 273 nsew signal input
rlabel metal2 s 31114 199200 31170 200000 6 io_out_vliw[28]
port 274 nsew signal input
rlabel metal2 s 32126 199200 32182 200000 6 io_out_vliw[29]
port 275 nsew signal input
rlabel metal2 s 4802 199200 4858 200000 6 io_out_vliw[2]
port 276 nsew signal input
rlabel metal2 s 33138 199200 33194 200000 6 io_out_vliw[30]
port 277 nsew signal input
rlabel metal2 s 34150 199200 34206 200000 6 io_out_vliw[31]
port 278 nsew signal input
rlabel metal2 s 35162 199200 35218 200000 6 io_out_vliw[32]
port 279 nsew signal input
rlabel metal2 s 36174 199200 36230 200000 6 io_out_vliw[33]
port 280 nsew signal input
rlabel metal2 s 37186 199200 37242 200000 6 io_out_vliw[34]
port 281 nsew signal input
rlabel metal2 s 38198 199200 38254 200000 6 io_out_vliw[35]
port 282 nsew signal input
rlabel metal2 s 5814 199200 5870 200000 6 io_out_vliw[3]
port 283 nsew signal input
rlabel metal2 s 6826 199200 6882 200000 6 io_out_vliw[4]
port 284 nsew signal input
rlabel metal2 s 7838 199200 7894 200000 6 io_out_vliw[5]
port 285 nsew signal input
rlabel metal2 s 8850 199200 8906 200000 6 io_out_vliw[6]
port 286 nsew signal input
rlabel metal2 s 9862 199200 9918 200000 6 io_out_vliw[7]
port 287 nsew signal input
rlabel metal2 s 10874 199200 10930 200000 6 io_out_vliw[8]
port 288 nsew signal input
rlabel metal2 s 11886 199200 11942 200000 6 io_out_vliw[9]
port 289 nsew signal input
rlabel metal3 s 39200 100648 40000 100768 6 io_out_z80[0]
port 290 nsew signal input
rlabel metal3 s 39200 108808 40000 108928 6 io_out_z80[10]
port 291 nsew signal input
rlabel metal3 s 39200 109624 40000 109744 6 io_out_z80[11]
port 292 nsew signal input
rlabel metal3 s 39200 110440 40000 110560 6 io_out_z80[12]
port 293 nsew signal input
rlabel metal3 s 39200 111256 40000 111376 6 io_out_z80[13]
port 294 nsew signal input
rlabel metal3 s 39200 112072 40000 112192 6 io_out_z80[14]
port 295 nsew signal input
rlabel metal3 s 39200 112888 40000 113008 6 io_out_z80[15]
port 296 nsew signal input
rlabel metal3 s 39200 113704 40000 113824 6 io_out_z80[16]
port 297 nsew signal input
rlabel metal3 s 39200 114520 40000 114640 6 io_out_z80[17]
port 298 nsew signal input
rlabel metal3 s 39200 115336 40000 115456 6 io_out_z80[18]
port 299 nsew signal input
rlabel metal3 s 39200 116152 40000 116272 6 io_out_z80[19]
port 300 nsew signal input
rlabel metal3 s 39200 101464 40000 101584 6 io_out_z80[1]
port 301 nsew signal input
rlabel metal3 s 39200 116968 40000 117088 6 io_out_z80[20]
port 302 nsew signal input
rlabel metal3 s 39200 117784 40000 117904 6 io_out_z80[21]
port 303 nsew signal input
rlabel metal3 s 39200 118600 40000 118720 6 io_out_z80[22]
port 304 nsew signal input
rlabel metal3 s 39200 119416 40000 119536 6 io_out_z80[23]
port 305 nsew signal input
rlabel metal3 s 39200 120232 40000 120352 6 io_out_z80[24]
port 306 nsew signal input
rlabel metal3 s 39200 121048 40000 121168 6 io_out_z80[25]
port 307 nsew signal input
rlabel metal3 s 39200 121864 40000 121984 6 io_out_z80[26]
port 308 nsew signal input
rlabel metal3 s 39200 122680 40000 122800 6 io_out_z80[27]
port 309 nsew signal input
rlabel metal3 s 39200 123496 40000 123616 6 io_out_z80[28]
port 310 nsew signal input
rlabel metal3 s 39200 124312 40000 124432 6 io_out_z80[29]
port 311 nsew signal input
rlabel metal3 s 39200 102280 40000 102400 6 io_out_z80[2]
port 312 nsew signal input
rlabel metal3 s 39200 125128 40000 125248 6 io_out_z80[30]
port 313 nsew signal input
rlabel metal3 s 39200 125944 40000 126064 6 io_out_z80[31]
port 314 nsew signal input
rlabel metal3 s 39200 126760 40000 126880 6 io_out_z80[32]
port 315 nsew signal input
rlabel metal3 s 39200 127576 40000 127696 6 io_out_z80[33]
port 316 nsew signal input
rlabel metal3 s 39200 128392 40000 128512 6 io_out_z80[34]
port 317 nsew signal input
rlabel metal3 s 39200 129208 40000 129328 6 io_out_z80[35]
port 318 nsew signal input
rlabel metal3 s 39200 103096 40000 103216 6 io_out_z80[3]
port 319 nsew signal input
rlabel metal3 s 39200 103912 40000 104032 6 io_out_z80[4]
port 320 nsew signal input
rlabel metal3 s 39200 104728 40000 104848 6 io_out_z80[5]
port 321 nsew signal input
rlabel metal3 s 39200 105544 40000 105664 6 io_out_z80[6]
port 322 nsew signal input
rlabel metal3 s 39200 106360 40000 106480 6 io_out_z80[7]
port 323 nsew signal input
rlabel metal3 s 39200 107176 40000 107296 6 io_out_z80[8]
port 324 nsew signal input
rlabel metal3 s 39200 107992 40000 108112 6 io_out_z80[9]
port 325 nsew signal input
rlabel metal3 s 39200 68008 40000 68128 6 la_data_out[0]
port 326 nsew signal output
rlabel metal3 s 39200 76168 40000 76288 6 la_data_out[10]
port 327 nsew signal output
rlabel metal3 s 39200 76984 40000 77104 6 la_data_out[11]
port 328 nsew signal output
rlabel metal3 s 39200 77800 40000 77920 6 la_data_out[12]
port 329 nsew signal output
rlabel metal3 s 39200 78616 40000 78736 6 la_data_out[13]
port 330 nsew signal output
rlabel metal3 s 39200 79432 40000 79552 6 la_data_out[14]
port 331 nsew signal output
rlabel metal3 s 39200 80248 40000 80368 6 la_data_out[15]
port 332 nsew signal output
rlabel metal3 s 39200 81064 40000 81184 6 la_data_out[16]
port 333 nsew signal output
rlabel metal3 s 39200 81880 40000 82000 6 la_data_out[17]
port 334 nsew signal output
rlabel metal3 s 39200 82696 40000 82816 6 la_data_out[18]
port 335 nsew signal output
rlabel metal3 s 39200 83512 40000 83632 6 la_data_out[19]
port 336 nsew signal output
rlabel metal3 s 39200 68824 40000 68944 6 la_data_out[1]
port 337 nsew signal output
rlabel metal3 s 39200 84328 40000 84448 6 la_data_out[20]
port 338 nsew signal output
rlabel metal3 s 39200 85144 40000 85264 6 la_data_out[21]
port 339 nsew signal output
rlabel metal3 s 39200 85960 40000 86080 6 la_data_out[22]
port 340 nsew signal output
rlabel metal3 s 39200 86776 40000 86896 6 la_data_out[23]
port 341 nsew signal output
rlabel metal3 s 39200 87592 40000 87712 6 la_data_out[24]
port 342 nsew signal output
rlabel metal3 s 39200 88408 40000 88528 6 la_data_out[25]
port 343 nsew signal output
rlabel metal3 s 39200 89224 40000 89344 6 la_data_out[26]
port 344 nsew signal output
rlabel metal3 s 39200 90040 40000 90160 6 la_data_out[27]
port 345 nsew signal output
rlabel metal3 s 39200 90856 40000 90976 6 la_data_out[28]
port 346 nsew signal output
rlabel metal3 s 39200 91672 40000 91792 6 la_data_out[29]
port 347 nsew signal output
rlabel metal3 s 39200 69640 40000 69760 6 la_data_out[2]
port 348 nsew signal output
rlabel metal3 s 39200 92488 40000 92608 6 la_data_out[30]
port 349 nsew signal output
rlabel metal3 s 39200 93304 40000 93424 6 la_data_out[31]
port 350 nsew signal output
rlabel metal3 s 39200 94120 40000 94240 6 la_data_out[32]
port 351 nsew signal output
rlabel metal3 s 39200 94936 40000 95056 6 la_data_out[33]
port 352 nsew signal output
rlabel metal3 s 39200 95752 40000 95872 6 la_data_out[34]
port 353 nsew signal output
rlabel metal3 s 39200 96568 40000 96688 6 la_data_out[35]
port 354 nsew signal output
rlabel metal3 s 39200 97384 40000 97504 6 la_data_out[36]
port 355 nsew signal output
rlabel metal3 s 39200 98200 40000 98320 6 la_data_out[37]
port 356 nsew signal output
rlabel metal3 s 39200 99016 40000 99136 6 la_data_out[38]
port 357 nsew signal output
rlabel metal3 s 39200 99832 40000 99952 6 la_data_out[39]
port 358 nsew signal output
rlabel metal3 s 39200 70456 40000 70576 6 la_data_out[3]
port 359 nsew signal output
rlabel metal3 s 39200 71272 40000 71392 6 la_data_out[4]
port 360 nsew signal output
rlabel metal3 s 39200 72088 40000 72208 6 la_data_out[5]
port 361 nsew signal output
rlabel metal3 s 39200 72904 40000 73024 6 la_data_out[6]
port 362 nsew signal output
rlabel metal3 s 39200 73720 40000 73840 6 la_data_out[7]
port 363 nsew signal output
rlabel metal3 s 39200 74536 40000 74656 6 la_data_out[8]
port 364 nsew signal output
rlabel metal3 s 39200 75352 40000 75472 6 la_data_out[9]
port 365 nsew signal output
rlabel metal2 s 39210 199200 39266 200000 6 rst_scrapcpu
port 366 nsew signal output
rlabel metal2 s 1766 199200 1822 200000 6 rst_vliw
port 367 nsew signal output
rlabel metal3 s 39200 130024 40000 130144 6 rst_z80
port 368 nsew signal output
rlabel metal4 s 4208 2128 4528 197520 6 vccd1
port 369 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 197520 6 vccd1
port 369 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 197520 6 vssd1
port 370 nsew ground bidirectional
rlabel metal3 s 0 78616 800 78736 6 wb_clk_i
port 371 nsew signal input
rlabel metal3 s 0 79704 800 79824 6 wb_rst_i
port 372 nsew signal input
rlabel metal3 s 0 118872 800 118992 6 wbs_ack_o
port 373 nsew signal output
rlabel metal2 s 1398 0 1454 800 6 wbs_adr_i[0]
port 374 nsew signal input
rlabel metal2 s 13358 0 13414 800 6 wbs_adr_i[10]
port 375 nsew signal input
rlabel metal2 s 14554 0 14610 800 6 wbs_adr_i[11]
port 376 nsew signal input
rlabel metal2 s 15750 0 15806 800 6 wbs_adr_i[12]
port 377 nsew signal input
rlabel metal2 s 16946 0 17002 800 6 wbs_adr_i[13]
port 378 nsew signal input
rlabel metal2 s 18142 0 18198 800 6 wbs_adr_i[14]
port 379 nsew signal input
rlabel metal2 s 19338 0 19394 800 6 wbs_adr_i[15]
port 380 nsew signal input
rlabel metal2 s 20534 0 20590 800 6 wbs_adr_i[16]
port 381 nsew signal input
rlabel metal2 s 21730 0 21786 800 6 wbs_adr_i[17]
port 382 nsew signal input
rlabel metal2 s 22926 0 22982 800 6 wbs_adr_i[18]
port 383 nsew signal input
rlabel metal2 s 24122 0 24178 800 6 wbs_adr_i[19]
port 384 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 wbs_adr_i[1]
port 385 nsew signal input
rlabel metal2 s 25318 0 25374 800 6 wbs_adr_i[20]
port 386 nsew signal input
rlabel metal2 s 26514 0 26570 800 6 wbs_adr_i[21]
port 387 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 wbs_adr_i[22]
port 388 nsew signal input
rlabel metal2 s 28906 0 28962 800 6 wbs_adr_i[23]
port 389 nsew signal input
rlabel metal2 s 30102 0 30158 800 6 wbs_adr_i[24]
port 390 nsew signal input
rlabel metal2 s 31298 0 31354 800 6 wbs_adr_i[25]
port 391 nsew signal input
rlabel metal2 s 32494 0 32550 800 6 wbs_adr_i[26]
port 392 nsew signal input
rlabel metal2 s 33690 0 33746 800 6 wbs_adr_i[27]
port 393 nsew signal input
rlabel metal2 s 34886 0 34942 800 6 wbs_adr_i[28]
port 394 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 wbs_adr_i[29]
port 395 nsew signal input
rlabel metal2 s 3790 0 3846 800 6 wbs_adr_i[2]
port 396 nsew signal input
rlabel metal2 s 37278 0 37334 800 6 wbs_adr_i[30]
port 397 nsew signal input
rlabel metal2 s 38474 0 38530 800 6 wbs_adr_i[31]
port 398 nsew signal input
rlabel metal2 s 4986 0 5042 800 6 wbs_adr_i[3]
port 399 nsew signal input
rlabel metal2 s 6182 0 6238 800 6 wbs_adr_i[4]
port 400 nsew signal input
rlabel metal2 s 7378 0 7434 800 6 wbs_adr_i[5]
port 401 nsew signal input
rlabel metal2 s 8574 0 8630 800 6 wbs_adr_i[6]
port 402 nsew signal input
rlabel metal2 s 9770 0 9826 800 6 wbs_adr_i[7]
port 403 nsew signal input
rlabel metal2 s 10966 0 11022 800 6 wbs_adr_i[8]
port 404 nsew signal input
rlabel metal2 s 12162 0 12218 800 6 wbs_adr_i[9]
port 405 nsew signal input
rlabel metal3 s 0 116696 800 116816 6 wbs_cyc_i
port 406 nsew signal input
rlabel metal3 s 0 80792 800 80912 6 wbs_dat_i[0]
port 407 nsew signal input
rlabel metal3 s 0 91672 800 91792 6 wbs_dat_i[10]
port 408 nsew signal input
rlabel metal3 s 0 92760 800 92880 6 wbs_dat_i[11]
port 409 nsew signal input
rlabel metal3 s 0 93848 800 93968 6 wbs_dat_i[12]
port 410 nsew signal input
rlabel metal3 s 0 94936 800 95056 6 wbs_dat_i[13]
port 411 nsew signal input
rlabel metal3 s 0 96024 800 96144 6 wbs_dat_i[14]
port 412 nsew signal input
rlabel metal3 s 0 97112 800 97232 6 wbs_dat_i[15]
port 413 nsew signal input
rlabel metal3 s 0 98200 800 98320 6 wbs_dat_i[16]
port 414 nsew signal input
rlabel metal3 s 0 99288 800 99408 6 wbs_dat_i[17]
port 415 nsew signal input
rlabel metal3 s 0 100376 800 100496 6 wbs_dat_i[18]
port 416 nsew signal input
rlabel metal3 s 0 101464 800 101584 6 wbs_dat_i[19]
port 417 nsew signal input
rlabel metal3 s 0 81880 800 82000 6 wbs_dat_i[1]
port 418 nsew signal input
rlabel metal3 s 0 102552 800 102672 6 wbs_dat_i[20]
port 419 nsew signal input
rlabel metal3 s 0 103640 800 103760 6 wbs_dat_i[21]
port 420 nsew signal input
rlabel metal3 s 0 104728 800 104848 6 wbs_dat_i[22]
port 421 nsew signal input
rlabel metal3 s 0 105816 800 105936 6 wbs_dat_i[23]
port 422 nsew signal input
rlabel metal3 s 0 106904 800 107024 6 wbs_dat_i[24]
port 423 nsew signal input
rlabel metal3 s 0 107992 800 108112 6 wbs_dat_i[25]
port 424 nsew signal input
rlabel metal3 s 0 109080 800 109200 6 wbs_dat_i[26]
port 425 nsew signal input
rlabel metal3 s 0 110168 800 110288 6 wbs_dat_i[27]
port 426 nsew signal input
rlabel metal3 s 0 111256 800 111376 6 wbs_dat_i[28]
port 427 nsew signal input
rlabel metal3 s 0 112344 800 112464 6 wbs_dat_i[29]
port 428 nsew signal input
rlabel metal3 s 0 82968 800 83088 6 wbs_dat_i[2]
port 429 nsew signal input
rlabel metal3 s 0 113432 800 113552 6 wbs_dat_i[30]
port 430 nsew signal input
rlabel metal3 s 0 114520 800 114640 6 wbs_dat_i[31]
port 431 nsew signal input
rlabel metal3 s 0 84056 800 84176 6 wbs_dat_i[3]
port 432 nsew signal input
rlabel metal3 s 0 85144 800 85264 6 wbs_dat_i[4]
port 433 nsew signal input
rlabel metal3 s 0 86232 800 86352 6 wbs_dat_i[5]
port 434 nsew signal input
rlabel metal3 s 0 87320 800 87440 6 wbs_dat_i[6]
port 435 nsew signal input
rlabel metal3 s 0 88408 800 88528 6 wbs_dat_i[7]
port 436 nsew signal input
rlabel metal3 s 0 89496 800 89616 6 wbs_dat_i[8]
port 437 nsew signal input
rlabel metal3 s 0 90584 800 90704 6 wbs_dat_i[9]
port 438 nsew signal input
rlabel metal3 s 39200 41896 40000 42016 6 wbs_dat_o[0]
port 439 nsew signal output
rlabel metal3 s 39200 50056 40000 50176 6 wbs_dat_o[10]
port 440 nsew signal output
rlabel metal3 s 39200 50872 40000 50992 6 wbs_dat_o[11]
port 441 nsew signal output
rlabel metal3 s 39200 51688 40000 51808 6 wbs_dat_o[12]
port 442 nsew signal output
rlabel metal3 s 39200 52504 40000 52624 6 wbs_dat_o[13]
port 443 nsew signal output
rlabel metal3 s 39200 53320 40000 53440 6 wbs_dat_o[14]
port 444 nsew signal output
rlabel metal3 s 39200 54136 40000 54256 6 wbs_dat_o[15]
port 445 nsew signal output
rlabel metal3 s 39200 54952 40000 55072 6 wbs_dat_o[16]
port 446 nsew signal output
rlabel metal3 s 39200 55768 40000 55888 6 wbs_dat_o[17]
port 447 nsew signal output
rlabel metal3 s 39200 56584 40000 56704 6 wbs_dat_o[18]
port 448 nsew signal output
rlabel metal3 s 39200 57400 40000 57520 6 wbs_dat_o[19]
port 449 nsew signal output
rlabel metal3 s 39200 42712 40000 42832 6 wbs_dat_o[1]
port 450 nsew signal output
rlabel metal3 s 39200 58216 40000 58336 6 wbs_dat_o[20]
port 451 nsew signal output
rlabel metal3 s 39200 59032 40000 59152 6 wbs_dat_o[21]
port 452 nsew signal output
rlabel metal3 s 39200 59848 40000 59968 6 wbs_dat_o[22]
port 453 nsew signal output
rlabel metal3 s 39200 60664 40000 60784 6 wbs_dat_o[23]
port 454 nsew signal output
rlabel metal3 s 39200 61480 40000 61600 6 wbs_dat_o[24]
port 455 nsew signal output
rlabel metal3 s 39200 62296 40000 62416 6 wbs_dat_o[25]
port 456 nsew signal output
rlabel metal3 s 39200 63112 40000 63232 6 wbs_dat_o[26]
port 457 nsew signal output
rlabel metal3 s 39200 63928 40000 64048 6 wbs_dat_o[27]
port 458 nsew signal output
rlabel metal3 s 39200 64744 40000 64864 6 wbs_dat_o[28]
port 459 nsew signal output
rlabel metal3 s 39200 65560 40000 65680 6 wbs_dat_o[29]
port 460 nsew signal output
rlabel metal3 s 39200 43528 40000 43648 6 wbs_dat_o[2]
port 461 nsew signal output
rlabel metal3 s 39200 66376 40000 66496 6 wbs_dat_o[30]
port 462 nsew signal output
rlabel metal3 s 39200 67192 40000 67312 6 wbs_dat_o[31]
port 463 nsew signal output
rlabel metal3 s 39200 44344 40000 44464 6 wbs_dat_o[3]
port 464 nsew signal output
rlabel metal3 s 39200 45160 40000 45280 6 wbs_dat_o[4]
port 465 nsew signal output
rlabel metal3 s 39200 45976 40000 46096 6 wbs_dat_o[5]
port 466 nsew signal output
rlabel metal3 s 39200 46792 40000 46912 6 wbs_dat_o[6]
port 467 nsew signal output
rlabel metal3 s 39200 47608 40000 47728 6 wbs_dat_o[7]
port 468 nsew signal output
rlabel metal3 s 39200 48424 40000 48544 6 wbs_dat_o[8]
port 469 nsew signal output
rlabel metal3 s 39200 49240 40000 49360 6 wbs_dat_o[9]
port 470 nsew signal output
rlabel metal3 s 0 117784 800 117904 6 wbs_stb_i
port 471 nsew signal input
rlabel metal3 s 0 115608 800 115728 6 wbs_we_i
port 472 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 40000 200000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 6687402
string GDS_FILE /home/tholin/Desktop/ci2406-rej-pommedeterrible-tholin/openlane/Multiplexer/runs/24_05_31_21_33/results/signoff/multiplexer.magic.gds
string GDS_START 373516
<< end >>

