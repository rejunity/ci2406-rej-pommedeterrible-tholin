// This is the unpowered netlist.
module wrapped_6502 (io_oeb,
    rst_n,
    wb_clk_i,
    custom_settings,
    io_in,
    io_out);
 output io_oeb;
 input rst_n;
 input wb_clk_i;
 input [1:0] custom_settings;
 input [35:0] io_in;
 output [35:0] io_out;

 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire \MOS6502.ABH[0] ;
 wire \MOS6502.ABH[1] ;
 wire \MOS6502.ABH[2] ;
 wire \MOS6502.ABH[3] ;
 wire \MOS6502.ABH[4] ;
 wire \MOS6502.ABH[5] ;
 wire \MOS6502.ABH[6] ;
 wire \MOS6502.ABH[7] ;
 wire \MOS6502.ABL[0] ;
 wire \MOS6502.ABL[1] ;
 wire \MOS6502.ABL[2] ;
 wire \MOS6502.ABL[3] ;
 wire \MOS6502.ABL[4] ;
 wire \MOS6502.ABL[5] ;
 wire \MOS6502.ABL[6] ;
 wire \MOS6502.ABL[7] ;
 wire \MOS6502.ADD[0] ;
 wire \MOS6502.ADD[1] ;
 wire \MOS6502.ADD[2] ;
 wire \MOS6502.ADD[3] ;
 wire \MOS6502.ADD[4] ;
 wire \MOS6502.ADD[5] ;
 wire \MOS6502.ADD[6] ;
 wire \MOS6502.ADD[7] ;
 wire \MOS6502.ALU.AI7 ;
 wire \MOS6502.ALU.BI7 ;
 wire \MOS6502.ALU.CO ;
 wire \MOS6502.ALU.HC ;
 wire \MOS6502.AXYS[0][0] ;
 wire \MOS6502.AXYS[0][1] ;
 wire \MOS6502.AXYS[0][2] ;
 wire \MOS6502.AXYS[0][3] ;
 wire \MOS6502.AXYS[0][4] ;
 wire \MOS6502.AXYS[0][5] ;
 wire \MOS6502.AXYS[0][6] ;
 wire \MOS6502.AXYS[0][7] ;
 wire \MOS6502.AXYS[1][0] ;
 wire \MOS6502.AXYS[1][1] ;
 wire \MOS6502.AXYS[1][2] ;
 wire \MOS6502.AXYS[1][3] ;
 wire \MOS6502.AXYS[1][4] ;
 wire \MOS6502.AXYS[1][5] ;
 wire \MOS6502.AXYS[1][6] ;
 wire \MOS6502.AXYS[1][7] ;
 wire \MOS6502.AXYS[2][0] ;
 wire \MOS6502.AXYS[2][1] ;
 wire \MOS6502.AXYS[2][2] ;
 wire \MOS6502.AXYS[2][3] ;
 wire \MOS6502.AXYS[2][4] ;
 wire \MOS6502.AXYS[2][5] ;
 wire \MOS6502.AXYS[2][6] ;
 wire \MOS6502.AXYS[2][7] ;
 wire \MOS6502.AXYS[3][0] ;
 wire \MOS6502.AXYS[3][1] ;
 wire \MOS6502.AXYS[3][2] ;
 wire \MOS6502.AXYS[3][3] ;
 wire \MOS6502.AXYS[3][4] ;
 wire \MOS6502.AXYS[3][5] ;
 wire \MOS6502.AXYS[3][6] ;
 wire \MOS6502.AXYS[3][7] ;
 wire \MOS6502.DIHOLD[0] ;
 wire \MOS6502.DIHOLD[1] ;
 wire \MOS6502.DIHOLD[2] ;
 wire \MOS6502.DIHOLD[3] ;
 wire \MOS6502.DIHOLD[4] ;
 wire \MOS6502.DIHOLD[5] ;
 wire \MOS6502.DIHOLD[6] ;
 wire \MOS6502.DIHOLD[7] ;
 wire \MOS6502.DI[0] ;
 wire \MOS6502.DI[1] ;
 wire \MOS6502.DI[2] ;
 wire \MOS6502.DI[3] ;
 wire \MOS6502.DI[4] ;
 wire \MOS6502.DI[5] ;
 wire \MOS6502.DI[6] ;
 wire \MOS6502.DI[7] ;
 wire \MOS6502.IRHOLD[0] ;
 wire \MOS6502.IRHOLD[1] ;
 wire \MOS6502.IRHOLD[2] ;
 wire \MOS6502.IRHOLD[3] ;
 wire \MOS6502.IRHOLD[4] ;
 wire \MOS6502.IRHOLD[5] ;
 wire \MOS6502.IRHOLD[6] ;
 wire \MOS6502.IRHOLD[7] ;
 wire \MOS6502.IRHOLD_valid ;
 wire \MOS6502.NMI_1 ;
 wire \MOS6502.NMI_edge ;
 wire \MOS6502.PC[0] ;
 wire \MOS6502.PC[10] ;
 wire \MOS6502.PC[11] ;
 wire \MOS6502.PC[12] ;
 wire \MOS6502.PC[13] ;
 wire \MOS6502.PC[14] ;
 wire \MOS6502.PC[15] ;
 wire \MOS6502.PC[1] ;
 wire \MOS6502.PC[2] ;
 wire \MOS6502.PC[3] ;
 wire \MOS6502.PC[4] ;
 wire \MOS6502.PC[5] ;
 wire \MOS6502.PC[6] ;
 wire \MOS6502.PC[7] ;
 wire \MOS6502.PC[8] ;
 wire \MOS6502.PC[9] ;
 wire \MOS6502.adc_bcd ;
 wire \MOS6502.adc_sbc ;
 wire \MOS6502.adj_bcd ;
 wire \MOS6502.backwards ;
 wire \MOS6502.bit_ins ;
 wire \MOS6502.clc ;
 wire \MOS6502.cld ;
 wire \MOS6502.cli ;
 wire \MOS6502.clv ;
 wire \MOS6502.compare ;
 wire \MOS6502.cond_code[0] ;
 wire \MOS6502.cond_code[1] ;
 wire \MOS6502.cond_code[2] ;
 wire \MOS6502.dst_reg[0] ;
 wire \MOS6502.dst_reg[1] ;
 wire \MOS6502.inc ;
 wire \MOS6502.index_y ;
 wire \MOS6502.load_only ;
 wire \MOS6502.load_reg ;
 wire \MOS6502.op[0] ;
 wire \MOS6502.op[1] ;
 wire \MOS6502.op[2] ;
 wire \MOS6502.op[3] ;
 wire \MOS6502.php ;
 wire \MOS6502.plp ;
 wire \MOS6502.res ;
 wire \MOS6502.rotate ;
 wire \MOS6502.sec ;
 wire \MOS6502.sed ;
 wire \MOS6502.sei ;
 wire \MOS6502.shift ;
 wire \MOS6502.shift_right ;
 wire \MOS6502.src_reg[0] ;
 wire \MOS6502.src_reg[1] ;
 wire \MOS6502.state[0] ;
 wire \MOS6502.state[1] ;
 wire \MOS6502.state[2] ;
 wire \MOS6502.state[3] ;
 wire \MOS6502.state[4] ;
 wire \MOS6502.state[5] ;
 wire \MOS6502.store ;
 wire \MOS6502.write_back ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire clknet_0_wb_clk_i;
 wire clknet_4_0_0_wb_clk_i;
 wire clknet_4_10_0_wb_clk_i;
 wire clknet_4_11_0_wb_clk_i;
 wire clknet_4_12_0_wb_clk_i;
 wire clknet_4_13_0_wb_clk_i;
 wire clknet_4_14_0_wb_clk_i;
 wire clknet_4_15_0_wb_clk_i;
 wire clknet_4_1_0_wb_clk_i;
 wire clknet_4_2_0_wb_clk_i;
 wire clknet_4_3_0_wb_clk_i;
 wire clknet_4_4_0_wb_clk_i;
 wire clknet_4_5_0_wb_clk_i;
 wire clknet_4_6_0_wb_clk_i;
 wire clknet_4_7_0_wb_clk_i;
 wire clknet_4_8_0_wb_clk_i;
 wire clknet_4_9_0_wb_clk_i;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__1026__A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__1039__A (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__1053__A (.DIODE(_0451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1054__B (.DIODE(_0451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1075__D (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__1087__A2 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__1088__A2 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__1090__B (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__1129__A (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__1132__A (.DIODE(_0534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1135__A (.DIODE(_0534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1146__S (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__1147__B2 (.DIODE(_0549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1148__B2 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__1156__S (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__1157__B2 (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1163__S (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__1164__B2 (.DIODE(_0564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1170__S (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__1171__B2 (.DIODE(_0570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1178__S (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__1179__B2 (.DIODE(_0577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1187__S (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__1188__B2 (.DIODE(_0585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1189__A1 (.DIODE(\MOS6502.ADD[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1194__S (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__1195__B2 (.DIODE(_0591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1203__S (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__1204__B2 (.DIODE(_0599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1208__A2 (.DIODE(_0549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1209__A1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__1210__A2 (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1212__A2 (.DIODE(_0564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1214__A2 (.DIODE(_0570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1216__A2 (.DIODE(_0577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1217__A1 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__1218__A2 (.DIODE(_0585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1220__A2 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__1223__A2 (.DIODE(_0599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1225__A (.DIODE(_0451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1231__B1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__1234__C1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__1235__A (.DIODE(_0429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1235__B (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__1239__B (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__1243__A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__1246__B2 (.DIODE(_0630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1247__A1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__1247__B1 (.DIODE(_0428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1248__A0 (.DIODE(_0577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1249__A (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__1251__A0 (.DIODE(_0585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1252__A (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__1253__A (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__1256__A0 (.DIODE(_0599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1257__A (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__1258__A (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__1259__A0 (.DIODE(_0591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1260__A (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__1263__A0 (.DIODE(_0570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1264__A0 (.DIODE(_0564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1265__A (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__1266__A (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__1268__A0 (.DIODE(_0549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1269__A (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__1270__A (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__1271__A0 (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1272__A (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__1283__A (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__1284__A (.DIODE(_0632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1296__A (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__1326__A1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__1330__A1 (.DIODE(_0450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1331__B (.DIODE(\MOS6502.ALU.CO ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1332__A1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__1332__B2 (.DIODE(_0534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1339__B1 (.DIODE(_0723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1352__A1 (.DIODE(_0450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1362__A0 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__1362__A1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__1362__A2 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__1362__A3 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__1365__B (.DIODE(_0723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1367__A1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__1379__B (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__1380__B1 (.DIODE(_0630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1381__A1 (.DIODE(_0723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1382__A1 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__1424__B2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__1427__B2 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__1430__B2 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__1431__B2 (.DIODE(\MOS6502.ADD[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1434__B2 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__1436__A1 (.DIODE(_0428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1442__B2 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__1444__B2 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__1445__B2 (.DIODE(\MOS6502.ADD[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1447__B (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__1448__B (.DIODE(_0630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1451__A2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__1452__A2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__1457__D (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__1458__C (.DIODE(_0723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1461__A2 (.DIODE(_0723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1461__B2 (.DIODE(_0549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1462__A (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__1466__A2 (.DIODE(_0630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1467__C (.DIODE(_0835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1469__B (.DIODE(_0723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1470__A2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__1470__B1 (.DIODE(_0549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1471__A1 (.DIODE(\MOS6502.ADD[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1481__B1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__1483__A2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__1484__B1 (.DIODE(\MOS6502.ALU.CO ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1485__A1 (.DIODE(_0630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1495__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__1496__C (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__1497__A1 (.DIODE(_0450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1497__B1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__1498__A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__1500__A (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__1502__A (.DIODE(_0451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1502__B (.DIODE(_0599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1503__A2 (.DIODE(_0450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1510__B1 (.DIODE(_0451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1511__A1 (.DIODE(_0451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1511__A2 (.DIODE(_0591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1513__A (.DIODE(\MOS6502.ADD[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1514__A (.DIODE(\MOS6502.ADD[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1517__A (.DIODE(_0450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1517__B (.DIODE(_0585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1518__A1 (.DIODE(_0450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1521__A1 (.DIODE(\MOS6502.ADD[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1524__B1 (.DIODE(_0450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1525__A1 (.DIODE(_0451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1525__A2 (.DIODE(_0577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1527__A (.DIODE(_0451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1527__B (.DIODE(_0570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1528__A2 (.DIODE(_0450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1530__B (.DIODE(\MOS6502.ALU.CO ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1531__A1 (.DIODE(\MOS6502.ALU.CO ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1534__A (.DIODE(_0451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1535__A1 (.DIODE(_0451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1535__A2 (.DIODE(_0564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1541__A0 (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1541__S (.DIODE(_0451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1545__A (.DIODE(\MOS6502.ALU.CO ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1545__B (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__1546__A1 (.DIODE(\MOS6502.ADD[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1548__A (.DIODE(_0451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1549__A1 (.DIODE(_0451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1549__A2 (.DIODE(_0549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1559__B1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__1568__S (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__1572__A2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__1572__B1 (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1574__A2 (.DIODE(_0723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1574__B2 (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1583__A2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__1583__B1 (.DIODE(_0564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1585__A2 (.DIODE(_0723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1585__B2 (.DIODE(_0564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1594__A2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__1594__B1 (.DIODE(_0570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1596__A2 (.DIODE(_0723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1596__B2 (.DIODE(_0570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1609__A2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__1609__B1 (.DIODE(_0585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1610__A1 (.DIODE(\MOS6502.ADD[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1612__A2 (.DIODE(_0723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1612__B2 (.DIODE(_0585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1620__A2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__1620__B1 (.DIODE(_0577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1629__A2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__1629__B1 (.DIODE(_0591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1631__A2 (.DIODE(_0723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1631__B2 (.DIODE(_0591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1641__A2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__1641__B1 (.DIODE(_0599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1644__A2 (.DIODE(_0723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1644__B2 (.DIODE(_0599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1664__A2 (.DIODE(_0723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1664__B2 (.DIODE(_0577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1678__C1 (.DIODE(_0630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1695__C1 (.DIODE(_0630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1699__A0 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__1699__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__1700__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__1702__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__1703__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__1704__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__1705__A (.DIODE(_0429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1706__A1 (.DIODE(_0429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1706__A2 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__1708__A (.DIODE(_0429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1709__B2 (.DIODE(_0429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1710__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__1711__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__1712__A0 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__1712__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__1713__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__1717__A (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__1717__B (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__1718__A (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__1718__B (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__1720__B (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__1722__B1 (.DIODE(_0723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1728__B (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__1729__B1 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__1731__A2 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__1738__A1 (.DIODE(_0428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1740__A (.DIODE(\MOS6502.ADD[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1743__A1 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__1744__A1 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__1746__B1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__1750__A1 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__1752__B1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__1756__A1 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__1758__B1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__1762__A1 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__1764__B1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__1768__A1 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__1769__A1 (.DIODE(\MOS6502.ADD[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1769__C1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__1773__A1 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__1776__A (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__1777__A2 (.DIODE(_0534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1777__C1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__1778__A (.DIODE(_0599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1781__A1 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__1783__A2 (.DIODE(_0534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1783__C1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__1784__A (.DIODE(_0591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1787__A1 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__1789__A1 (.DIODE(\MOS6502.ADD[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1789__A2 (.DIODE(_0534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1789__C1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__1790__A (.DIODE(_0585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1793__A1 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__1795__A2 (.DIODE(_0534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1795__C1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__1796__A (.DIODE(_0577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1799__A1 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__1801__A2 (.DIODE(_0534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1801__C1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__1802__A (.DIODE(_0570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1805__A1 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__1807__A2 (.DIODE(_0534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1807__C1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__1808__A (.DIODE(_0564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1811__A1 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__1812__A2 (.DIODE(_0534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1812__C1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__1813__A1 (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1815__B1_N (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__1817__A1 (.DIODE(\MOS6502.ADD[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1817__A2 (.DIODE(_0534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1817__C1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__1818__A1 (.DIODE(_0549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1820__B2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__1824__B (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__1826__D (.DIODE(_0723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1830__A (.DIODE(_0429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1830__D (.DIODE(_0835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1832__S (.DIODE(_0274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1833__A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__1834__S (.DIODE(_0274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1835__A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__1836__S (.DIODE(_0274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1837__A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__1838__S (.DIODE(_0274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1839__A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__1840__S (.DIODE(_0274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1841__A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__1842__S (.DIODE(_0274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1843__A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__1844__S (.DIODE(_0274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1845__A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__1846__S (.DIODE(_0274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1847__A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__1848__S (.DIODE(_0274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1849__A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__1850__S (.DIODE(_0274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1851__A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__1852__S (.DIODE(_0274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1853__A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__1854__S (.DIODE(_0274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1855__A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__1856__S (.DIODE(_0274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1857__A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__1858__S (.DIODE(_0274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1859__A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__1860__S (.DIODE(_0274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1861__A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__1862__S (.DIODE(_0274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1863__A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__1864__B (.DIODE(_0599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1865__B (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__1866__B (.DIODE(_0585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1868__B (.DIODE(_0570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1869__A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__1870__A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__1870__B (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__1871__A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__1871__B (.DIODE(_0549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1873__A (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__1876__S (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__1877__A1 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__1878__A1 (.DIODE(_0599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1880__A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__1883__C1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__1886__A2 (.DIODE(_0591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1888__A (.DIODE(\MOS6502.ADD[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1888__D (.DIODE(\MOS6502.ADD[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1891__B1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__1893__A2 (.DIODE(_0630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1895__A (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__1896__A0 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__1896__A1 (.DIODE(_0549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1898__A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__1899__B2 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__1901__A1 (.DIODE(\MOS6502.ADD[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1902__A1 (.DIODE(_0585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1904__C1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__1905__A1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__1906__A1 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__1906__S (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__1909__A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__1912__A (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__1914__B2 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__1915__A2 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__1916__A0 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__1916__S (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__1918__A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__1919__A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__1919__B (.DIODE(_0835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1920__A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__1920__B (.DIODE(_0835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1921__A (.DIODE(_0429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1922__A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__1922__B (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__1924__B1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__1926__C1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__1927__A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__1927__A3 (.DIODE(_0835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1927__B1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__1930__C1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__1931__A1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__1931__A3 (.DIODE(_0835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1931__B1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__1934__C1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__1935__A1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__1935__A3 (.DIODE(_0835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1935__B1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__1937__A1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__1937__A3 (.DIODE(_0835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1939__A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__1939__A3 (.DIODE(_0835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1939__B1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__1941__A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__1941__B (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__1942__B1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__1969__B1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__1975__C1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__1983__C1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__1987__C1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__1994__A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__2003__A (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__2014__C1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__2023__C1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__2035__A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__2038__C1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__2045__A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__2047__A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__2051__A1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__2051__C1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__2053__B2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__2055__C_N (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__2056__A1 (.DIODE(_0428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2057__A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__2058__B1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__2067__B1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout52_A (.DIODE(_0632_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout63_A (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout73_A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout74_A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout75_A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout76_A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout77_A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout78_A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold147_A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold160_A (.DIODE(\MOS6502.ADD[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold167_A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold191_A (.DIODE(\MOS6502.ALU.CO ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold200_A (.DIODE(\MOS6502.ADD[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold214_A (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold217_A (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold223_A (.DIODE(_0564_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold225_A (.DIODE(_0591_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold229_A (.DIODE(_0577_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold232_A (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold234_A (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold236_A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_output15_A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_output16_A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_output27_A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_output35_A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_output36_A (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_output37_A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_output38_A (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_output39_A (.DIODE(net39));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_114 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_8 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_163 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_34 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_6 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__inv_2 _1025_ (.A(\MOS6502.NMI_edge ),
    .Y(_0428_));
 sky130_fd_sc_hd__inv_2 _1026_ (.A(net78),
    .Y(_0429_));
 sky130_fd_sc_hd__inv_2 _1027_ (.A(net269),
    .Y(_0430_));
 sky130_fd_sc_hd__inv_2 _1028_ (.A(net297),
    .Y(_0431_));
 sky130_fd_sc_hd__inv_2 _1029_ (.A(net235),
    .Y(_0432_));
 sky130_fd_sc_hd__inv_2 _1030_ (.A(\MOS6502.rotate ),
    .Y(_0433_));
 sky130_fd_sc_hd__inv_2 _1031_ (.A(net198),
    .Y(_0434_));
 sky130_fd_sc_hd__inv_2 _1032_ (.A(\MOS6502.load_only ),
    .Y(_0435_));
 sky130_fd_sc_hd__inv_2 _1033_ (.A(net233),
    .Y(_0436_));
 sky130_fd_sc_hd__inv_2 _1034_ (.A(net177),
    .Y(_0437_));
 sky130_fd_sc_hd__inv_2 _1035_ (.A(\MOS6502.ABL[1] ),
    .Y(_0438_));
 sky130_fd_sc_hd__inv_2 _1036_ (.A(net322),
    .Y(_0439_));
 sky130_fd_sc_hd__inv_2 _1037_ (.A(\MOS6502.state[4] ),
    .Y(_0440_));
 sky130_fd_sc_hd__inv_2 _1038_ (.A(net74),
    .Y(_0441_));
 sky130_fd_sc_hd__inv_2 _1039_ (.A(net11),
    .Y(_0442_));
 sky130_fd_sc_hd__and2b_1 _1040_ (.A_N(\MOS6502.state[4] ),
    .B(net322),
    .X(_0443_));
 sky130_fd_sc_hd__nand2b_1 _1041_ (.A_N(\MOS6502.state[4] ),
    .B(\MOS6502.state[5] ),
    .Y(_0444_));
 sky130_fd_sc_hd__or4b_2 _1042_ (.A(net68),
    .B(net69),
    .C(net71),
    .D_N(net70),
    .X(_0445_));
 sky130_fd_sc_hd__nor2_2 _1043_ (.A(net67),
    .B(_0445_),
    .Y(_0446_));
 sky130_fd_sc_hd__and2b_1 _1044_ (.A_N(\MOS6502.state[5] ),
    .B(\MOS6502.state[4] ),
    .X(_0447_));
 sky130_fd_sc_hd__nand2b_2 _1045_ (.A_N(\MOS6502.state[5] ),
    .B(\MOS6502.state[4] ),
    .Y(_0448_));
 sky130_fd_sc_hd__or4bb_4 _1046_ (.A(net69),
    .B(net71),
    .C_N(net70),
    .D_N(net68),
    .X(_0449_));
 sky130_fd_sc_hd__nor2_4 _1047_ (.A(net66),
    .B(_0449_),
    .Y(_0450_));
 sky130_fd_sc_hd__or2_4 _1048_ (.A(_0448_),
    .B(_0449_),
    .X(_0451_));
 sky130_fd_sc_hd__or4bb_4 _1049_ (.A(net68),
    .B(net70),
    .C_N(net71),
    .D_N(net69),
    .X(_0452_));
 sky130_fd_sc_hd__nor2_1 _1050_ (.A(net67),
    .B(_0452_),
    .Y(_0453_));
 sky130_fd_sc_hd__nor2_1 _1051_ (.A(net67),
    .B(_0449_),
    .Y(_0454_));
 sky130_fd_sc_hd__a21o_1 _1052_ (.A1(_0449_),
    .A2(_0452_),
    .B1(_0444_),
    .X(_0455_));
 sky130_fd_sc_hd__nand2_1 _1053_ (.A(_0451_),
    .B(_0455_),
    .Y(_0456_));
 sky130_fd_sc_hd__and3b_2 _1054_ (.A_N(_0446_),
    .B(_0451_),
    .C(_0455_),
    .X(_0457_));
 sky130_fd_sc_hd__or4b_2 _1055_ (.A(net69),
    .B(net70),
    .C(net71),
    .D_N(net68),
    .X(_0458_));
 sky130_fd_sc_hd__nor2_2 _1056_ (.A(\MOS6502.state[4] ),
    .B(_0458_),
    .Y(_0459_));
 sky130_fd_sc_hd__or3_4 _1057_ (.A(net282),
    .B(\MOS6502.state[4] ),
    .C(_0458_),
    .X(_0460_));
 sky130_fd_sc_hd__nand2_4 _1058_ (.A(_0457_),
    .B(_0460_),
    .Y(_0461_));
 sky130_fd_sc_hd__or2_1 _1059_ (.A(\MOS6502.state[5] ),
    .B(\MOS6502.state[4] ),
    .X(_0462_));
 sky130_fd_sc_hd__nand4b_4 _1060_ (.A_N(net71),
    .B(net70),
    .C(\MOS6502.state[2] ),
    .D(\MOS6502.state[3] ),
    .Y(_0463_));
 sky130_fd_sc_hd__nor2_1 _1061_ (.A(net65),
    .B(_0463_),
    .Y(_0464_));
 sky130_fd_sc_hd__nor2_1 _1062_ (.A(_0445_),
    .B(net65),
    .Y(_0465_));
 sky130_fd_sc_hd__a21oi_1 _1063_ (.A1(_0445_),
    .A2(_0463_),
    .B1(net65),
    .Y(_0466_));
 sky130_fd_sc_hd__or4bb_2 _1064_ (.A(\MOS6502.state[3] ),
    .B(net69),
    .C_N(net70),
    .D_N(net71),
    .X(_0467_));
 sky130_fd_sc_hd__nor2_2 _1065_ (.A(net66),
    .B(_0467_),
    .Y(_0468_));
 sky130_fd_sc_hd__nor3_1 _1066_ (.A(net68),
    .B(net69),
    .C(net70),
    .Y(_0469_));
 sky130_fd_sc_hd__or4_2 _1067_ (.A(net68),
    .B(\MOS6502.state[2] ),
    .C(\MOS6502.state[1] ),
    .D(\MOS6502.state[0] ),
    .X(_0470_));
 sky130_fd_sc_hd__nand2_1 _1068_ (.A(\MOS6502.state[5] ),
    .B(\MOS6502.state[4] ),
    .Y(_0471_));
 sky130_fd_sc_hd__nor2_1 _1069_ (.A(_0470_),
    .B(_0471_),
    .Y(_0472_));
 sky130_fd_sc_hd__or3_4 _1070_ (.A(_0466_),
    .B(_0468_),
    .C(_0472_),
    .X(_0473_));
 sky130_fd_sc_hd__nand2_1 _1071_ (.A(net68),
    .B(net69),
    .Y(_0474_));
 sky130_fd_sc_hd__or4bb_4 _1072_ (.A(net70),
    .B(net71),
    .C_N(net68),
    .D_N(net69),
    .X(_0475_));
 sky130_fd_sc_hd__nor2_2 _1073_ (.A(net65),
    .B(_0475_),
    .Y(_0476_));
 sky130_fd_sc_hd__or2_4 _1074_ (.A(net65),
    .B(_0475_),
    .X(_0477_));
 sky130_fd_sc_hd__nor4_1 _1075_ (.A(_0466_),
    .B(_0468_),
    .C(_0472_),
    .D(net55),
    .Y(_0478_));
 sky130_fd_sc_hd__nand4_2 _1076_ (.A(net68),
    .B(net69),
    .C(net70),
    .D(net71),
    .Y(_0479_));
 sky130_fd_sc_hd__nor2_1 _1077_ (.A(net66),
    .B(_0479_),
    .Y(_0480_));
 sky130_fd_sc_hd__nor2_1 _1078_ (.A(net67),
    .B(_0475_),
    .Y(_0481_));
 sky130_fd_sc_hd__o22a_1 _1079_ (.A1(net67),
    .A2(_0475_),
    .B1(_0479_),
    .B2(net66),
    .X(_0482_));
 sky130_fd_sc_hd__nor2_2 _1080_ (.A(net66),
    .B(_0475_),
    .Y(_0483_));
 sky130_fd_sc_hd__nand4b_4 _1081_ (.A_N(net69),
    .B(net70),
    .C(net71),
    .D(net68),
    .Y(_0484_));
 sky130_fd_sc_hd__nor2_2 _1082_ (.A(net65),
    .B(_0484_),
    .Y(_0485_));
 sky130_fd_sc_hd__o22ai_4 _1083_ (.A1(net66),
    .A2(_0475_),
    .B1(_0484_),
    .B2(net65),
    .Y(_0486_));
 sky130_fd_sc_hd__nor2_2 _1084_ (.A(_0448_),
    .B(_0463_),
    .Y(_0487_));
 sky130_fd_sc_hd__nor4b_4 _1085_ (.A(_0459_),
    .B(_0487_),
    .C(_0486_),
    .D_N(_0482_),
    .Y(_0488_));
 sky130_fd_sc_hd__and4_2 _1086_ (.A(\MOS6502.src_reg[1] ),
    .B(_0457_),
    .C(net51),
    .D(_0488_),
    .X(_0489_));
 sky130_fd_sc_hd__a211oi_4 _1087_ (.A1(\MOS6502.dst_reg[1] ),
    .A2(net55),
    .B1(_0489_),
    .C1(_0473_),
    .Y(_0490_));
 sky130_fd_sc_hd__a211o_4 _1088_ (.A1(\MOS6502.dst_reg[1] ),
    .A2(net55),
    .B1(_0489_),
    .C1(_0473_),
    .X(_0491_));
 sky130_fd_sc_hd__nand4b_4 _1089_ (.A_N(net145),
    .B(_0457_),
    .C(net51),
    .D(_0488_),
    .Y(_0492_));
 sky130_fd_sc_hd__and2_1 _1090_ (.A(\MOS6502.dst_reg[0] ),
    .B(net55),
    .X(_0493_));
 sky130_fd_sc_hd__a211o_4 _1091_ (.A1(\MOS6502.index_y ),
    .A2(_0473_),
    .B1(net51),
    .C1(_0493_),
    .X(_0494_));
 sky130_fd_sc_hd__and2_2 _1092_ (.A(_0492_),
    .B(_0494_),
    .X(_0495_));
 sky130_fd_sc_hd__nand2_8 _1093_ (.A(_0492_),
    .B(_0494_),
    .Y(_0496_));
 sky130_fd_sc_hd__mux2_1 _1094_ (.A0(net89),
    .A1(net129),
    .S(_0496_),
    .X(_0497_));
 sky130_fd_sc_hd__mux2_1 _1095_ (.A0(net101),
    .A1(net105),
    .S(_0496_),
    .X(_0498_));
 sky130_fd_sc_hd__mux2_1 _1096_ (.A0(_0497_),
    .A1(_0498_),
    .S(_0491_),
    .X(_0499_));
 sky130_fd_sc_hd__and4bb_1 _1097_ (.A_N(net69),
    .B_N(net70),
    .C(net71),
    .D(net68),
    .X(_0500_));
 sky130_fd_sc_hd__or4bb_4 _1098_ (.A(net69),
    .B(net70),
    .C_N(net71),
    .D_N(net68),
    .X(_0501_));
 sky130_fd_sc_hd__nor2_1 _1099_ (.A(net65),
    .B(_0501_),
    .Y(_0502_));
 sky130_fd_sc_hd__nor2_1 _1100_ (.A(net66),
    .B(_0484_),
    .Y(_0503_));
 sky130_fd_sc_hd__o22ai_4 _1101_ (.A1(net66),
    .A2(_0484_),
    .B1(_0501_),
    .B2(net65),
    .Y(_0504_));
 sky130_fd_sc_hd__nor2_1 _1102_ (.A(net67),
    .B(_0484_),
    .Y(_0505_));
 sky130_fd_sc_hd__and4b_1 _1103_ (.A_N(net68),
    .B(net69),
    .C(net70),
    .D(net71),
    .X(_0506_));
 sky130_fd_sc_hd__and2_4 _1104_ (.A(_0443_),
    .B(_0506_),
    .X(_0507_));
 sky130_fd_sc_hd__or3_1 _1105_ (.A(_0504_),
    .B(_0505_),
    .C(_0507_),
    .X(_0508_));
 sky130_fd_sc_hd__nor2_2 _1106_ (.A(_0449_),
    .B(net65),
    .Y(_0509_));
 sky130_fd_sc_hd__or4bb_2 _1107_ (.A(net68),
    .B(net71),
    .C_N(net70),
    .D_N(net69),
    .X(_0510_));
 sky130_fd_sc_hd__nor2_2 _1108_ (.A(net67),
    .B(_0510_),
    .Y(_0511_));
 sky130_fd_sc_hd__a21bo_1 _1109_ (.A1(\MOS6502.state[5] ),
    .A2(_0459_),
    .B1_N(_0482_),
    .X(_0512_));
 sky130_fd_sc_hd__or4_1 _1110_ (.A(_0508_),
    .B(_0509_),
    .C(_0511_),
    .D(_0512_),
    .X(_0513_));
 sky130_fd_sc_hd__nand2_1 _1111_ (.A(net323),
    .B(_0469_),
    .Y(_0514_));
 sky130_fd_sc_hd__nor2_1 _1112_ (.A(net66),
    .B(_0514_),
    .Y(_0515_));
 sky130_fd_sc_hd__nor2_1 _1113_ (.A(net67),
    .B(_0501_),
    .Y(_0516_));
 sky130_fd_sc_hd__or4b_2 _1114_ (.A(\MOS6502.state[3] ),
    .B(net70),
    .C(net71),
    .D_N(\MOS6502.state[2] ),
    .X(_0517_));
 sky130_fd_sc_hd__nor2_2 _1115_ (.A(net66),
    .B(_0517_),
    .Y(_0518_));
 sky130_fd_sc_hd__or3_1 _1116_ (.A(_0515_),
    .B(_0516_),
    .C(_0518_),
    .X(_0519_));
 sky130_fd_sc_hd__nor2_2 _1117_ (.A(net65),
    .B(_0467_),
    .Y(_0520_));
 sky130_fd_sc_hd__and3_1 _1118_ (.A(_0439_),
    .B(\MOS6502.state[4] ),
    .C(_0506_),
    .X(_0521_));
 sky130_fd_sc_hd__or2_1 _1119_ (.A(_0520_),
    .B(_0521_),
    .X(_0522_));
 sky130_fd_sc_hd__nor2_1 _1120_ (.A(net65),
    .B(_0514_),
    .Y(_0523_));
 sky130_fd_sc_hd__nor2_1 _1121_ (.A(net66),
    .B(_0501_),
    .Y(_0524_));
 sky130_fd_sc_hd__or2_1 _1122_ (.A(_0523_),
    .B(_0524_),
    .X(_0525_));
 sky130_fd_sc_hd__or3_4 _1123_ (.A(_0519_),
    .B(_0522_),
    .C(_0525_),
    .X(_0526_));
 sky130_fd_sc_hd__nor2_2 _1124_ (.A(net65),
    .B(_0510_),
    .Y(_0527_));
 sky130_fd_sc_hd__nor2_1 _1125_ (.A(net66),
    .B(_0470_),
    .Y(_0528_));
 sky130_fd_sc_hd__nor2_1 _1126_ (.A(_0471_),
    .B(_0514_),
    .Y(_0529_));
 sky130_fd_sc_hd__nor2_2 _1127_ (.A(_0462_),
    .B(_0479_),
    .Y(_0530_));
 sky130_fd_sc_hd__or2_1 _1128_ (.A(_0468_),
    .B(_0530_),
    .X(_0531_));
 sky130_fd_sc_hd__or4_1 _1129_ (.A(net53),
    .B(_0528_),
    .C(_0529_),
    .D(_0531_),
    .X(_0532_));
 sky130_fd_sc_hd__or3_4 _1130_ (.A(_0513_),
    .B(_0526_),
    .C(_0532_),
    .X(_0533_));
 sky130_fd_sc_hd__and3_4 _1131_ (.A(_0439_),
    .B(_0440_),
    .C(_0506_),
    .X(_0534_));
 sky130_fd_sc_hd__inv_2 _1132_ (.A(_0534_),
    .Y(_0535_));
 sky130_fd_sc_hd__nor2_1 _1133_ (.A(net66),
    .B(_0452_),
    .Y(_0536_));
 sky130_fd_sc_hd__nor2_1 _1134_ (.A(net65),
    .B(_0517_),
    .Y(_0537_));
 sky130_fd_sc_hd__or3_4 _1135_ (.A(_0534_),
    .B(_0536_),
    .C(_0537_),
    .X(_0538_));
 sky130_fd_sc_hd__nor2_1 _1136_ (.A(net67),
    .B(_0467_),
    .Y(_0539_));
 sky130_fd_sc_hd__nor2_2 _1137_ (.A(net67),
    .B(_0517_),
    .Y(_0540_));
 sky130_fd_sc_hd__or2_1 _1138_ (.A(net67),
    .B(_0517_),
    .X(_0541_));
 sky130_fd_sc_hd__or2_2 _1139_ (.A(_0539_),
    .B(_0540_),
    .X(_0542_));
 sky130_fd_sc_hd__nor2_8 _1140_ (.A(net67),
    .B(_0463_),
    .Y(_0543_));
 sky130_fd_sc_hd__or2_2 _1141_ (.A(net67),
    .B(_0463_),
    .X(_0544_));
 sky130_fd_sc_hd__or3_4 _1142_ (.A(_0538_),
    .B(_0542_),
    .C(_0543_),
    .X(_0545_));
 sky130_fd_sc_hd__nor2_1 _1143_ (.A(_0445_),
    .B(net66),
    .Y(_0546_));
 sky130_fd_sc_hd__nor2_1 _1144_ (.A(net67),
    .B(_0479_),
    .Y(_0547_));
 sky130_fd_sc_hd__or2_4 _1145_ (.A(_0546_),
    .B(_0547_),
    .X(_0548_));
 sky130_fd_sc_hd__mux2_4 _1146_ (.A0(net310),
    .A1(net192),
    .S(net78),
    .X(_0549_));
 sky130_fd_sc_hd__a22o_1 _1147_ (.A1(net279),
    .A2(_0545_),
    .B1(_0548_),
    .B2(_0549_),
    .X(_0550_));
 sky130_fd_sc_hd__a221o_1 _1148_ (.A1(_0461_),
    .A2(_0499_),
    .B1(_0533_),
    .B2(net244),
    .C1(_0550_),
    .X(_0551_));
 sky130_fd_sc_hd__nor4_4 _1149_ (.A(_0461_),
    .B(_0533_),
    .C(_0545_),
    .D(_0548_),
    .Y(_0552_));
 sky130_fd_sc_hd__mux2_2 _1150_ (.A0(_0551_),
    .A1(net209),
    .S(net47),
    .X(net17));
 sky130_fd_sc_hd__mux2_1 _1151_ (.A0(\MOS6502.AXYS[1][6] ),
    .A1(\MOS6502.AXYS[0][6] ),
    .S(_0496_),
    .X(_0553_));
 sky130_fd_sc_hd__nand2_1 _1152_ (.A(\MOS6502.AXYS[3][6] ),
    .B(_0495_),
    .Y(_0554_));
 sky130_fd_sc_hd__a21oi_1 _1153_ (.A1(\MOS6502.AXYS[2][6] ),
    .A2(_0496_),
    .B1(_0490_),
    .Y(_0555_));
 sky130_fd_sc_hd__a2bb2o_1 _1154_ (.A1_N(_0491_),
    .A2_N(_0553_),
    .B1(_0554_),
    .B2(_0555_),
    .X(_0556_));
 sky130_fd_sc_hd__inv_2 _1155_ (.A(_0556_),
    .Y(_0557_));
 sky130_fd_sc_hd__mux2_4 _1156_ (.A0(net300),
    .A1(\MOS6502.DI[6] ),
    .S(net78),
    .X(_0558_));
 sky130_fd_sc_hd__a22o_1 _1157_ (.A1(net262),
    .A2(_0545_),
    .B1(_0548_),
    .B2(_0558_),
    .X(_0559_));
 sky130_fd_sc_hd__a221o_1 _1158_ (.A1(\MOS6502.ADD[6] ),
    .A2(_0533_),
    .B1(_0557_),
    .B2(_0461_),
    .C1(_0559_),
    .X(_0560_));
 sky130_fd_sc_hd__a21o_1 _1159_ (.A1(net211),
    .A2(_0552_),
    .B1(_0560_),
    .X(net46));
 sky130_fd_sc_hd__mux2_1 _1160_ (.A0(\MOS6502.AXYS[1][5] ),
    .A1(\MOS6502.AXYS[0][5] ),
    .S(_0496_),
    .X(_0561_));
 sky130_fd_sc_hd__mux2_1 _1161_ (.A0(\MOS6502.AXYS[3][5] ),
    .A1(\MOS6502.AXYS[2][5] ),
    .S(_0496_),
    .X(_0562_));
 sky130_fd_sc_hd__mux2_1 _1162_ (.A0(_0561_),
    .A1(_0562_),
    .S(_0491_),
    .X(_0563_));
 sky130_fd_sc_hd__mux2_4 _1163_ (.A0(net306),
    .A1(\MOS6502.DI[5] ),
    .S(net78),
    .X(_0564_));
 sky130_fd_sc_hd__a22o_1 _1164_ (.A1(net267),
    .A2(_0545_),
    .B1(_0548_),
    .B2(_0564_),
    .X(_0565_));
 sky130_fd_sc_hd__a221o_1 _1165_ (.A1(net264),
    .A2(_0533_),
    .B1(_0563_),
    .B2(_0461_),
    .C1(_0565_),
    .X(_0566_));
 sky130_fd_sc_hd__a21o_1 _1166_ (.A1(net225),
    .A2(_0552_),
    .B1(_0566_),
    .X(net45));
 sky130_fd_sc_hd__mux2_1 _1167_ (.A0(\MOS6502.AXYS[1][4] ),
    .A1(\MOS6502.AXYS[0][4] ),
    .S(_0496_),
    .X(_0567_));
 sky130_fd_sc_hd__mux2_1 _1168_ (.A0(\MOS6502.AXYS[3][4] ),
    .A1(\MOS6502.AXYS[2][4] ),
    .S(_0496_),
    .X(_0568_));
 sky130_fd_sc_hd__mux2_1 _1169_ (.A0(_0567_),
    .A1(_0568_),
    .S(_0491_),
    .X(_0569_));
 sky130_fd_sc_hd__mux2_4 _1170_ (.A0(net296),
    .A1(net180),
    .S(net78),
    .X(_0570_));
 sky130_fd_sc_hd__a22o_1 _1171_ (.A1(net266),
    .A2(_0545_),
    .B1(_0548_),
    .B2(_0570_),
    .X(_0571_));
 sky130_fd_sc_hd__a221o_1 _1172_ (.A1(net255),
    .A2(_0533_),
    .B1(_0569_),
    .B2(_0461_),
    .C1(_0571_),
    .X(_0572_));
 sky130_fd_sc_hd__a21o_1 _1173_ (.A1(net221),
    .A2(_0552_),
    .B1(_0572_),
    .X(net44));
 sky130_fd_sc_hd__and3_1 _1174_ (.A(\MOS6502.AXYS[1][3] ),
    .B(_0492_),
    .C(_0494_),
    .X(_0573_));
 sky130_fd_sc_hd__mux2_1 _1175_ (.A0(\MOS6502.AXYS[3][3] ),
    .A1(\MOS6502.AXYS[2][3] ),
    .S(_0496_),
    .X(_0574_));
 sky130_fd_sc_hd__a211o_1 _1176_ (.A1(\MOS6502.AXYS[0][3] ),
    .A2(_0496_),
    .B1(_0573_),
    .C1(_0491_),
    .X(_0575_));
 sky130_fd_sc_hd__o21a_1 _1177_ (.A1(_0490_),
    .A2(_0574_),
    .B1(_0575_),
    .X(_0576_));
 sky130_fd_sc_hd__mux2_4 _1178_ (.A0(net312),
    .A1(\MOS6502.DI[3] ),
    .S(net78),
    .X(_0577_));
 sky130_fd_sc_hd__a22o_1 _1179_ (.A1(net270),
    .A2(_0545_),
    .B1(_0548_),
    .B2(_0577_),
    .X(_0578_));
 sky130_fd_sc_hd__a221o_1 _1180_ (.A1(\MOS6502.ADD[3] ),
    .A2(_0533_),
    .B1(_0576_),
    .B2(_0461_),
    .C1(_0578_),
    .X(_0579_));
 sky130_fd_sc_hd__a21o_1 _1181_ (.A1(net213),
    .A2(_0552_),
    .B1(_0579_),
    .X(net43));
 sky130_fd_sc_hd__a21o_1 _1182_ (.A1(_0492_),
    .A2(_0494_),
    .B1(\MOS6502.AXYS[0][2] ),
    .X(_0580_));
 sky130_fd_sc_hd__a21o_1 _1183_ (.A1(_0492_),
    .A2(_0494_),
    .B1(\MOS6502.AXYS[2][2] ),
    .X(_0581_));
 sky130_fd_sc_hd__o211ai_2 _1184_ (.A1(\MOS6502.AXYS[1][2] ),
    .A2(_0496_),
    .B1(_0580_),
    .C1(_0490_),
    .Y(_0582_));
 sky130_fd_sc_hd__o211ai_1 _1185_ (.A1(\MOS6502.AXYS[3][2] ),
    .A2(_0496_),
    .B1(_0581_),
    .C1(_0491_),
    .Y(_0583_));
 sky130_fd_sc_hd__nand2_1 _1186_ (.A(_0582_),
    .B(_0583_),
    .Y(_0584_));
 sky130_fd_sc_hd__mux2_4 _1187_ (.A0(net305),
    .A1(net186),
    .S(net78),
    .X(_0585_));
 sky130_fd_sc_hd__a22o_1 _1188_ (.A1(net274),
    .A2(_0545_),
    .B1(_0548_),
    .B2(_0585_),
    .X(_0586_));
 sky130_fd_sc_hd__a221o_1 _1189_ (.A1(\MOS6502.ADD[2] ),
    .A2(_0533_),
    .B1(_0584_),
    .B2(_0461_),
    .C1(_0586_),
    .X(_0587_));
 sky130_fd_sc_hd__a21o_1 _1190_ (.A1(net217),
    .A2(_0552_),
    .B1(_0587_),
    .X(net42));
 sky130_fd_sc_hd__mux2_1 _1191_ (.A0(\MOS6502.AXYS[0][1] ),
    .A1(\MOS6502.AXYS[1][1] ),
    .S(_0495_),
    .X(_0588_));
 sky130_fd_sc_hd__mux2_1 _1192_ (.A0(\MOS6502.AXYS[2][1] ),
    .A1(\MOS6502.AXYS[3][1] ),
    .S(_0495_),
    .X(_0589_));
 sky130_fd_sc_hd__mux2_1 _1193_ (.A0(_0588_),
    .A1(_0589_),
    .S(_0491_),
    .X(_0590_));
 sky130_fd_sc_hd__mux2_4 _1194_ (.A0(net308),
    .A1(\MOS6502.DI[1] ),
    .S(net78),
    .X(_0591_));
 sky130_fd_sc_hd__a22o_1 _1195_ (.A1(\MOS6502.ABL[1] ),
    .A2(_0545_),
    .B1(_0548_),
    .B2(_0591_),
    .X(_0592_));
 sky130_fd_sc_hd__a221o_1 _1196_ (.A1(net261),
    .A2(_0533_),
    .B1(_0590_),
    .B2(_0461_),
    .C1(_0592_),
    .X(_0593_));
 sky130_fd_sc_hd__a21o_1 _1197_ (.A1(net219),
    .A2(_0552_),
    .B1(_0593_),
    .X(net41));
 sky130_fd_sc_hd__a21o_1 _1198_ (.A1(_0492_),
    .A2(_0494_),
    .B1(\MOS6502.AXYS[0][0] ),
    .X(_0594_));
 sky130_fd_sc_hd__a21o_1 _1199_ (.A1(_0492_),
    .A2(_0494_),
    .B1(\MOS6502.AXYS[2][0] ),
    .X(_0595_));
 sky130_fd_sc_hd__o211ai_2 _1200_ (.A1(\MOS6502.AXYS[1][0] ),
    .A2(_0496_),
    .B1(_0594_),
    .C1(_0490_),
    .Y(_0596_));
 sky130_fd_sc_hd__o211ai_2 _1201_ (.A1(\MOS6502.AXYS[3][0] ),
    .A2(_0496_),
    .B1(_0595_),
    .C1(_0491_),
    .Y(_0597_));
 sky130_fd_sc_hd__nand2_1 _1202_ (.A(_0596_),
    .B(_0597_),
    .Y(_0598_));
 sky130_fd_sc_hd__mux2_4 _1203_ (.A0(net304),
    .A1(net178),
    .S(net78),
    .X(_0599_));
 sky130_fd_sc_hd__a22o_1 _1204_ (.A1(net260),
    .A2(_0545_),
    .B1(_0548_),
    .B2(_0599_),
    .X(_0600_));
 sky130_fd_sc_hd__a221o_1 _1205_ (.A1(net259),
    .A2(_0533_),
    .B1(_0598_),
    .B2(_0461_),
    .C1(_0600_),
    .X(_0601_));
 sky130_fd_sc_hd__a21o_2 _1206_ (.A1(net223),
    .A2(_0552_),
    .B1(_0601_),
    .X(net40));
 sky130_fd_sc_hd__or3_4 _1207_ (.A(_0527_),
    .B(_0542_),
    .C(_0543_),
    .X(_0602_));
 sky130_fd_sc_hd__a22o_1 _1208_ (.A1(_0526_),
    .A2(_0549_),
    .B1(_0602_),
    .B2(net288),
    .X(_0603_));
 sky130_fd_sc_hd__a221o_1 _1209_ (.A1(net244),
    .A2(_0538_),
    .B1(net47),
    .B2(net200),
    .C1(_0603_),
    .X(net25));
 sky130_fd_sc_hd__a22o_1 _1210_ (.A1(_0526_),
    .A2(_0558_),
    .B1(_0602_),
    .B2(net290),
    .X(_0604_));
 sky130_fd_sc_hd__a221o_1 _1211_ (.A1(net277),
    .A2(_0538_),
    .B1(net47),
    .B2(net202),
    .C1(_0604_),
    .X(net24));
 sky130_fd_sc_hd__a22o_1 _1212_ (.A1(_0526_),
    .A2(_0564_),
    .B1(_0602_),
    .B2(net295),
    .X(_0605_));
 sky130_fd_sc_hd__a221o_1 _1213_ (.A1(net264),
    .A2(_0538_),
    .B1(net47),
    .B2(net196),
    .C1(_0605_),
    .X(net23));
 sky130_fd_sc_hd__a22o_1 _1214_ (.A1(_0526_),
    .A2(_0570_),
    .B1(_0602_),
    .B2(net291),
    .X(_0606_));
 sky130_fd_sc_hd__a221o_1 _1215_ (.A1(net255),
    .A2(_0538_),
    .B1(net47),
    .B2(net190),
    .C1(_0606_),
    .X(net22));
 sky130_fd_sc_hd__a22o_1 _1216_ (.A1(_0526_),
    .A2(_0577_),
    .B1(_0602_),
    .B2(net293),
    .X(_0607_));
 sky130_fd_sc_hd__a221o_2 _1217_ (.A1(net278),
    .A2(_0538_),
    .B1(net47),
    .B2(net194),
    .C1(_0607_),
    .X(net21));
 sky130_fd_sc_hd__a22o_1 _1218_ (.A1(_0526_),
    .A2(_0585_),
    .B1(_0602_),
    .B2(net302),
    .X(_0608_));
 sky130_fd_sc_hd__a221o_2 _1219_ (.A1(net284),
    .A2(_0538_),
    .B1(net47),
    .B2(net188),
    .C1(_0608_),
    .X(net20));
 sky130_fd_sc_hd__a22o_1 _1220_ (.A1(_0526_),
    .A2(net309),
    .B1(_0602_),
    .B2(net311),
    .X(_0609_));
 sky130_fd_sc_hd__a221o_2 _1221_ (.A1(net261),
    .A2(_0538_),
    .B1(net47),
    .B2(net182),
    .C1(_0609_),
    .X(net19));
 sky130_fd_sc_hd__a221o_1 _1222_ (.A1(\MOS6502.ADD[0] ),
    .A2(_0538_),
    .B1(_0602_),
    .B2(\MOS6502.ABH[0] ),
    .C1(_0513_),
    .X(_0610_));
 sky130_fd_sc_hd__a211o_1 _1223_ (.A1(_0526_),
    .A2(_0599_),
    .B1(_0610_),
    .C1(_0461_),
    .X(_0611_));
 sky130_fd_sc_hd__a21o_1 _1224_ (.A1(net184),
    .A2(_0552_),
    .B1(_0611_),
    .X(net18));
 sky130_fd_sc_hd__nand2_4 _1225_ (.A(_0451_),
    .B(_0460_),
    .Y(_0612_));
 sky130_fd_sc_hd__or2_1 _1226_ (.A(_0446_),
    .B(_0509_),
    .X(_0613_));
 sky130_fd_sc_hd__or3_4 _1227_ (.A(_0504_),
    .B(_0612_),
    .C(_0613_),
    .X(_0614_));
 sky130_fd_sc_hd__nor2_2 _1228_ (.A(_0543_),
    .B(_0614_),
    .Y(_0615_));
 sky130_fd_sc_hd__or4_2 _1229_ (.A(_0523_),
    .B(_0529_),
    .C(_0537_),
    .D(_0547_),
    .X(_0616_));
 sky130_fd_sc_hd__o31a_1 _1230_ (.A1(_0515_),
    .A2(_0536_),
    .A3(_0616_),
    .B1(\MOS6502.store ),
    .X(_0617_));
 sky130_fd_sc_hd__o31ai_4 _1231_ (.A1(_0543_),
    .A2(_0614_),
    .A3(_0617_),
    .B1(net77),
    .Y(net15));
 sky130_fd_sc_hd__and3b_2 _1232_ (.A_N(net2),
    .B(net1),
    .C(clknet_4_10_0_wb_clk_i),
    .X(_0618_));
 sky130_fd_sc_hd__nor2_2 _1233_ (.A(clknet_4_10_0_wb_clk_i),
    .B(net1),
    .Y(_0619_));
 sky130_fd_sc_hd__a211oi_2 _1234_ (.A1(net2),
    .A2(_0619_),
    .B1(_0618_),
    .C1(net15),
    .Y(net35));
 sky130_fd_sc_hd__nor2_1 _1235_ (.A(_0429_),
    .B(net72),
    .Y(_0620_));
 sky130_fd_sc_hd__and4b_2 _1236_ (.A_N(net70),
    .B(net71),
    .C(net68),
    .D(net69),
    .X(_0621_));
 sky130_fd_sc_hd__o21a_1 _1237_ (.A1(_0443_),
    .A2(_0447_),
    .B1(_0621_),
    .X(_0622_));
 sky130_fd_sc_hd__or4_1 _1238_ (.A(_0515_),
    .B(_0536_),
    .C(_0543_),
    .D(_0622_),
    .X(_0623_));
 sky130_fd_sc_hd__or2_1 _1239_ (.A(net215),
    .B(net275),
    .X(_0624_));
 sky130_fd_sc_hd__a21oi_1 _1240_ (.A1(_0436_),
    .A2(_0520_),
    .B1(_0518_),
    .Y(_0625_));
 sky130_fd_sc_hd__nor2_1 _1241_ (.A(_0624_),
    .B(_0625_),
    .Y(_0626_));
 sky130_fd_sc_hd__a211o_1 _1242_ (.A1(_0436_),
    .A2(_0616_),
    .B1(_0623_),
    .C1(_0626_),
    .X(_0627_));
 sky130_fd_sc_hd__nor2_1 _1243_ (.A(net78),
    .B(_0441_),
    .Y(_0628_));
 sky130_fd_sc_hd__a32o_1 _1244_ (.A1(_0443_),
    .A2(_0621_),
    .A3(net56),
    .B1(_0481_),
    .B2(net61),
    .X(_0629_));
 sky130_fd_sc_hd__and3_4 _1245_ (.A(_0439_),
    .B(_0440_),
    .C(_0621_),
    .X(_0630_));
 sky130_fd_sc_hd__a22o_1 _1246_ (.A1(net63),
    .A2(_0627_),
    .B1(net58),
    .B2(_0630_),
    .X(_0631_));
 sky130_fd_sc_hd__o21a_1 _1247_ (.A1(net37),
    .A2(_0442_),
    .B1(_0428_),
    .X(_0632_));
 sky130_fd_sc_hd__mux2_1 _1248_ (.A0(_0577_),
    .A1(net85),
    .S(net236),
    .X(_0633_));
 sky130_fd_sc_hd__and2_2 _1249_ (.A(net52),
    .B(_0633_),
    .X(_0634_));
 sky130_fd_sc_hd__inv_2 _1250_ (.A(_0634_),
    .Y(_0635_));
 sky130_fd_sc_hd__mux2_1 _1251_ (.A0(_0585_),
    .A1(\MOS6502.IRHOLD[2] ),
    .S(\MOS6502.IRHOLD_valid ),
    .X(_0636_));
 sky130_fd_sc_hd__and2_2 _1252_ (.A(net52),
    .B(_0636_),
    .X(_0637_));
 sky130_fd_sc_hd__nand2_2 _1253_ (.A(net52),
    .B(_0636_),
    .Y(_0638_));
 sky130_fd_sc_hd__nand2_1 _1254_ (.A(_0634_),
    .B(_0638_),
    .Y(_0639_));
 sky130_fd_sc_hd__inv_2 _1255_ (.A(_0639_),
    .Y(_0640_));
 sky130_fd_sc_hd__mux2_1 _1256_ (.A0(_0599_),
    .A1(\MOS6502.IRHOLD[0] ),
    .S(\MOS6502.IRHOLD_valid ),
    .X(_0641_));
 sky130_fd_sc_hd__and2_1 _1257_ (.A(net52),
    .B(_0641_),
    .X(_0642_));
 sky130_fd_sc_hd__nand2_2 _1258_ (.A(net52),
    .B(_0641_),
    .Y(_0643_));
 sky130_fd_sc_hd__mux2_1 _1259_ (.A0(_0591_),
    .A1(net87),
    .S(\MOS6502.IRHOLD_valid ),
    .X(_0644_));
 sky130_fd_sc_hd__and2_2 _1260_ (.A(net52),
    .B(_0644_),
    .X(_0645_));
 sky130_fd_sc_hd__or2_2 _1261_ (.A(_0642_),
    .B(_0645_),
    .X(_0646_));
 sky130_fd_sc_hd__or2_2 _1262_ (.A(_0639_),
    .B(_0646_),
    .X(_0647_));
 sky130_fd_sc_hd__mux2_2 _1263_ (.A0(_0570_),
    .A1(net325),
    .S(net236),
    .X(_0648_));
 sky130_fd_sc_hd__mux2_1 _1264_ (.A0(_0564_),
    .A1(net111),
    .S(\MOS6502.IRHOLD_valid ),
    .X(_0649_));
 sky130_fd_sc_hd__and2_4 _1265_ (.A(net52),
    .B(_0649_),
    .X(_0650_));
 sky130_fd_sc_hd__nand2_4 _1266_ (.A(net52),
    .B(_0649_),
    .Y(_0651_));
 sky130_fd_sc_hd__or2_1 _1267_ (.A(_0648_),
    .B(_0651_),
    .X(_0652_));
 sky130_fd_sc_hd__mux2_4 _1268_ (.A0(_0549_),
    .A1(net91),
    .S(\MOS6502.IRHOLD_valid ),
    .X(_0653_));
 sky130_fd_sc_hd__and2_2 _1269_ (.A(net52),
    .B(_0653_),
    .X(_0654_));
 sky130_fd_sc_hd__nand2_4 _1270_ (.A(net52),
    .B(_0653_),
    .Y(_0655_));
 sky130_fd_sc_hd__mux2_1 _1271_ (.A0(_0558_),
    .A1(net137),
    .S(\MOS6502.IRHOLD_valid ),
    .X(_0656_));
 sky130_fd_sc_hd__and2_4 _1272_ (.A(net52),
    .B(_0656_),
    .X(_0657_));
 sky130_fd_sc_hd__and2b_1 _1273_ (.A_N(_0653_),
    .B(_0657_),
    .X(_0658_));
 sky130_fd_sc_hd__nand2b_1 _1274_ (.A_N(_0653_),
    .B(_0657_),
    .Y(_0659_));
 sky130_fd_sc_hd__or2_1 _1275_ (.A(_0652_),
    .B(_0659_),
    .X(_0660_));
 sky130_fd_sc_hd__inv_2 _1276_ (.A(_0660_),
    .Y(_0661_));
 sky130_fd_sc_hd__nand2_1 _1277_ (.A(_0634_),
    .B(_0637_),
    .Y(_0662_));
 sky130_fd_sc_hd__or2_1 _1278_ (.A(_0646_),
    .B(_0662_),
    .X(_0663_));
 sky130_fd_sc_hd__nor2_1 _1279_ (.A(_0660_),
    .B(_0663_),
    .Y(_0664_));
 sky130_fd_sc_hd__o32a_1 _1280_ (.A1(_0647_),
    .A2(_0652_),
    .A3(_0654_),
    .B1(_0660_),
    .B2(_0663_),
    .X(_0665_));
 sky130_fd_sc_hd__nor2_1 _1281_ (.A(_0639_),
    .B(_0642_),
    .Y(_0666_));
 sky130_fd_sc_hd__o31a_1 _1282_ (.A1(_0645_),
    .A2(_0648_),
    .A3(_0654_),
    .B1(_0666_),
    .X(_0667_));
 sky130_fd_sc_hd__and2_2 _1283_ (.A(net52),
    .B(_0648_),
    .X(_0668_));
 sky130_fd_sc_hd__nand2_2 _1284_ (.A(_0632_),
    .B(_0648_),
    .Y(_0669_));
 sky130_fd_sc_hd__nand2_1 _1285_ (.A(_0651_),
    .B(_0669_),
    .Y(_0670_));
 sky130_fd_sc_hd__nor2_1 _1286_ (.A(_0659_),
    .B(_0670_),
    .Y(_0671_));
 sky130_fd_sc_hd__or3_1 _1287_ (.A(_0659_),
    .B(_0663_),
    .C(_0670_),
    .X(_0672_));
 sky130_fd_sc_hd__inv_2 _1288_ (.A(_0672_),
    .Y(_0673_));
 sky130_fd_sc_hd__nor2_2 _1289_ (.A(_0643_),
    .B(_0645_),
    .Y(_0674_));
 sky130_fd_sc_hd__or2_2 _1290_ (.A(_0643_),
    .B(_0645_),
    .X(_0675_));
 sky130_fd_sc_hd__a211o_1 _1291_ (.A1(_0638_),
    .A2(_0675_),
    .B1(_0669_),
    .C1(_0635_),
    .X(_0676_));
 sky130_fd_sc_hd__or4_1 _1292_ (.A(_0637_),
    .B(_0646_),
    .C(_0654_),
    .D(_0670_),
    .X(_0677_));
 sky130_fd_sc_hd__nor2_1 _1293_ (.A(_0634_),
    .B(_0637_),
    .Y(_0678_));
 sky130_fd_sc_hd__or2_1 _1294_ (.A(_0634_),
    .B(_0637_),
    .X(_0679_));
 sky130_fd_sc_hd__and2_1 _1295_ (.A(_0476_),
    .B(net63),
    .X(_0680_));
 sky130_fd_sc_hd__nand2_2 _1296_ (.A(net55),
    .B(net63),
    .Y(_0681_));
 sky130_fd_sc_hd__or2_1 _1297_ (.A(_0634_),
    .B(_0638_),
    .X(_0682_));
 sky130_fd_sc_hd__o211a_1 _1298_ (.A1(_0675_),
    .A2(_0679_),
    .B1(_0680_),
    .C1(_0682_),
    .X(_0683_));
 sky130_fd_sc_hd__and3_1 _1299_ (.A(_0676_),
    .B(_0677_),
    .C(_0683_),
    .X(_0684_));
 sky130_fd_sc_hd__and4b_1 _1300_ (.A_N(_0667_),
    .B(_0672_),
    .C(_0684_),
    .D(_0665_),
    .X(_0685_));
 sky130_fd_sc_hd__or2_1 _1301_ (.A(_0654_),
    .B(_0657_),
    .X(_0686_));
 sky130_fd_sc_hd__or2_2 _1302_ (.A(_0652_),
    .B(_0686_),
    .X(_0687_));
 sky130_fd_sc_hd__inv_2 _1303_ (.A(_0687_),
    .Y(_0688_));
 sky130_fd_sc_hd__o21a_1 _1304_ (.A1(_0648_),
    .A2(_0655_),
    .B1(_0687_),
    .X(_0689_));
 sky130_fd_sc_hd__and2_2 _1305_ (.A(_0643_),
    .B(_0645_),
    .X(_0690_));
 sky130_fd_sc_hd__nand2_1 _1306_ (.A(_0643_),
    .B(_0645_),
    .Y(_0691_));
 sky130_fd_sc_hd__nor2_1 _1307_ (.A(_0674_),
    .B(_0690_),
    .Y(_0692_));
 sky130_fd_sc_hd__o32a_1 _1308_ (.A1(_0662_),
    .A2(_0668_),
    .A3(_0692_),
    .B1(_0689_),
    .B2(_0663_),
    .X(_0693_));
 sky130_fd_sc_hd__or2_1 _1309_ (.A(_0646_),
    .B(_0679_),
    .X(_0694_));
 sky130_fd_sc_hd__a31o_1 _1310_ (.A1(_0660_),
    .A2(_0669_),
    .A3(_0687_),
    .B1(_0694_),
    .X(_0695_));
 sky130_fd_sc_hd__and3_1 _1311_ (.A(_0685_),
    .B(_0693_),
    .C(_0695_),
    .X(_0696_));
 sky130_fd_sc_hd__or3_1 _1312_ (.A(_0629_),
    .B(_0631_),
    .C(_0696_),
    .X(_0697_));
 sky130_fd_sc_hd__nor2_1 _1313_ (.A(_0681_),
    .B(_0694_),
    .Y(_0698_));
 sky130_fd_sc_hd__a22o_1 _1314_ (.A1(_0453_),
    .A2(net58),
    .B1(_0671_),
    .B2(_0698_),
    .X(_0699_));
 sky130_fd_sc_hd__a32o_1 _1315_ (.A1(_0518_),
    .A2(net63),
    .A3(_0624_),
    .B1(net58),
    .B2(_0536_),
    .X(_0700_));
 sky130_fd_sc_hd__or3_1 _1316_ (.A(_0697_),
    .B(_0699_),
    .C(_0700_),
    .X(_0701_));
 sky130_fd_sc_hd__nor2_1 _1317_ (.A(_0681_),
    .B(_0682_),
    .Y(_0702_));
 sky130_fd_sc_hd__a22o_1 _1318_ (.A1(_0547_),
    .A2(net58),
    .B1(_0669_),
    .B2(_0702_),
    .X(_0703_));
 sky130_fd_sc_hd__a221o_1 _1319_ (.A1(_0464_),
    .A2(net63),
    .B1(net59),
    .B2(_0530_),
    .C1(_0703_),
    .X(_0704_));
 sky130_fd_sc_hd__nor2_1 _1320_ (.A(net66),
    .B(_0510_),
    .Y(_0705_));
 sky130_fd_sc_hd__a22o_1 _1321_ (.A1(_0521_),
    .A2(net57),
    .B1(_0705_),
    .B2(net61),
    .X(_0706_));
 sky130_fd_sc_hd__a22o_1 _1322_ (.A1(_0511_),
    .A2(net62),
    .B1(net56),
    .B2(_0507_),
    .X(_0707_));
 sky130_fd_sc_hd__or3_1 _1323_ (.A(_0704_),
    .B(_0706_),
    .C(_0707_),
    .X(_0708_));
 sky130_fd_sc_hd__a32o_1 _1324_ (.A1(net233),
    .A2(_0616_),
    .A3(net63),
    .B1(net58),
    .B2(_0539_),
    .X(_0709_));
 sky130_fd_sc_hd__a22o_1 _1325_ (.A1(_0454_),
    .A2(net62),
    .B1(net57),
    .B2(_0505_),
    .X(_0710_));
 sky130_fd_sc_hd__a221o_1 _1326_ (.A1(net54),
    .A2(net62),
    .B1(net57),
    .B2(_0485_),
    .C1(_0710_),
    .X(_0711_));
 sky130_fd_sc_hd__a22o_1 _1327_ (.A1(_0487_),
    .A2(net61),
    .B1(net56),
    .B2(_0480_),
    .X(_0712_));
 sky130_fd_sc_hd__a22o_1 _1328_ (.A1(_0546_),
    .A2(net61),
    .B1(net56),
    .B2(_0468_),
    .X(_0713_));
 sky130_fd_sc_hd__a221o_1 _1329_ (.A1(_0465_),
    .A2(net61),
    .B1(net56),
    .B2(_0520_),
    .C1(_0713_),
    .X(_0714_));
 sky130_fd_sc_hd__a22o_1 _1330_ (.A1(_0450_),
    .A2(net61),
    .B1(net56),
    .B2(_0503_),
    .X(_0715_));
 sky130_fd_sc_hd__xor2_2 _1331_ (.A(\MOS6502.backwards ),
    .B(\MOS6502.ALU.CO ),
    .X(_0716_));
 sky130_fd_sc_hd__a32o_1 _1332_ (.A1(net53),
    .A2(net62),
    .A3(_0716_),
    .B1(net56),
    .B2(_0534_),
    .X(_0717_));
 sky130_fd_sc_hd__or4_1 _1333_ (.A(_0712_),
    .B(_0714_),
    .C(_0715_),
    .D(_0717_),
    .X(_0718_));
 sky130_fd_sc_hd__or4_1 _1334_ (.A(_0708_),
    .B(_0709_),
    .C(_0711_),
    .D(_0718_),
    .X(_0719_));
 sky130_fd_sc_hd__nor2_1 _1335_ (.A(net67),
    .B(_0514_),
    .Y(_0720_));
 sky130_fd_sc_hd__or3_1 _1336_ (.A(_0635_),
    .B(_0677_),
    .C(_0681_),
    .X(_0721_));
 sky130_fd_sc_hd__a21bo_1 _1337_ (.A1(net58),
    .A2(_0720_),
    .B1_N(_0721_),
    .X(_0722_));
 sky130_fd_sc_hd__nor2_8 _1338_ (.A(_0452_),
    .B(net65),
    .Y(_0723_));
 sky130_fd_sc_hd__a22o_1 _1339_ (.A1(_0668_),
    .A2(_0698_),
    .B1(_0723_),
    .B2(net58),
    .X(_0724_));
 sky130_fd_sc_hd__and2_1 _1340_ (.A(_0516_),
    .B(net56),
    .X(_0725_));
 sky130_fd_sc_hd__a221o_1 _1341_ (.A1(_0459_),
    .A2(net61),
    .B1(net56),
    .B2(_0502_),
    .C1(_0725_),
    .X(_0726_));
 sky130_fd_sc_hd__a22o_1 _1342_ (.A1(_0472_),
    .A2(net62),
    .B1(net56),
    .B2(_0529_),
    .X(_0727_));
 sky130_fd_sc_hd__a221o_1 _1343_ (.A1(_0528_),
    .A2(net62),
    .B1(net57),
    .B2(_0515_),
    .C1(_0727_),
    .X(_0728_));
 sky130_fd_sc_hd__nor2_1 _1344_ (.A(net65),
    .B(_0470_),
    .Y(_0729_));
 sky130_fd_sc_hd__nor2_1 _1345_ (.A(net66),
    .B(_0458_),
    .Y(_0730_));
 sky130_fd_sc_hd__or2_1 _1346_ (.A(_0729_),
    .B(_0730_),
    .X(_0731_));
 sky130_fd_sc_hd__a32o_1 _1347_ (.A1(_0447_),
    .A2(_0621_),
    .A3(net56),
    .B1(_0483_),
    .B2(net61),
    .X(_0732_));
 sky130_fd_sc_hd__a221o_1 _1348_ (.A1(_0525_),
    .A2(net57),
    .B1(_0731_),
    .B2(net61),
    .C1(_0732_),
    .X(_0733_));
 sky130_fd_sc_hd__or4_1 _1349_ (.A(_0724_),
    .B(_0726_),
    .C(_0728_),
    .D(_0733_),
    .X(_0734_));
 sky130_fd_sc_hd__or4_1 _1350_ (.A(_0701_),
    .B(_0719_),
    .C(_0722_),
    .D(_0734_),
    .X(_0001_));
 sky130_fd_sc_hd__a22o_1 _1351_ (.A1(_0454_),
    .A2(net58),
    .B1(_0661_),
    .B2(_0698_),
    .X(_0735_));
 sky130_fd_sc_hd__a22o_1 _1352_ (.A1(_0450_),
    .A2(net58),
    .B1(_0688_),
    .B2(_0698_),
    .X(_0736_));
 sky130_fd_sc_hd__or2_1 _1353_ (.A(_0735_),
    .B(_0736_),
    .X(_0737_));
 sky130_fd_sc_hd__a22o_1 _1354_ (.A1(_0539_),
    .A2(net63),
    .B1(net58),
    .B2(_0543_),
    .X(_0738_));
 sky130_fd_sc_hd__or4_1 _1355_ (.A(_0647_),
    .B(_0652_),
    .C(_0654_),
    .D(_0681_),
    .X(_0739_));
 sky130_fd_sc_hd__a21bo_1 _1356_ (.A1(_0487_),
    .A2(net58),
    .B1_N(_0739_),
    .X(_0740_));
 sky130_fd_sc_hd__or2_1 _1357_ (.A(_0738_),
    .B(_0740_),
    .X(_0741_));
 sky130_fd_sc_hd__o21a_1 _1358_ (.A1(_0485_),
    .A2(_0524_),
    .B1(net61),
    .X(_0742_));
 sky130_fd_sc_hd__a221o_1 _1359_ (.A1(_0673_),
    .A2(_0680_),
    .B1(_0705_),
    .B2(net57),
    .C1(_0742_),
    .X(_0743_));
 sky130_fd_sc_hd__and3_1 _1360_ (.A(_0674_),
    .B(_0678_),
    .C(_0680_),
    .X(_0744_));
 sky130_fd_sc_hd__a22o_1 _1361_ (.A1(_0464_),
    .A2(net58),
    .B1(_0669_),
    .B2(_0744_),
    .X(_0745_));
 sky130_fd_sc_hd__mux4_1 _1362_ (.A0(net39),
    .A1(net16),
    .A2(net38),
    .A3(net27),
    .S0(\MOS6502.cond_code[2] ),
    .S1(\MOS6502.cond_code[1] ),
    .X(_0746_));
 sky130_fd_sc_hd__xnor2_1 _1363_ (.A(net171),
    .B(_0746_),
    .Y(_0747_));
 sky130_fd_sc_hd__inv_2 _1364_ (.A(_0747_),
    .Y(_0748_));
 sky130_fd_sc_hd__and3_1 _1365_ (.A(net62),
    .B(_0723_),
    .C(_0747_),
    .X(_0749_));
 sky130_fd_sc_hd__a22o_1 _1366_ (.A1(_0453_),
    .A2(net62),
    .B1(net57),
    .B2(_0511_),
    .X(_0750_));
 sky130_fd_sc_hd__a211o_1 _1367_ (.A1(net53),
    .A2(net57),
    .B1(_0749_),
    .C1(_0750_),
    .X(_0751_));
 sky130_fd_sc_hd__or3_1 _1368_ (.A(_0741_),
    .B(_0743_),
    .C(_0745_),
    .X(_0752_));
 sky130_fd_sc_hd__or3_1 _1369_ (.A(_0737_),
    .B(_0751_),
    .C(_0752_),
    .X(_0753_));
 sky130_fd_sc_hd__a22o_1 _1370_ (.A1(_0502_),
    .A2(net63),
    .B1(net58),
    .B2(_0509_),
    .X(_0754_));
 sky130_fd_sc_hd__a22o_1 _1371_ (.A1(_0446_),
    .A2(net58),
    .B1(_0720_),
    .B2(net63),
    .X(_0755_));
 sky130_fd_sc_hd__a22o_1 _1372_ (.A1(_0546_),
    .A2(net58),
    .B1(_0668_),
    .B2(_0744_),
    .X(_0756_));
 sky130_fd_sc_hd__a2111oi_1 _1373_ (.A1(_0465_),
    .A2(net58),
    .B1(_0754_),
    .C1(_0755_),
    .D1(_0756_),
    .Y(_0757_));
 sky130_fd_sc_hd__o21ai_1 _1374_ (.A1(_0676_),
    .A2(_0681_),
    .B1(_0757_),
    .Y(_0758_));
 sky130_fd_sc_hd__or3_1 _1375_ (.A(_0719_),
    .B(_0753_),
    .C(_0758_),
    .X(_0002_));
 sky130_fd_sc_hd__a22o_1 _1376_ (.A1(_0540_),
    .A2(net59),
    .B1(_0667_),
    .B2(_0680_),
    .X(_0759_));
 sky130_fd_sc_hd__nor2_1 _1377_ (.A(net67),
    .B(_0470_),
    .Y(_0760_));
 sky130_fd_sc_hd__or4_1 _1378_ (.A(_0446_),
    .B(_0516_),
    .C(_0540_),
    .D(_0760_),
    .X(_0761_));
 sky130_fd_sc_hd__and2b_1 _1379_ (.A_N(_0716_),
    .B(net53),
    .X(_0762_));
 sky130_fd_sc_hd__a211o_1 _1380_ (.A1(_0439_),
    .A2(_0506_),
    .B1(_0630_),
    .C1(_0762_),
    .X(_0763_));
 sky130_fd_sc_hd__a211o_1 _1381_ (.A1(_0723_),
    .A2(_0748_),
    .B1(_0761_),
    .C1(_0763_),
    .X(_0764_));
 sky130_fd_sc_hd__a22o_1 _1382_ (.A1(net55),
    .A2(net56),
    .B1(_0764_),
    .B2(net61),
    .X(_0765_));
 sky130_fd_sc_hd__a22o_1 _1383_ (.A1(_0503_),
    .A2(net61),
    .B1(net56),
    .B2(_0483_),
    .X(_0766_));
 sky130_fd_sc_hd__a221o_1 _1384_ (.A1(_0468_),
    .A2(net62),
    .B1(net57),
    .B2(_0518_),
    .C1(_0766_),
    .X(_0767_));
 sky130_fd_sc_hd__a22o_1 _1385_ (.A1(_0505_),
    .A2(net62),
    .B1(net57),
    .B2(_0481_),
    .X(_0768_));
 sky130_fd_sc_hd__o211a_1 _1386_ (.A1(net233),
    .A2(_0624_),
    .B1(net63),
    .C1(_0520_),
    .X(_0769_));
 sky130_fd_sc_hd__a211o_1 _1387_ (.A1(_0537_),
    .A2(net56),
    .B1(_0768_),
    .C1(_0769_),
    .X(_0770_));
 sky130_fd_sc_hd__or4_1 _1388_ (.A(_0759_),
    .B(_0765_),
    .C(_0767_),
    .D(_0770_),
    .X(_0771_));
 sky130_fd_sc_hd__or2_1 _1389_ (.A(_0712_),
    .B(_0732_),
    .X(_0772_));
 sky130_fd_sc_hd__or4_1 _1390_ (.A(_0717_),
    .B(_0724_),
    .C(_0751_),
    .D(_0772_),
    .X(_0773_));
 sky130_fd_sc_hd__or4_1 _1391_ (.A(_0708_),
    .B(_0752_),
    .C(_0771_),
    .D(_0773_),
    .X(_0774_));
 sky130_fd_sc_hd__or2_1 _1392_ (.A(_0701_),
    .B(_0774_),
    .X(_0003_));
 sky130_fd_sc_hd__nor2_1 _1393_ (.A(_0681_),
    .B(_0693_),
    .Y(_0775_));
 sky130_fd_sc_hd__a22o_1 _1394_ (.A1(_0664_),
    .A2(_0680_),
    .B1(_0730_),
    .B2(net57),
    .X(_0776_));
 sky130_fd_sc_hd__a32o_1 _1395_ (.A1(net282),
    .A2(_0459_),
    .A3(net56),
    .B1(net61),
    .B2(_0507_),
    .X(_0777_));
 sky130_fd_sc_hd__or2_1 _1396_ (.A(_0776_),
    .B(_0777_),
    .X(_0778_));
 sky130_fd_sc_hd__a22o_1 _1397_ (.A1(_0472_),
    .A2(net59),
    .B1(_0668_),
    .B2(_0702_),
    .X(_0779_));
 sky130_fd_sc_hd__a221o_1 _1398_ (.A1(_0530_),
    .A2(net62),
    .B1(net57),
    .B2(_0528_),
    .C1(_0779_),
    .X(_0780_));
 sky130_fd_sc_hd__a22o_1 _1399_ (.A1(_0480_),
    .A2(net61),
    .B1(net56),
    .B2(_0760_),
    .X(_0781_));
 sky130_fd_sc_hd__a211o_1 _1400_ (.A1(net57),
    .A2(_0729_),
    .B1(_0780_),
    .C1(_0781_),
    .X(_0782_));
 sky130_fd_sc_hd__or4_1 _1401_ (.A(_0771_),
    .B(_0775_),
    .C(_0778_),
    .D(_0782_),
    .X(_0783_));
 sky130_fd_sc_hd__or4_1 _1402_ (.A(_0001_),
    .B(_0753_),
    .C(_0758_),
    .D(_0783_),
    .X(_0784_));
 sky130_fd_sc_hd__a221o_1 _1403_ (.A1(_0524_),
    .A2(net57),
    .B1(_0730_),
    .B2(net61),
    .C1(_0715_),
    .X(_0785_));
 sky130_fd_sc_hd__or2_1 _1404_ (.A(_0772_),
    .B(_0785_),
    .X(_0786_));
 sky130_fd_sc_hd__or4_1 _1405_ (.A(_0711_),
    .B(_0754_),
    .C(_0766_),
    .D(_0768_),
    .X(_0787_));
 sky130_fd_sc_hd__or3_1 _1406_ (.A(_0726_),
    .B(_0786_),
    .C(_0787_),
    .X(_0788_));
 sky130_fd_sc_hd__or4_1 _1407_ (.A(_0704_),
    .B(_0745_),
    .C(_0765_),
    .D(_0788_),
    .X(_0789_));
 sky130_fd_sc_hd__or4_1 _1408_ (.A(_0737_),
    .B(_0741_),
    .C(_0778_),
    .D(_0789_),
    .X(_0790_));
 sky130_fd_sc_hd__or3b_1 _1409_ (.A(_0697_),
    .B(_0790_),
    .C_N(_0784_),
    .X(_0004_));
 sky130_fd_sc_hd__or4_1 _1410_ (.A(_0700_),
    .B(_0706_),
    .C(_0713_),
    .D(_0767_),
    .X(_0791_));
 sky130_fd_sc_hd__or4_1 _1411_ (.A(_0728_),
    .B(_0756_),
    .C(_0786_),
    .D(_0791_),
    .X(_0792_));
 sky130_fd_sc_hd__or3_1 _1412_ (.A(_0736_),
    .B(_0740_),
    .C(_0792_),
    .X(_0793_));
 sky130_fd_sc_hd__or4_1 _1413_ (.A(_0743_),
    .B(_0776_),
    .C(_0780_),
    .D(_0793_),
    .X(_0005_));
 sky130_fd_sc_hd__or4_1 _1414_ (.A(_0629_),
    .B(_0707_),
    .C(_0750_),
    .D(_0768_),
    .X(_0794_));
 sky130_fd_sc_hd__a311o_1 _1415_ (.A1(net282),
    .A2(_0459_),
    .A3(net61),
    .B1(_0725_),
    .C1(_0777_),
    .X(_0795_));
 sky130_fd_sc_hd__or4_1 _1416_ (.A(_0710_),
    .B(_0727_),
    .C(_0794_),
    .D(_0795_),
    .X(_0796_));
 sky130_fd_sc_hd__or4_1 _1417_ (.A(_0709_),
    .B(_0738_),
    .C(_0755_),
    .D(_0781_),
    .X(_0797_));
 sky130_fd_sc_hd__or4_1 _1418_ (.A(_0703_),
    .B(_0779_),
    .C(_0796_),
    .D(_0797_),
    .X(_0798_));
 sky130_fd_sc_hd__or2_1 _1419_ (.A(_0722_),
    .B(_0798_),
    .X(_0799_));
 sky130_fd_sc_hd__or4_1 _1420_ (.A(_0699_),
    .B(_0735_),
    .C(_0759_),
    .D(_0799_),
    .X(_0006_));
 sky130_fd_sc_hd__or2_1 _1421_ (.A(_0446_),
    .B(_0543_),
    .X(_0800_));
 sky130_fd_sc_hd__a21boi_4 _1422_ (.A1(\MOS6502.php ),
    .A2(_0544_),
    .B1_N(_0800_),
    .Y(_0801_));
 sky130_fd_sc_hd__a21o_2 _1423_ (.A1(\MOS6502.php ),
    .A2(_0446_),
    .B1(_0509_),
    .X(_0802_));
 sky130_fd_sc_hd__a22o_1 _1424_ (.A1(\MOS6502.PC[8] ),
    .A2(_0612_),
    .B1(_0802_),
    .B2(net16),
    .X(_0803_));
 sky130_fd_sc_hd__a22o_1 _1425_ (.A1(\MOS6502.PC[0] ),
    .A2(_0504_),
    .B1(_0801_),
    .B2(\MOS6502.ADD[0] ),
    .X(_0804_));
 sky130_fd_sc_hd__a211o_1 _1426_ (.A1(_0598_),
    .A2(_0615_),
    .B1(_0803_),
    .C1(_0804_),
    .X(net26));
 sky130_fd_sc_hd__a22o_1 _1427_ (.A1(\MOS6502.PC[1] ),
    .A2(_0504_),
    .B1(_0802_),
    .B2(net27),
    .X(_0805_));
 sky130_fd_sc_hd__a22o_1 _1428_ (.A1(\MOS6502.PC[9] ),
    .A2(_0612_),
    .B1(_0801_),
    .B2(\MOS6502.ADD[1] ),
    .X(_0806_));
 sky130_fd_sc_hd__a211o_1 _1429_ (.A1(_0590_),
    .A2(_0615_),
    .B1(_0805_),
    .C1(_0806_),
    .X(net28));
 sky130_fd_sc_hd__a22o_1 _1430_ (.A1(\MOS6502.PC[2] ),
    .A2(_0504_),
    .B1(_0802_),
    .B2(net37),
    .X(_0807_));
 sky130_fd_sc_hd__a22o_1 _1431_ (.A1(\MOS6502.PC[10] ),
    .A2(_0612_),
    .B1(_0801_),
    .B2(\MOS6502.ADD[2] ),
    .X(_0808_));
 sky130_fd_sc_hd__a211o_1 _1432_ (.A1(_0584_),
    .A2(_0615_),
    .B1(_0807_),
    .C1(_0808_),
    .X(net29));
 sky130_fd_sc_hd__and2_1 _1433_ (.A(\MOS6502.PC[3] ),
    .B(_0504_),
    .X(_0809_));
 sky130_fd_sc_hd__a221o_1 _1434_ (.A1(\MOS6502.PC[11] ),
    .A2(_0612_),
    .B1(_0802_),
    .B2(net36),
    .C1(_0809_),
    .X(_0810_));
 sky130_fd_sc_hd__a221o_1 _1435_ (.A1(_0576_),
    .A2(_0615_),
    .B1(_0801_),
    .B2(\MOS6502.ADD[3] ),
    .C1(_0810_),
    .X(net30));
 sky130_fd_sc_hd__a32o_1 _1436_ (.A1(_0428_),
    .A2(_0442_),
    .A3(_0509_),
    .B1(_0446_),
    .B2(\MOS6502.php ),
    .X(_0811_));
 sky130_fd_sc_hd__a221o_1 _1437_ (.A1(\MOS6502.PC[4] ),
    .A2(_0504_),
    .B1(_0800_),
    .B2(\MOS6502.ADD[4] ),
    .C1(_0811_),
    .X(_0812_));
 sky130_fd_sc_hd__a221o_1 _1438_ (.A1(\MOS6502.PC[12] ),
    .A2(_0612_),
    .B1(_0615_),
    .B2(_0569_),
    .C1(_0812_),
    .X(net31));
 sky130_fd_sc_hd__a221o_1 _1439_ (.A1(\MOS6502.PC[5] ),
    .A2(_0504_),
    .B1(_0800_),
    .B2(\MOS6502.ADD[5] ),
    .C1(_0802_),
    .X(_0813_));
 sky130_fd_sc_hd__a221o_1 _1440_ (.A1(\MOS6502.PC[13] ),
    .A2(_0612_),
    .B1(_0615_),
    .B2(_0563_),
    .C1(_0813_),
    .X(net32));
 sky130_fd_sc_hd__and2_1 _1441_ (.A(\MOS6502.PC[6] ),
    .B(_0504_),
    .X(_0814_));
 sky130_fd_sc_hd__a221o_1 _1442_ (.A1(\MOS6502.PC[14] ),
    .A2(_0612_),
    .B1(_0802_),
    .B2(net38),
    .C1(_0814_),
    .X(_0815_));
 sky130_fd_sc_hd__a221o_1 _1443_ (.A1(_0557_),
    .A2(_0615_),
    .B1(_0801_),
    .B2(\MOS6502.ADD[6] ),
    .C1(_0815_),
    .X(net33));
 sky130_fd_sc_hd__a22o_1 _1444_ (.A1(\MOS6502.PC[7] ),
    .A2(_0504_),
    .B1(_0802_),
    .B2(net39),
    .X(_0816_));
 sky130_fd_sc_hd__a221o_1 _1445_ (.A1(\MOS6502.PC[15] ),
    .A2(_0612_),
    .B1(_0801_),
    .B2(\MOS6502.ADD[7] ),
    .C1(_0816_),
    .X(_0817_));
 sky130_fd_sc_hd__a21o_1 _1446_ (.A1(_0499_),
    .A2(_0615_),
    .B1(_0817_),
    .X(net34));
 sky130_fd_sc_hd__and2_1 _1447_ (.A(net198),
    .B(net36),
    .X(_0000_));
 sky130_fd_sc_hd__or2_4 _1448_ (.A(_0542_),
    .B(_0630_),
    .X(_0818_));
 sky130_fd_sc_hd__and2_1 _1449_ (.A(net206),
    .B(_0818_),
    .X(_0819_));
 sky130_fd_sc_hd__nand2_2 _1450_ (.A(net206),
    .B(_0818_),
    .Y(_0820_));
 sky130_fd_sc_hd__a221oi_4 _1451_ (.A1(\MOS6502.backwards ),
    .A2(net53),
    .B1(_0818_),
    .B2(\MOS6502.op[2] ),
    .C1(_0614_),
    .Y(_0821_));
 sky130_fd_sc_hd__a221o_2 _1452_ (.A1(\MOS6502.backwards ),
    .A2(net53),
    .B1(_0818_),
    .B2(\MOS6502.op[2] ),
    .C1(_0614_),
    .X(_0822_));
 sky130_fd_sc_hd__and2_2 _1453_ (.A(net253),
    .B(_0818_),
    .X(_0823_));
 sky130_fd_sc_hd__nand2_2 _1454_ (.A(net253),
    .B(_0818_),
    .Y(_0824_));
 sky130_fd_sc_hd__or4_4 _1455_ (.A(_0508_),
    .B(_0509_),
    .C(_0511_),
    .D(_0530_),
    .X(_0825_));
 sky130_fd_sc_hd__nand2_1 _1456_ (.A(net283),
    .B(_0477_),
    .Y(_0826_));
 sky130_fd_sc_hd__or4_2 _1457_ (.A(_0487_),
    .B(_0511_),
    .C(_0523_),
    .D(net53),
    .X(_0827_));
 sky130_fd_sc_hd__or4_1 _1458_ (.A(_0483_),
    .B(_0613_),
    .C(_0723_),
    .D(_0826_),
    .X(_0828_));
 sky130_fd_sc_hd__or4_1 _1459_ (.A(_0456_),
    .B(_0502_),
    .C(_0542_),
    .D(_0720_),
    .X(_0829_));
 sky130_fd_sc_hd__nor4_4 _1460_ (.A(_0825_),
    .B(_0827_),
    .C(_0828_),
    .D(_0829_),
    .Y(_0830_));
 sky130_fd_sc_hd__a22o_1 _1461_ (.A1(\MOS6502.PC[7] ),
    .A2(_0723_),
    .B1(_0830_),
    .B2(_0549_),
    .X(_0831_));
 sky130_fd_sc_hd__nor3_2 _1462_ (.A(net55),
    .B(_0523_),
    .C(_0818_),
    .Y(_0832_));
 sky130_fd_sc_hd__a21oi_4 _1463_ (.A1(\MOS6502.op[0] ),
    .A2(_0818_),
    .B1(_0832_),
    .Y(_0833_));
 sky130_fd_sc_hd__a21o_2 _1464_ (.A1(\MOS6502.op[0] ),
    .A2(_0818_),
    .B1(_0832_),
    .X(_0834_));
 sky130_fd_sc_hd__or2_4 _1465_ (.A(_0487_),
    .B(_0720_),
    .X(_0835_));
 sky130_fd_sc_hd__a211o_1 _1466_ (.A1(_0435_),
    .A2(_0630_),
    .B1(_0540_),
    .C1(_0483_),
    .X(_0836_));
 sky130_fd_sc_hd__or4_4 _1467_ (.A(_0461_),
    .B(_0473_),
    .C(_0835_),
    .D(_0836_),
    .X(_0837_));
 sky130_fd_sc_hd__inv_2 _1468_ (.A(_0837_),
    .Y(_0838_));
 sky130_fd_sc_hd__or2_4 _1469_ (.A(_0539_),
    .B(_0723_),
    .X(_0839_));
 sky130_fd_sc_hd__a22o_1 _1470_ (.A1(\MOS6502.ABH[7] ),
    .A2(net53),
    .B1(_0549_),
    .B2(_0839_),
    .X(_0840_));
 sky130_fd_sc_hd__a221o_2 _1471_ (.A1(\MOS6502.ADD[7] ),
    .A2(_0825_),
    .B1(_0837_),
    .B2(_0499_),
    .C1(_0840_),
    .X(_0841_));
 sky130_fd_sc_hd__nand2_1 _1472_ (.A(\MOS6502.op[1] ),
    .B(_0818_),
    .Y(_0842_));
 sky130_fd_sc_hd__and2b_2 _1473_ (.A_N(_0832_),
    .B(_0842_),
    .X(_0843_));
 sky130_fd_sc_hd__nand2b_1 _1474_ (.A_N(_0832_),
    .B(_0842_),
    .Y(_0844_));
 sky130_fd_sc_hd__nor2_2 _1475_ (.A(_0833_),
    .B(_0843_),
    .Y(_0845_));
 sky130_fd_sc_hd__and3_1 _1476_ (.A(_0831_),
    .B(_0841_),
    .C(_0843_),
    .X(_0846_));
 sky130_fd_sc_hd__a21oi_1 _1477_ (.A1(_0831_),
    .A2(_0841_),
    .B1(_0834_),
    .Y(_0847_));
 sky130_fd_sc_hd__a21o_1 _1478_ (.A1(_0831_),
    .A2(_0833_),
    .B1(_0841_),
    .X(_0848_));
 sky130_fd_sc_hd__o311a_1 _1479_ (.A1(_0845_),
    .A2(_0846_),
    .A3(_0847_),
    .B1(_0848_),
    .C1(_0824_),
    .X(_0849_));
 sky130_fd_sc_hd__o21ai_1 _1480_ (.A1(\MOS6502.shift ),
    .A2(\MOS6502.load_only ),
    .B1(_0433_),
    .Y(_0850_));
 sky130_fd_sc_hd__a22o_1 _1481_ (.A1(_0433_),
    .A2(\MOS6502.compare ),
    .B1(net16),
    .B2(_0850_),
    .X(_0851_));
 sky130_fd_sc_hd__nor2_1 _1482_ (.A(\MOS6502.rotate ),
    .B(\MOS6502.shift ),
    .Y(_0852_));
 sky130_fd_sc_hd__a22o_1 _1483_ (.A1(\MOS6502.rotate ),
    .A2(net16),
    .B1(_0852_),
    .B2(\MOS6502.inc ),
    .X(_0853_));
 sky130_fd_sc_hd__o31a_1 _1484_ (.A1(_0518_),
    .A2(_0520_),
    .A3(_0527_),
    .B1(\MOS6502.ALU.CO ),
    .X(_0854_));
 sky130_fd_sc_hd__a22o_1 _1485_ (.A1(_0630_),
    .A2(_0851_),
    .B1(_0853_),
    .B2(_0542_),
    .X(_0855_));
 sky130_fd_sc_hd__or4_1 _1486_ (.A(_0487_),
    .B(_0505_),
    .C(_0507_),
    .D(_0511_),
    .X(_0856_));
 sky130_fd_sc_hd__or4b_1 _1487_ (.A(_0530_),
    .B(_0546_),
    .C(_0856_),
    .D_N(_0455_),
    .X(_0857_));
 sky130_fd_sc_hd__or3_1 _1488_ (.A(_0854_),
    .B(_0855_),
    .C(_0857_),
    .X(_0858_));
 sky130_fd_sc_hd__a21oi_1 _1489_ (.A1(_0823_),
    .A2(_0858_),
    .B1(_0849_),
    .Y(_0859_));
 sky130_fd_sc_hd__o21a_1 _1490_ (.A1(_0822_),
    .A2(_0859_),
    .B1(_0819_),
    .X(_0860_));
 sky130_fd_sc_hd__nand2_2 _1491_ (.A(_0820_),
    .B(_0821_),
    .Y(_0861_));
 sky130_fd_sc_hd__nor2_1 _1492_ (.A(_0831_),
    .B(_0861_),
    .Y(_0862_));
 sky130_fd_sc_hd__a211o_1 _1493_ (.A1(_0822_),
    .A2(_0831_),
    .B1(_0860_),
    .C1(_0862_),
    .X(_0863_));
 sky130_fd_sc_hd__inv_2 _1494_ (.A(_0863_),
    .Y(_0864_));
 sky130_fd_sc_hd__mux2_1 _1495_ (.A0(net169),
    .A1(_0864_),
    .S(net79),
    .X(_0007_));
 sky130_fd_sc_hd__and3b_1 _1496_ (.A_N(\MOS6502.plp ),
    .B(\MOS6502.load_reg ),
    .C(net55),
    .X(_0865_));
 sky130_fd_sc_hd__o41a_2 _1497_ (.A1(_0450_),
    .A2(_0486_),
    .A3(_0512_),
    .A4(_0865_),
    .B1(net78),
    .X(_0866_));
 sky130_fd_sc_hd__and2_2 _1498_ (.A(net14),
    .B(_0866_),
    .X(_0867_));
 sky130_fd_sc_hd__and3_1 _1499_ (.A(_0491_),
    .B(_0496_),
    .C(_0867_),
    .X(_0868_));
 sky130_fd_sc_hd__or2_4 _1500_ (.A(net72),
    .B(_0868_),
    .X(_0869_));
 sky130_fd_sc_hd__inv_2 _1501_ (.A(_0869_),
    .Y(_0870_));
 sky130_fd_sc_hd__or2_1 _1502_ (.A(_0451_),
    .B(_0599_),
    .X(_0871_));
 sky130_fd_sc_hd__o211a_1 _1503_ (.A1(\MOS6502.ADD[0] ),
    .A2(_0450_),
    .B1(_0867_),
    .C1(_0871_),
    .X(_0872_));
 sky130_fd_sc_hd__mux2_1 _1504_ (.A0(net149),
    .A1(_0872_),
    .S(_0869_),
    .X(_0008_));
 sky130_fd_sc_hd__and3_1 _1505_ (.A(\MOS6502.adc_bcd ),
    .B(\MOS6502.adj_bcd ),
    .C(\MOS6502.ALU.HC ),
    .X(_0873_));
 sky130_fd_sc_hd__nand2b_1 _1506_ (.A_N(\MOS6502.adc_bcd ),
    .B(\MOS6502.adj_bcd ),
    .Y(_0874_));
 sky130_fd_sc_hd__nor2_1 _1507_ (.A(\MOS6502.ALU.HC ),
    .B(_0874_),
    .Y(_0875_));
 sky130_fd_sc_hd__o21a_1 _1508_ (.A1(_0873_),
    .A2(_0875_),
    .B1(\MOS6502.ADD[1] ),
    .X(_0876_));
 sky130_fd_sc_hd__nor3_1 _1509_ (.A(\MOS6502.ADD[1] ),
    .B(_0873_),
    .C(_0875_),
    .Y(_0877_));
 sky130_fd_sc_hd__o21ai_1 _1510_ (.A1(_0876_),
    .A2(_0877_),
    .B1(_0451_),
    .Y(_0878_));
 sky130_fd_sc_hd__o211a_1 _1511_ (.A1(_0451_),
    .A2(_0591_),
    .B1(_0867_),
    .C1(_0878_),
    .X(_0879_));
 sky130_fd_sc_hd__mux2_1 _1512_ (.A0(net93),
    .A1(_0879_),
    .S(_0869_),
    .X(_0009_));
 sky130_fd_sc_hd__nand2_1 _1513_ (.A(\MOS6502.ADD[2] ),
    .B(_0873_),
    .Y(_0880_));
 sky130_fd_sc_hd__or2_1 _1514_ (.A(\MOS6502.ADD[2] ),
    .B(_0873_),
    .X(_0881_));
 sky130_fd_sc_hd__and3_1 _1515_ (.A(_0876_),
    .B(_0880_),
    .C(_0881_),
    .X(_0882_));
 sky130_fd_sc_hd__a21oi_1 _1516_ (.A1(_0880_),
    .A2(_0881_),
    .B1(_0876_),
    .Y(_0883_));
 sky130_fd_sc_hd__nand2_1 _1517_ (.A(_0450_),
    .B(_0585_),
    .Y(_0884_));
 sky130_fd_sc_hd__o31a_1 _1518_ (.A1(_0450_),
    .A2(_0882_),
    .A3(_0883_),
    .B1(_0884_),
    .X(_0885_));
 sky130_fd_sc_hd__and2b_1 _1519_ (.A_N(_0885_),
    .B(_0867_),
    .X(_0886_));
 sky130_fd_sc_hd__a22o_1 _1520_ (.A1(net159),
    .A2(_0870_),
    .B1(_0886_),
    .B2(_0868_),
    .X(_0010_));
 sky130_fd_sc_hd__a21o_1 _1521_ (.A1(\MOS6502.ADD[2] ),
    .A2(_0873_),
    .B1(_0882_),
    .X(_0887_));
 sky130_fd_sc_hd__xnor2_1 _1522_ (.A(\MOS6502.ADD[3] ),
    .B(_0875_),
    .Y(_0888_));
 sky130_fd_sc_hd__nor2_1 _1523_ (.A(_0887_),
    .B(_0888_),
    .Y(_0889_));
 sky130_fd_sc_hd__a21o_1 _1524_ (.A1(_0887_),
    .A2(_0888_),
    .B1(_0450_),
    .X(_0890_));
 sky130_fd_sc_hd__o221a_1 _1525_ (.A1(_0451_),
    .A2(_0577_),
    .B1(_0889_),
    .B2(_0890_),
    .C1(_0867_),
    .X(_0891_));
 sky130_fd_sc_hd__mux2_1 _1526_ (.A0(net127),
    .A1(_0891_),
    .S(_0869_),
    .X(_0011_));
 sky130_fd_sc_hd__or2_1 _1527_ (.A(_0451_),
    .B(_0570_),
    .X(_0892_));
 sky130_fd_sc_hd__o211a_1 _1528_ (.A1(\MOS6502.ADD[4] ),
    .A2(_0450_),
    .B1(_0867_),
    .C1(_0892_),
    .X(_0893_));
 sky130_fd_sc_hd__mux2_1 _1529_ (.A0(net135),
    .A1(_0893_),
    .S(_0869_),
    .X(_0012_));
 sky130_fd_sc_hd__and3_1 _1530_ (.A(\MOS6502.adc_bcd ),
    .B(\MOS6502.ALU.CO ),
    .C(\MOS6502.adj_bcd ),
    .X(_0894_));
 sky130_fd_sc_hd__o21ba_1 _1531_ (.A1(\MOS6502.ALU.CO ),
    .A2(_0874_),
    .B1_N(_0894_),
    .X(_0895_));
 sky130_fd_sc_hd__and2b_1 _1532_ (.A_N(_0895_),
    .B(\MOS6502.ADD[5] ),
    .X(_0896_));
 sky130_fd_sc_hd__xor2_1 _1533_ (.A(\MOS6502.ADD[5] ),
    .B(_0895_),
    .X(_0897_));
 sky130_fd_sc_hd__nand2_1 _1534_ (.A(_0451_),
    .B(_0897_),
    .Y(_0898_));
 sky130_fd_sc_hd__o211a_1 _1535_ (.A1(_0451_),
    .A2(_0564_),
    .B1(_0867_),
    .C1(_0898_),
    .X(_0899_));
 sky130_fd_sc_hd__mux2_1 _1536_ (.A0(net125),
    .A1(_0899_),
    .S(_0869_),
    .X(_0013_));
 sky130_fd_sc_hd__nand2_1 _1537_ (.A(\MOS6502.ADD[6] ),
    .B(_0894_),
    .Y(_0900_));
 sky130_fd_sc_hd__or2_1 _1538_ (.A(\MOS6502.ADD[6] ),
    .B(_0894_),
    .X(_0901_));
 sky130_fd_sc_hd__nand2_1 _1539_ (.A(_0900_),
    .B(_0901_),
    .Y(_0902_));
 sky130_fd_sc_hd__xnor2_1 _1540_ (.A(_0896_),
    .B(_0902_),
    .Y(_0903_));
 sky130_fd_sc_hd__mux2_1 _1541_ (.A0(_0558_),
    .A1(_0903_),
    .S(_0451_),
    .X(_0904_));
 sky130_fd_sc_hd__and2_1 _1542_ (.A(_0867_),
    .B(_0904_),
    .X(_0905_));
 sky130_fd_sc_hd__a22o_1 _1543_ (.A1(net151),
    .A2(_0870_),
    .B1(_0905_),
    .B2(_0868_),
    .X(_0014_));
 sky130_fd_sc_hd__a21bo_1 _1544_ (.A1(_0896_),
    .A2(_0901_),
    .B1_N(_0900_),
    .X(_0906_));
 sky130_fd_sc_hd__xnor2_1 _1545_ (.A(\MOS6502.ALU.CO ),
    .B(net244),
    .Y(_0907_));
 sky130_fd_sc_hd__mux2_1 _1546_ (.A0(_0907_),
    .A1(\MOS6502.ADD[7] ),
    .S(_0874_),
    .X(_0908_));
 sky130_fd_sc_hd__xnor2_1 _1547_ (.A(_0906_),
    .B(_0908_),
    .Y(_0909_));
 sky130_fd_sc_hd__nand2_1 _1548_ (.A(_0451_),
    .B(_0909_),
    .Y(_0910_));
 sky130_fd_sc_hd__o211a_1 _1549_ (.A1(_0451_),
    .A2(_0549_),
    .B1(_0867_),
    .C1(_0910_),
    .X(_0911_));
 sky130_fd_sc_hd__mux2_1 _1550_ (.A0(net105),
    .A1(_0911_),
    .S(_0869_),
    .X(_0015_));
 sky130_fd_sc_hd__and2_1 _1551_ (.A(net74),
    .B(net3),
    .X(_0016_));
 sky130_fd_sc_hd__and2_1 _1552_ (.A(net74),
    .B(net4),
    .X(_0017_));
 sky130_fd_sc_hd__and2_1 _1553_ (.A(net75),
    .B(net5),
    .X(_0018_));
 sky130_fd_sc_hd__and2_1 _1554_ (.A(net75),
    .B(net6),
    .X(_0019_));
 sky130_fd_sc_hd__and2_1 _1555_ (.A(net75),
    .B(net7),
    .X(_0020_));
 sky130_fd_sc_hd__and2_1 _1556_ (.A(net75),
    .B(net8),
    .X(_0021_));
 sky130_fd_sc_hd__and2_1 _1557_ (.A(net75),
    .B(net9),
    .X(_0022_));
 sky130_fd_sc_hd__and2_1 _1558_ (.A(net75),
    .B(net10),
    .X(_0023_));
 sky130_fd_sc_hd__a31o_4 _1559_ (.A1(_0490_),
    .A2(_0495_),
    .A3(_0866_),
    .B1(net72),
    .X(_0912_));
 sky130_fd_sc_hd__mux2_1 _1560_ (.A0(net161),
    .A1(_0872_),
    .S(_0912_),
    .X(_0024_));
 sky130_fd_sc_hd__mux2_1 _1561_ (.A0(net139),
    .A1(_0879_),
    .S(_0912_),
    .X(_0025_));
 sky130_fd_sc_hd__mux2_1 _1562_ (.A0(net143),
    .A1(_0886_),
    .S(_0912_),
    .X(_0026_));
 sky130_fd_sc_hd__mux2_1 _1563_ (.A0(net153),
    .A1(_0891_),
    .S(_0912_),
    .X(_0027_));
 sky130_fd_sc_hd__mux2_1 _1564_ (.A0(net99),
    .A1(_0893_),
    .S(_0912_),
    .X(_0028_));
 sky130_fd_sc_hd__mux2_1 _1565_ (.A0(net115),
    .A1(_0899_),
    .S(_0912_),
    .X(_0029_));
 sky130_fd_sc_hd__mux2_1 _1566_ (.A0(net103),
    .A1(_0905_),
    .S(_0912_),
    .X(_0030_));
 sky130_fd_sc_hd__mux2_1 _1567_ (.A0(net89),
    .A1(_0911_),
    .S(_0912_),
    .X(_0031_));
 sky130_fd_sc_hd__mux2_1 _1568_ (.A0(\MOS6502.backwards ),
    .A1(net192),
    .S(net78),
    .X(_0032_));
 sky130_fd_sc_hd__or2_1 _1569_ (.A(_0859_),
    .B(_0863_),
    .X(_0913_));
 sky130_fd_sc_hd__nand2_1 _1570_ (.A(_0859_),
    .B(_0863_),
    .Y(_0914_));
 sky130_fd_sc_hd__and2_1 _1571_ (.A(_0913_),
    .B(_0914_),
    .X(_0915_));
 sky130_fd_sc_hd__a22o_1 _1572_ (.A1(\MOS6502.ABH[6] ),
    .A2(net53),
    .B1(_0558_),
    .B2(_0839_),
    .X(_0916_));
 sky130_fd_sc_hd__a221o_1 _1573_ (.A1(\MOS6502.ADD[6] ),
    .A2(_0825_),
    .B1(_0837_),
    .B2(_0557_),
    .C1(_0916_),
    .X(_0917_));
 sky130_fd_sc_hd__a22o_1 _1574_ (.A1(\MOS6502.PC[6] ),
    .A2(_0723_),
    .B1(_0830_),
    .B2(_0558_),
    .X(_0918_));
 sky130_fd_sc_hd__a21oi_1 _1575_ (.A1(_0917_),
    .A2(_0918_),
    .B1(_0834_),
    .Y(_0919_));
 sky130_fd_sc_hd__a311o_1 _1576_ (.A1(_0843_),
    .A2(_0917_),
    .A3(_0918_),
    .B1(_0919_),
    .C1(_0845_),
    .X(_0920_));
 sky130_fd_sc_hd__a21oi_1 _1577_ (.A1(_0833_),
    .A2(_0918_),
    .B1(_0917_),
    .Y(_0921_));
 sky130_fd_sc_hd__nor2_1 _1578_ (.A(_0823_),
    .B(_0921_),
    .Y(_0922_));
 sky130_fd_sc_hd__a22o_1 _1579_ (.A1(_0823_),
    .A2(_0841_),
    .B1(_0920_),
    .B2(_0922_),
    .X(_0923_));
 sky130_fd_sc_hd__a21o_1 _1580_ (.A1(_0821_),
    .A2(_0923_),
    .B1(_0820_),
    .X(_0924_));
 sky130_fd_sc_hd__mux2_1 _1581_ (.A0(_0861_),
    .A1(_0821_),
    .S(_0918_),
    .X(_0925_));
 sky130_fd_sc_hd__and3_1 _1582_ (.A(_0923_),
    .B(_0924_),
    .C(_0925_),
    .X(_0926_));
 sky130_fd_sc_hd__a22o_1 _1583_ (.A1(\MOS6502.ABH[5] ),
    .A2(net53),
    .B1(_0564_),
    .B2(_0839_),
    .X(_0927_));
 sky130_fd_sc_hd__a221o_1 _1584_ (.A1(\MOS6502.ADD[5] ),
    .A2(_0825_),
    .B1(_0837_),
    .B2(_0563_),
    .C1(_0927_),
    .X(_0928_));
 sky130_fd_sc_hd__a22o_1 _1585_ (.A1(\MOS6502.PC[5] ),
    .A2(_0723_),
    .B1(_0830_),
    .B2(_0564_),
    .X(_0929_));
 sky130_fd_sc_hd__a21oi_1 _1586_ (.A1(_0928_),
    .A2(_0929_),
    .B1(_0834_),
    .Y(_0930_));
 sky130_fd_sc_hd__a31o_1 _1587_ (.A1(_0843_),
    .A2(_0928_),
    .A3(_0929_),
    .B1(_0845_),
    .X(_0931_));
 sky130_fd_sc_hd__a21o_1 _1588_ (.A1(_0833_),
    .A2(_0929_),
    .B1(_0928_),
    .X(_0932_));
 sky130_fd_sc_hd__o211a_1 _1589_ (.A1(_0930_),
    .A2(_0931_),
    .B1(_0932_),
    .C1(_0824_),
    .X(_0933_));
 sky130_fd_sc_hd__a21o_1 _1590_ (.A1(_0823_),
    .A2(_0917_),
    .B1(_0933_),
    .X(_0934_));
 sky130_fd_sc_hd__a21o_1 _1591_ (.A1(_0821_),
    .A2(_0934_),
    .B1(_0820_),
    .X(_0935_));
 sky130_fd_sc_hd__mux2_1 _1592_ (.A0(_0861_),
    .A1(_0821_),
    .S(_0929_),
    .X(_0936_));
 sky130_fd_sc_hd__and3_1 _1593_ (.A(_0934_),
    .B(_0935_),
    .C(_0936_),
    .X(_0937_));
 sky130_fd_sc_hd__a22o_1 _1594_ (.A1(\MOS6502.ABH[4] ),
    .A2(net53),
    .B1(_0570_),
    .B2(_0839_),
    .X(_0938_));
 sky130_fd_sc_hd__a221o_1 _1595_ (.A1(\MOS6502.ADD[4] ),
    .A2(_0825_),
    .B1(_0837_),
    .B2(_0569_),
    .C1(_0938_),
    .X(_0939_));
 sky130_fd_sc_hd__a22o_1 _1596_ (.A1(\MOS6502.PC[4] ),
    .A2(_0723_),
    .B1(_0830_),
    .B2(_0570_),
    .X(_0940_));
 sky130_fd_sc_hd__a21oi_1 _1597_ (.A1(_0939_),
    .A2(_0940_),
    .B1(_0834_),
    .Y(_0941_));
 sky130_fd_sc_hd__a31o_1 _1598_ (.A1(_0843_),
    .A2(_0939_),
    .A3(_0940_),
    .B1(_0845_),
    .X(_0942_));
 sky130_fd_sc_hd__a21o_1 _1599_ (.A1(_0833_),
    .A2(_0940_),
    .B1(_0939_),
    .X(_0943_));
 sky130_fd_sc_hd__o211a_1 _1600_ (.A1(_0941_),
    .A2(_0942_),
    .B1(_0943_),
    .C1(_0824_),
    .X(_0944_));
 sky130_fd_sc_hd__a21oi_1 _1601_ (.A1(_0823_),
    .A2(_0928_),
    .B1(_0944_),
    .Y(_0945_));
 sky130_fd_sc_hd__o21a_1 _1602_ (.A1(_0822_),
    .A2(_0945_),
    .B1(_0819_),
    .X(_0946_));
 sky130_fd_sc_hd__nor2_1 _1603_ (.A(_0861_),
    .B(_0940_),
    .Y(_0947_));
 sky130_fd_sc_hd__a211o_1 _1604_ (.A1(_0822_),
    .A2(_0940_),
    .B1(_0946_),
    .C1(_0947_),
    .X(_0948_));
 sky130_fd_sc_hd__nor2_1 _1605_ (.A(_0945_),
    .B(_0948_),
    .Y(_0949_));
 sky130_fd_sc_hd__and2_1 _1606_ (.A(_0945_),
    .B(_0948_),
    .X(_0950_));
 sky130_fd_sc_hd__nor2_1 _1607_ (.A(_0949_),
    .B(_0950_),
    .Y(_0951_));
 sky130_fd_sc_hd__a21o_1 _1608_ (.A1(_0582_),
    .A2(_0583_),
    .B1(_0838_),
    .X(_0952_));
 sky130_fd_sc_hd__a22o_1 _1609_ (.A1(\MOS6502.ABH[2] ),
    .A2(net53),
    .B1(_0585_),
    .B2(_0839_),
    .X(_0953_));
 sky130_fd_sc_hd__a21oi_1 _1610_ (.A1(\MOS6502.ADD[2] ),
    .A2(_0825_),
    .B1(_0953_),
    .Y(_0954_));
 sky130_fd_sc_hd__nand2_1 _1611_ (.A(_0952_),
    .B(_0954_),
    .Y(_0955_));
 sky130_fd_sc_hd__a22o_1 _1612_ (.A1(\MOS6502.PC[2] ),
    .A2(_0723_),
    .B1(_0830_),
    .B2(_0585_),
    .X(_0956_));
 sky130_fd_sc_hd__inv_2 _1613_ (.A(_0956_),
    .Y(_0957_));
 sky130_fd_sc_hd__a21o_1 _1614_ (.A1(_0952_),
    .A2(_0954_),
    .B1(_0957_),
    .X(_0958_));
 sky130_fd_sc_hd__a211oi_1 _1615_ (.A1(_0952_),
    .A2(_0954_),
    .B1(_0957_),
    .C1(_0844_),
    .Y(_0959_));
 sky130_fd_sc_hd__a211o_1 _1616_ (.A1(_0833_),
    .A2(_0958_),
    .B1(_0959_),
    .C1(_0845_),
    .X(_0960_));
 sky130_fd_sc_hd__nor2_1 _1617_ (.A(_0834_),
    .B(_0957_),
    .Y(_0961_));
 sky130_fd_sc_hd__o21a_1 _1618_ (.A1(_0955_),
    .A2(_0961_),
    .B1(_0824_),
    .X(_0962_));
 sky130_fd_sc_hd__o211ai_4 _1619_ (.A1(_0490_),
    .A2(_0574_),
    .B1(_0575_),
    .C1(_0837_),
    .Y(_0963_));
 sky130_fd_sc_hd__a22o_1 _1620_ (.A1(\MOS6502.ABH[3] ),
    .A2(net53),
    .B1(_0577_),
    .B2(_0839_),
    .X(_0964_));
 sky130_fd_sc_hd__a21oi_1 _1621_ (.A1(\MOS6502.ADD[3] ),
    .A2(_0825_),
    .B1(_0964_),
    .Y(_0965_));
 sky130_fd_sc_hd__nand2_1 _1622_ (.A(_0963_),
    .B(_0965_),
    .Y(_0966_));
 sky130_fd_sc_hd__a22o_1 _1623_ (.A1(_0960_),
    .A2(_0962_),
    .B1(_0966_),
    .B2(_0823_),
    .X(_0967_));
 sky130_fd_sc_hd__a21o_1 _1624_ (.A1(_0821_),
    .A2(_0967_),
    .B1(_0820_),
    .X(_0968_));
 sky130_fd_sc_hd__mux2_1 _1625_ (.A0(_0861_),
    .A1(_0821_),
    .S(_0956_),
    .X(_0969_));
 sky130_fd_sc_hd__and3_1 _1626_ (.A(_0967_),
    .B(_0968_),
    .C(_0969_),
    .X(_0970_));
 sky130_fd_sc_hd__a21oi_1 _1627_ (.A1(_0968_),
    .A2(_0969_),
    .B1(_0967_),
    .Y(_0971_));
 sky130_fd_sc_hd__nor2_1 _1628_ (.A(_0970_),
    .B(_0971_),
    .Y(_0972_));
 sky130_fd_sc_hd__a22o_1 _1629_ (.A1(\MOS6502.ABH[1] ),
    .A2(net53),
    .B1(_0591_),
    .B2(_0839_),
    .X(_0973_));
 sky130_fd_sc_hd__a221o_1 _1630_ (.A1(\MOS6502.ADD[1] ),
    .A2(_0825_),
    .B1(_0837_),
    .B2(_0590_),
    .C1(_0973_),
    .X(_0974_));
 sky130_fd_sc_hd__a22oi_4 _1631_ (.A1(\MOS6502.PC[1] ),
    .A2(_0723_),
    .B1(_0830_),
    .B2(_0591_),
    .Y(_0975_));
 sky130_fd_sc_hd__or3b_1 _1632_ (.A(_0833_),
    .B(_0844_),
    .C_N(_0975_),
    .X(_0976_));
 sky130_fd_sc_hd__nor2_1 _1633_ (.A(_0834_),
    .B(_0975_),
    .Y(_0977_));
 sky130_fd_sc_hd__o31a_1 _1634_ (.A1(_0834_),
    .A2(_0842_),
    .A3(_0975_),
    .B1(_0976_),
    .X(_0978_));
 sky130_fd_sc_hd__mux2_1 _1635_ (.A0(_0977_),
    .A1(_0978_),
    .S(_0974_),
    .X(_0979_));
 sky130_fd_sc_hd__mux2_1 _1636_ (.A0(_0955_),
    .A1(_0979_),
    .S(_0824_),
    .X(_0980_));
 sky130_fd_sc_hd__a21o_1 _1637_ (.A1(_0821_),
    .A2(_0980_),
    .B1(_0820_),
    .X(_0981_));
 sky130_fd_sc_hd__mux2_1 _1638_ (.A0(_0821_),
    .A1(_0861_),
    .S(_0975_),
    .X(_0982_));
 sky130_fd_sc_hd__and3_1 _1639_ (.A(_0980_),
    .B(_0981_),
    .C(_0982_),
    .X(_0983_));
 sky130_fd_sc_hd__a21oi_1 _1640_ (.A1(_0596_),
    .A2(_0597_),
    .B1(_0838_),
    .Y(_0984_));
 sky130_fd_sc_hd__a22o_1 _1641_ (.A1(\MOS6502.ABH[0] ),
    .A2(net53),
    .B1(_0599_),
    .B2(_0839_),
    .X(_0985_));
 sky130_fd_sc_hd__a21o_1 _1642_ (.A1(\MOS6502.ADD[0] ),
    .A2(_0825_),
    .B1(_0985_),
    .X(_0986_));
 sky130_fd_sc_hd__or2_1 _1643_ (.A(_0984_),
    .B(_0986_),
    .X(_0987_));
 sky130_fd_sc_hd__a22o_1 _1644_ (.A1(\MOS6502.PC[0] ),
    .A2(_0723_),
    .B1(_0830_),
    .B2(_0599_),
    .X(_0988_));
 sky130_fd_sc_hd__o21a_1 _1645_ (.A1(_0984_),
    .A2(_0986_),
    .B1(_0988_),
    .X(_0989_));
 sky130_fd_sc_hd__a21o_1 _1646_ (.A1(_0843_),
    .A2(_0988_),
    .B1(_0845_),
    .X(_0990_));
 sky130_fd_sc_hd__o2bb2a_1 _1647_ (.A1_N(_0987_),
    .A2_N(_0990_),
    .B1(_0989_),
    .B2(_0834_),
    .X(_0991_));
 sky130_fd_sc_hd__o21ai_1 _1648_ (.A1(_0987_),
    .A2(_0988_),
    .B1(_0824_),
    .Y(_0992_));
 sky130_fd_sc_hd__o2bb2a_1 _1649_ (.A1_N(_0823_),
    .A2_N(_0974_),
    .B1(_0991_),
    .B2(_0992_),
    .X(_0993_));
 sky130_fd_sc_hd__nand2_1 _1650_ (.A(_0819_),
    .B(_0822_),
    .Y(_0994_));
 sky130_fd_sc_hd__nand2_1 _1651_ (.A(_0861_),
    .B(_0994_),
    .Y(_0995_));
 sky130_fd_sc_hd__mux2_1 _1652_ (.A0(_0995_),
    .A1(_0822_),
    .S(_0988_),
    .X(_0996_));
 sky130_fd_sc_hd__nor2_1 _1653_ (.A(_0993_),
    .B(_0996_),
    .Y(_0997_));
 sky130_fd_sc_hd__and3_1 _1654_ (.A(_0824_),
    .B(_0858_),
    .C(_0994_),
    .X(_0998_));
 sky130_fd_sc_hd__o21ai_1 _1655_ (.A1(_0819_),
    .A2(_0996_),
    .B1(_0993_),
    .Y(_0999_));
 sky130_fd_sc_hd__nand2b_1 _1656_ (.A_N(_0997_),
    .B(_0999_),
    .Y(_1000_));
 sky130_fd_sc_hd__a21o_1 _1657_ (.A1(_0998_),
    .A2(_0999_),
    .B1(_0997_),
    .X(_1001_));
 sky130_fd_sc_hd__a21o_1 _1658_ (.A1(_0981_),
    .A2(_0982_),
    .B1(_0980_),
    .X(_1002_));
 sky130_fd_sc_hd__nand2b_1 _1659_ (.A_N(_0983_),
    .B(_1002_),
    .Y(_1003_));
 sky130_fd_sc_hd__a21o_1 _1660_ (.A1(_1001_),
    .A2(_1002_),
    .B1(_0983_),
    .X(_1004_));
 sky130_fd_sc_hd__and2_1 _1661_ (.A(_0972_),
    .B(_1004_),
    .X(_1005_));
 sky130_fd_sc_hd__xor2_1 _1662_ (.A(_0972_),
    .B(_1004_),
    .X(_1006_));
 sky130_fd_sc_hd__xnor2_1 _1663_ (.A(_1001_),
    .B(_1003_),
    .Y(_1007_));
 sky130_fd_sc_hd__a22o_1 _1664_ (.A1(\MOS6502.PC[3] ),
    .A2(_0723_),
    .B1(_0830_),
    .B2(_0577_),
    .X(_1008_));
 sky130_fd_sc_hd__inv_2 _1665_ (.A(_1008_),
    .Y(_1009_));
 sky130_fd_sc_hd__a21o_1 _1666_ (.A1(_0963_),
    .A2(_0965_),
    .B1(_1009_),
    .X(_1010_));
 sky130_fd_sc_hd__a211oi_1 _1667_ (.A1(_0963_),
    .A2(_0965_),
    .B1(_1009_),
    .C1(_0844_),
    .Y(_1011_));
 sky130_fd_sc_hd__a211o_1 _1668_ (.A1(_0833_),
    .A2(_1010_),
    .B1(_1011_),
    .C1(_0845_),
    .X(_1012_));
 sky130_fd_sc_hd__nor2_1 _1669_ (.A(_0834_),
    .B(_1009_),
    .Y(_1013_));
 sky130_fd_sc_hd__o21a_1 _1670_ (.A1(_0966_),
    .A2(_1013_),
    .B1(_0824_),
    .X(_1014_));
 sky130_fd_sc_hd__a22o_1 _1671_ (.A1(_0823_),
    .A2(_0939_),
    .B1(_1012_),
    .B2(_1014_),
    .X(_1015_));
 sky130_fd_sc_hd__a21o_1 _1672_ (.A1(_0821_),
    .A2(_1015_),
    .B1(_0820_),
    .X(_1016_));
 sky130_fd_sc_hd__mux2_1 _1673_ (.A0(_0861_),
    .A1(_0821_),
    .S(_1008_),
    .X(_1017_));
 sky130_fd_sc_hd__and3_1 _1674_ (.A(_1015_),
    .B(_1016_),
    .C(_1017_),
    .X(_1018_));
 sky130_fd_sc_hd__a21oi_1 _1675_ (.A1(_1016_),
    .A2(_1017_),
    .B1(_1015_),
    .Y(_1019_));
 sky130_fd_sc_hd__nor2_1 _1676_ (.A(_1018_),
    .B(_1019_),
    .Y(_1020_));
 sky130_fd_sc_hd__a211o_1 _1677_ (.A1(_0972_),
    .A2(_1004_),
    .B1(_1020_),
    .C1(_0970_),
    .X(_1021_));
 sky130_fd_sc_hd__o2111a_1 _1678_ (.A1(_1006_),
    .A2(_1007_),
    .B1(_1021_),
    .C1(_0630_),
    .D1(\MOS6502.adc_bcd ),
    .X(_1022_));
 sky130_fd_sc_hd__o21a_1 _1679_ (.A1(_0970_),
    .A2(_1005_),
    .B1(_1020_),
    .X(_1023_));
 sky130_fd_sc_hd__or3_1 _1680_ (.A(_1018_),
    .B(_1022_),
    .C(_1023_),
    .X(_1024_));
 sky130_fd_sc_hd__o31a_1 _1681_ (.A1(_1018_),
    .A2(_1022_),
    .A3(_1023_),
    .B1(_0951_),
    .X(_0151_));
 sky130_fd_sc_hd__a21oi_1 _1682_ (.A1(_0935_),
    .A2(_0936_),
    .B1(_0934_),
    .Y(_0152_));
 sky130_fd_sc_hd__nor2_1 _1683_ (.A(_0937_),
    .B(_0152_),
    .Y(_0153_));
 sky130_fd_sc_hd__o21a_1 _1684_ (.A1(_0949_),
    .A2(_0151_),
    .B1(_0153_),
    .X(_0154_));
 sky130_fd_sc_hd__a21oi_1 _1685_ (.A1(_0924_),
    .A2(_0925_),
    .B1(_0923_),
    .Y(_0155_));
 sky130_fd_sc_hd__nor2_1 _1686_ (.A(_0926_),
    .B(_0155_),
    .Y(_0156_));
 sky130_fd_sc_hd__o21a_1 _1687_ (.A1(_0937_),
    .A2(_0154_),
    .B1(_0156_),
    .X(_0157_));
 sky130_fd_sc_hd__o21ai_1 _1688_ (.A1(_0926_),
    .A2(_0157_),
    .B1(_0915_),
    .Y(_0158_));
 sky130_fd_sc_hd__or3_1 _1689_ (.A(_0915_),
    .B(_0926_),
    .C(_0157_),
    .X(_0159_));
 sky130_fd_sc_hd__and2_1 _1690_ (.A(_0158_),
    .B(_0159_),
    .X(_0160_));
 sky130_fd_sc_hd__nor3_1 _1691_ (.A(_0949_),
    .B(_0151_),
    .C(_0153_),
    .Y(_0161_));
 sky130_fd_sc_hd__nor2_1 _1692_ (.A(_0154_),
    .B(_0161_),
    .Y(_0162_));
 sky130_fd_sc_hd__nor3_1 _1693_ (.A(_0937_),
    .B(_0154_),
    .C(_0156_),
    .Y(_0163_));
 sky130_fd_sc_hd__nor2_1 _1694_ (.A(_0157_),
    .B(_0163_),
    .Y(_0164_));
 sky130_fd_sc_hd__o211a_1 _1695_ (.A1(_0162_),
    .A2(_0164_),
    .B1(\MOS6502.adc_bcd ),
    .C1(_0630_),
    .X(_0165_));
 sky130_fd_sc_hd__a22oi_1 _1696_ (.A1(_0823_),
    .A2(_0987_),
    .B1(_0158_),
    .B2(_0913_),
    .Y(_0166_));
 sky130_fd_sc_hd__and4_1 _1697_ (.A(_0823_),
    .B(_0913_),
    .C(_0987_),
    .D(_0158_),
    .X(_0167_));
 sky130_fd_sc_hd__a211o_1 _1698_ (.A1(_0160_),
    .A2(_0165_),
    .B1(_0166_),
    .C1(_0167_),
    .X(_0168_));
 sky130_fd_sc_hd__mux2_1 _1699_ (.A0(net275),
    .A1(_0168_),
    .S(net79),
    .X(_0033_));
 sky130_fd_sc_hd__mux2_1 _1700_ (.A0(net173),
    .A1(_1024_),
    .S(net79),
    .X(_0034_));
 sky130_fd_sc_hd__xnor2_1 _1701_ (.A(_0998_),
    .B(_1000_),
    .Y(_0169_));
 sky130_fd_sc_hd__mux2_1 _1702_ (.A0(net259),
    .A1(_0169_),
    .S(net79),
    .X(_0035_));
 sky130_fd_sc_hd__mux2_1 _1703_ (.A0(net261),
    .A1(_1007_),
    .S(net79),
    .X(_0036_));
 sky130_fd_sc_hd__mux2_1 _1704_ (.A0(net284),
    .A1(_1006_),
    .S(net79),
    .X(_0037_));
 sky130_fd_sc_hd__nor2_1 _1705_ (.A(_0429_),
    .B(_1023_),
    .Y(_0170_));
 sky130_fd_sc_hd__a22o_1 _1706_ (.A1(_0429_),
    .A2(net278),
    .B1(_1021_),
    .B2(_0170_),
    .X(_0038_));
 sky130_fd_sc_hd__nor2_1 _1707_ (.A(_0951_),
    .B(_1024_),
    .Y(_0171_));
 sky130_fd_sc_hd__or2_1 _1708_ (.A(_0429_),
    .B(_0151_),
    .X(_0172_));
 sky130_fd_sc_hd__a2bb2o_1 _1709_ (.A1_N(_0172_),
    .A2_N(_0171_),
    .B1(net255),
    .B2(_0429_),
    .X(_0039_));
 sky130_fd_sc_hd__mux2_1 _1710_ (.A0(net264),
    .A1(_0162_),
    .S(net79),
    .X(_0040_));
 sky130_fd_sc_hd__mux2_1 _1711_ (.A0(net277),
    .A1(_0164_),
    .S(net79),
    .X(_0041_));
 sky130_fd_sc_hd__mux2_1 _1712_ (.A0(net244),
    .A1(_0160_),
    .S(net79),
    .X(_0042_));
 sky130_fd_sc_hd__mux2_1 _1713_ (.A0(net175),
    .A1(_0841_),
    .S(net79),
    .X(_0043_));
 sky130_fd_sc_hd__o22a_1 _1714_ (.A1(_0443_),
    .A2(_0447_),
    .B1(_0500_),
    .B2(_0621_),
    .X(_0173_));
 sky130_fd_sc_hd__or2_4 _1715_ (.A(_0521_),
    .B(_0173_),
    .X(_0174_));
 sky130_fd_sc_hd__or3_4 _1716_ (.A(_0521_),
    .B(_0527_),
    .C(_0173_),
    .X(_0175_));
 sky130_fd_sc_hd__nor3_2 _1717_ (.A(net55),
    .B(net54),
    .C(_0175_),
    .Y(_0176_));
 sky130_fd_sc_hd__and2_1 _1718_ (.A(net55),
    .B(net52),
    .X(_0177_));
 sky130_fd_sc_hd__o21a_1 _1719_ (.A1(_0176_),
    .A2(_0177_),
    .B1(net223),
    .X(_0178_));
 sky130_fd_sc_hd__nor2_2 _1720_ (.A(_0477_),
    .B(net52),
    .Y(_0179_));
 sky130_fd_sc_hd__a22o_1 _1721_ (.A1(\MOS6502.ADD[0] ),
    .A2(_0175_),
    .B1(_0179_),
    .B2(\MOS6502.ABL[0] ),
    .X(_0180_));
 sky130_fd_sc_hd__a2111o_1 _1722_ (.A1(_0443_),
    .A2(_0621_),
    .B1(_0723_),
    .C1(_0465_),
    .D1(_0485_),
    .X(_0181_));
 sky130_fd_sc_hd__or3_1 _1723_ (.A(_0516_),
    .B(_0524_),
    .C(_0181_),
    .X(_0182_));
 sky130_fd_sc_hd__or4_1 _1724_ (.A(_0729_),
    .B(_0763_),
    .C(_0177_),
    .D(_0182_),
    .X(_0183_));
 sky130_fd_sc_hd__o21ai_1 _1725_ (.A1(_0178_),
    .A2(_0180_),
    .B1(_0183_),
    .Y(_0184_));
 sky130_fd_sc_hd__or3_1 _1726_ (.A(_0178_),
    .B(_0180_),
    .C(_0183_),
    .X(_0185_));
 sky130_fd_sc_hd__a32o_1 _1727_ (.A1(_0620_),
    .A2(_0184_),
    .A3(_0185_),
    .B1(net60),
    .B2(net223),
    .X(_0044_));
 sky130_fd_sc_hd__nand2_1 _1728_ (.A(net219),
    .B(net52),
    .Y(_0186_));
 sky130_fd_sc_hd__a211o_1 _1729_ (.A1(_0535_),
    .A2(_0176_),
    .B1(net52),
    .C1(_0438_),
    .X(_0187_));
 sky130_fd_sc_hd__a21o_1 _1730_ (.A1(_0186_),
    .A2(_0187_),
    .B1(_0477_),
    .X(_0188_));
 sky130_fd_sc_hd__a22oi_2 _1731_ (.A1(_0437_),
    .A2(net54),
    .B1(_0175_),
    .B2(\MOS6502.ADD[1] ),
    .Y(_0189_));
 sky130_fd_sc_hd__nand2_1 _1732_ (.A(net219),
    .B(_0176_),
    .Y(_0190_));
 sky130_fd_sc_hd__a31o_1 _1733_ (.A1(_0188_),
    .A2(_0189_),
    .A3(_0190_),
    .B1(_0184_),
    .X(_0191_));
 sky130_fd_sc_hd__and4_1 _1734_ (.A(_0184_),
    .B(_0188_),
    .C(_0189_),
    .D(_0190_),
    .X(_0192_));
 sky130_fd_sc_hd__nand2_1 _1735_ (.A(_0620_),
    .B(_0191_),
    .Y(_0193_));
 sky130_fd_sc_hd__a2bb2o_1 _1736_ (.A1_N(_0192_),
    .A2_N(_0193_),
    .B1(net219),
    .B2(net60),
    .X(_0045_));
 sky130_fd_sc_hd__o21ai_1 _1737_ (.A1(_0176_),
    .A2(_0177_),
    .B1(net217),
    .Y(_0194_));
 sky130_fd_sc_hd__o21a_1 _1738_ (.A1(_0428_),
    .A2(net177),
    .B1(_0509_),
    .X(_0195_));
 sky130_fd_sc_hd__a21oi_1 _1739_ (.A1(\MOS6502.ABL[2] ),
    .A2(_0179_),
    .B1(_0195_),
    .Y(_0196_));
 sky130_fd_sc_hd__nand2_1 _1740_ (.A(\MOS6502.ADD[2] ),
    .B(_0175_),
    .Y(_0197_));
 sky130_fd_sc_hd__a31o_1 _1741_ (.A1(_0194_),
    .A2(_0196_),
    .A3(_0197_),
    .B1(_0191_),
    .X(_0198_));
 sky130_fd_sc_hd__nand4_1 _1742_ (.A(_0191_),
    .B(_0194_),
    .C(_0196_),
    .D(_0197_),
    .Y(_0199_));
 sky130_fd_sc_hd__a32o_1 _1743_ (.A1(net64),
    .A2(_0198_),
    .A3(_0199_),
    .B1(net60),
    .B2(net217),
    .X(_0046_));
 sky130_fd_sc_hd__o21bai_4 _1744_ (.A1(net55),
    .A2(_0175_),
    .B1_N(_0177_),
    .Y(_0200_));
 sky130_fd_sc_hd__nand2_1 _1745_ (.A(net213),
    .B(_0200_),
    .Y(_0201_));
 sky130_fd_sc_hd__a21oi_1 _1746_ (.A1(\MOS6502.ABL[3] ),
    .A2(_0179_),
    .B1(net54),
    .Y(_0202_));
 sky130_fd_sc_hd__nand2_1 _1747_ (.A(\MOS6502.ADD[3] ),
    .B(_0175_),
    .Y(_0203_));
 sky130_fd_sc_hd__a31o_1 _1748_ (.A1(_0201_),
    .A2(_0202_),
    .A3(_0203_),
    .B1(_0198_),
    .X(_0204_));
 sky130_fd_sc_hd__nand4_1 _1749_ (.A(_0198_),
    .B(_0201_),
    .C(_0202_),
    .D(_0203_),
    .Y(_0205_));
 sky130_fd_sc_hd__a32o_1 _1750_ (.A1(net64),
    .A2(_0204_),
    .A3(_0205_),
    .B1(net60),
    .B2(net213),
    .X(_0047_));
 sky130_fd_sc_hd__nand2_1 _1751_ (.A(net221),
    .B(_0200_),
    .Y(_0206_));
 sky130_fd_sc_hd__a21oi_1 _1752_ (.A1(\MOS6502.ABL[4] ),
    .A2(_0179_),
    .B1(net54),
    .Y(_0207_));
 sky130_fd_sc_hd__nand2_1 _1753_ (.A(\MOS6502.ADD[4] ),
    .B(_0175_),
    .Y(_0208_));
 sky130_fd_sc_hd__a31o_1 _1754_ (.A1(_0206_),
    .A2(_0207_),
    .A3(_0208_),
    .B1(_0204_),
    .X(_0209_));
 sky130_fd_sc_hd__nand4_1 _1755_ (.A(_0204_),
    .B(_0206_),
    .C(_0207_),
    .D(_0208_),
    .Y(_0210_));
 sky130_fd_sc_hd__a32o_1 _1756_ (.A1(net64),
    .A2(_0209_),
    .A3(_0210_),
    .B1(net60),
    .B2(net221),
    .X(_0048_));
 sky130_fd_sc_hd__nand2_1 _1757_ (.A(net225),
    .B(_0200_),
    .Y(_0211_));
 sky130_fd_sc_hd__a21oi_1 _1758_ (.A1(\MOS6502.ABL[5] ),
    .A2(_0179_),
    .B1(net54),
    .Y(_0212_));
 sky130_fd_sc_hd__nand2_1 _1759_ (.A(\MOS6502.ADD[5] ),
    .B(_0175_),
    .Y(_0213_));
 sky130_fd_sc_hd__nand4_1 _1760_ (.A(_0209_),
    .B(_0211_),
    .C(_0212_),
    .D(_0213_),
    .Y(_0214_));
 sky130_fd_sc_hd__a31o_1 _1761_ (.A1(_0211_),
    .A2(_0212_),
    .A3(_0213_),
    .B1(_0209_),
    .X(_0215_));
 sky130_fd_sc_hd__a32o_1 _1762_ (.A1(net64),
    .A2(_0214_),
    .A3(_0215_),
    .B1(net60),
    .B2(net225),
    .X(_0049_));
 sky130_fd_sc_hd__nand2_1 _1763_ (.A(net211),
    .B(_0200_),
    .Y(_0216_));
 sky130_fd_sc_hd__a21oi_1 _1764_ (.A1(\MOS6502.ABL[6] ),
    .A2(_0179_),
    .B1(net54),
    .Y(_0217_));
 sky130_fd_sc_hd__nand2_1 _1765_ (.A(\MOS6502.ADD[6] ),
    .B(_0175_),
    .Y(_0218_));
 sky130_fd_sc_hd__a31o_1 _1766_ (.A1(_0216_),
    .A2(_0217_),
    .A3(_0218_),
    .B1(_0215_),
    .X(_0219_));
 sky130_fd_sc_hd__nand4_1 _1767_ (.A(_0215_),
    .B(_0216_),
    .C(_0217_),
    .D(_0218_),
    .Y(_0220_));
 sky130_fd_sc_hd__a32o_1 _1768_ (.A1(net64),
    .A2(_0219_),
    .A3(_0220_),
    .B1(net60),
    .B2(net211),
    .X(_0050_));
 sky130_fd_sc_hd__a221o_1 _1769_ (.A1(\MOS6502.ADD[7] ),
    .A2(_0175_),
    .B1(_0179_),
    .B2(\MOS6502.ABL[7] ),
    .C1(net54),
    .X(_0221_));
 sky130_fd_sc_hd__a21oi_1 _1770_ (.A1(net209),
    .A2(_0200_),
    .B1(_0221_),
    .Y(_0222_));
 sky130_fd_sc_hd__nand2_1 _1771_ (.A(_0219_),
    .B(_0222_),
    .Y(_0223_));
 sky130_fd_sc_hd__or2_1 _1772_ (.A(_0219_),
    .B(_0222_),
    .X(_0224_));
 sky130_fd_sc_hd__a32o_1 _1773_ (.A1(net64),
    .A2(_0223_),
    .A3(_0224_),
    .B1(net60),
    .B2(net209),
    .X(_0051_));
 sky130_fd_sc_hd__a21o_2 _1774_ (.A1(_0535_),
    .A2(_0176_),
    .B1(_0177_),
    .X(_0225_));
 sky130_fd_sc_hd__nand2_1 _1775_ (.A(net184),
    .B(_0225_),
    .Y(_0226_));
 sky130_fd_sc_hd__or2_4 _1776_ (.A(net53),
    .B(_0179_),
    .X(_0227_));
 sky130_fd_sc_hd__a221oi_2 _1777_ (.A1(\MOS6502.ADD[0] ),
    .A2(_0534_),
    .B1(_0227_),
    .B2(\MOS6502.ABH[0] ),
    .C1(net54),
    .Y(_0228_));
 sky130_fd_sc_hd__nand2_1 _1778_ (.A(_0599_),
    .B(_0174_),
    .Y(_0229_));
 sky130_fd_sc_hd__a31o_1 _1779_ (.A1(_0226_),
    .A2(_0228_),
    .A3(_0229_),
    .B1(_0224_),
    .X(_0230_));
 sky130_fd_sc_hd__nand4_1 _1780_ (.A(_0224_),
    .B(_0226_),
    .C(_0228_),
    .D(_0229_),
    .Y(_0231_));
 sky130_fd_sc_hd__a32o_1 _1781_ (.A1(net64),
    .A2(_0230_),
    .A3(_0231_),
    .B1(net60),
    .B2(net184),
    .X(_0052_));
 sky130_fd_sc_hd__nand2_1 _1782_ (.A(net182),
    .B(_0225_),
    .Y(_0232_));
 sky130_fd_sc_hd__a221oi_2 _1783_ (.A1(\MOS6502.ADD[1] ),
    .A2(_0534_),
    .B1(_0227_),
    .B2(\MOS6502.ABH[1] ),
    .C1(net54),
    .Y(_0233_));
 sky130_fd_sc_hd__nand2_1 _1784_ (.A(_0591_),
    .B(_0174_),
    .Y(_0234_));
 sky130_fd_sc_hd__nand4_1 _1785_ (.A(_0230_),
    .B(_0232_),
    .C(_0233_),
    .D(_0234_),
    .Y(_0235_));
 sky130_fd_sc_hd__a31o_1 _1786_ (.A1(_0232_),
    .A2(_0233_),
    .A3(_0234_),
    .B1(_0230_),
    .X(_0236_));
 sky130_fd_sc_hd__a32o_1 _1787_ (.A1(net64),
    .A2(_0235_),
    .A3(_0236_),
    .B1(net60),
    .B2(net182),
    .X(_0053_));
 sky130_fd_sc_hd__nand2_1 _1788_ (.A(net188),
    .B(_0225_),
    .Y(_0237_));
 sky130_fd_sc_hd__a221oi_2 _1789_ (.A1(\MOS6502.ADD[2] ),
    .A2(_0534_),
    .B1(_0227_),
    .B2(\MOS6502.ABH[2] ),
    .C1(net54),
    .Y(_0238_));
 sky130_fd_sc_hd__nand2_1 _1790_ (.A(_0585_),
    .B(_0174_),
    .Y(_0239_));
 sky130_fd_sc_hd__a31o_1 _1791_ (.A1(_0237_),
    .A2(_0238_),
    .A3(_0239_),
    .B1(_0236_),
    .X(_0240_));
 sky130_fd_sc_hd__nand4_1 _1792_ (.A(_0236_),
    .B(_0237_),
    .C(_0238_),
    .D(_0239_),
    .Y(_0241_));
 sky130_fd_sc_hd__a32o_1 _1793_ (.A1(net64),
    .A2(_0240_),
    .A3(_0241_),
    .B1(net60),
    .B2(net188),
    .X(_0054_));
 sky130_fd_sc_hd__nand2_1 _1794_ (.A(net194),
    .B(_0225_),
    .Y(_0242_));
 sky130_fd_sc_hd__a221oi_2 _1795_ (.A1(\MOS6502.ADD[3] ),
    .A2(_0534_),
    .B1(_0227_),
    .B2(\MOS6502.ABH[3] ),
    .C1(net54),
    .Y(_0243_));
 sky130_fd_sc_hd__nand2_1 _1796_ (.A(_0577_),
    .B(_0174_),
    .Y(_0244_));
 sky130_fd_sc_hd__nand4_1 _1797_ (.A(_0240_),
    .B(_0242_),
    .C(_0243_),
    .D(_0244_),
    .Y(_0245_));
 sky130_fd_sc_hd__a31o_1 _1798_ (.A1(_0242_),
    .A2(_0243_),
    .A3(_0244_),
    .B1(_0240_),
    .X(_0246_));
 sky130_fd_sc_hd__a32o_1 _1799_ (.A1(net64),
    .A2(_0245_),
    .A3(_0246_),
    .B1(net60),
    .B2(net194),
    .X(_0055_));
 sky130_fd_sc_hd__nand2_1 _1800_ (.A(net190),
    .B(_0225_),
    .Y(_0247_));
 sky130_fd_sc_hd__a221oi_2 _1801_ (.A1(\MOS6502.ADD[4] ),
    .A2(_0534_),
    .B1(_0227_),
    .B2(\MOS6502.ABH[4] ),
    .C1(net54),
    .Y(_0248_));
 sky130_fd_sc_hd__nand2_1 _1802_ (.A(_0570_),
    .B(_0174_),
    .Y(_0249_));
 sky130_fd_sc_hd__a31o_1 _1803_ (.A1(_0247_),
    .A2(_0248_),
    .A3(_0249_),
    .B1(_0246_),
    .X(_0250_));
 sky130_fd_sc_hd__nand4_1 _1804_ (.A(_0246_),
    .B(_0247_),
    .C(_0248_),
    .D(_0249_),
    .Y(_0251_));
 sky130_fd_sc_hd__a32o_1 _1805_ (.A1(net64),
    .A2(_0250_),
    .A3(_0251_),
    .B1(net60),
    .B2(net190),
    .X(_0056_));
 sky130_fd_sc_hd__nand2_1 _1806_ (.A(net196),
    .B(_0225_),
    .Y(_0252_));
 sky130_fd_sc_hd__a221oi_2 _1807_ (.A1(\MOS6502.ADD[5] ),
    .A2(_0534_),
    .B1(_0227_),
    .B2(\MOS6502.ABH[5] ),
    .C1(net54),
    .Y(_0253_));
 sky130_fd_sc_hd__nand2_1 _1808_ (.A(_0564_),
    .B(_0174_),
    .Y(_0254_));
 sky130_fd_sc_hd__nand4_1 _1809_ (.A(_0250_),
    .B(_0252_),
    .C(_0253_),
    .D(_0254_),
    .Y(_0255_));
 sky130_fd_sc_hd__a31o_1 _1810_ (.A1(_0252_),
    .A2(_0253_),
    .A3(_0254_),
    .B1(_0250_),
    .X(_0256_));
 sky130_fd_sc_hd__a32o_1 _1811_ (.A1(net64),
    .A2(_0255_),
    .A3(_0256_),
    .B1(net60),
    .B2(net196),
    .X(_0057_));
 sky130_fd_sc_hd__a221o_1 _1812_ (.A1(\MOS6502.ADD[6] ),
    .A2(_0534_),
    .B1(_0227_),
    .B2(\MOS6502.ABH[6] ),
    .C1(net54),
    .X(_0257_));
 sky130_fd_sc_hd__a221oi_2 _1813_ (.A1(_0558_),
    .A2(_0174_),
    .B1(_0225_),
    .B2(net202),
    .C1(_0257_),
    .Y(_0258_));
 sky130_fd_sc_hd__or2_1 _1814_ (.A(_0256_),
    .B(_0258_),
    .X(_0259_));
 sky130_fd_sc_hd__a21boi_1 _1815_ (.A1(_0256_),
    .A2(_0258_),
    .B1_N(net64),
    .Y(_0260_));
 sky130_fd_sc_hd__a22o_1 _1816_ (.A1(net202),
    .A2(net60),
    .B1(_0259_),
    .B2(_0260_),
    .X(_0058_));
 sky130_fd_sc_hd__a221o_1 _1817_ (.A1(\MOS6502.ADD[7] ),
    .A2(_0534_),
    .B1(_0227_),
    .B2(\MOS6502.ABH[7] ),
    .C1(net54),
    .X(_0261_));
 sky130_fd_sc_hd__a221o_1 _1818_ (.A1(_0549_),
    .A2(_0174_),
    .B1(_0225_),
    .B2(net200),
    .C1(_0261_),
    .X(_0262_));
 sky130_fd_sc_hd__xnor2_1 _1819_ (.A(_0259_),
    .B(_0262_),
    .Y(_0263_));
 sky130_fd_sc_hd__a22o_1 _1820_ (.A1(net200),
    .A2(net60),
    .B1(_0263_),
    .B2(net64),
    .X(_0059_));
 sky130_fd_sc_hd__or3b_1 _1821_ (.A(net68),
    .B(net71),
    .C_N(net69),
    .X(_0264_));
 sky130_fd_sc_hd__o211a_1 _1822_ (.A1(_0440_),
    .A2(_0264_),
    .B1(_0458_),
    .C1(_0449_),
    .X(_0265_));
 sky130_fd_sc_hd__a21o_1 _1823_ (.A1(\MOS6502.state[5] ),
    .A2(\MOS6502.state[4] ),
    .B1(_0265_),
    .X(_0266_));
 sky130_fd_sc_hd__or3b_1 _1824_ (.A(_0453_),
    .B(net55),
    .C_N(_0266_),
    .X(_0267_));
 sky130_fd_sc_hd__or4_1 _1825_ (.A(_0466_),
    .B(_0486_),
    .C(_0827_),
    .D(_0267_),
    .X(_0268_));
 sky130_fd_sc_hd__or4_1 _1826_ (.A(_0469_),
    .B(_0481_),
    .C(_0543_),
    .D(_0723_),
    .X(_0269_));
 sky130_fd_sc_hd__or3_1 _1827_ (.A(_0531_),
    .B(_0548_),
    .C(_0269_),
    .X(_0270_));
 sky130_fd_sc_hd__or4_1 _1828_ (.A(_0522_),
    .B(_0538_),
    .C(_0268_),
    .D(_0270_),
    .X(_0271_));
 sky130_fd_sc_hd__or4_1 _1829_ (.A(_0508_),
    .B(_0818_),
    .C(_0173_),
    .D(_0271_),
    .X(_0272_));
 sky130_fd_sc_hd__or4_1 _1830_ (.A(_0429_),
    .B(_0480_),
    .C(_0760_),
    .D(_0835_),
    .X(_0273_));
 sky130_fd_sc_hd__and2b_4 _1831_ (.A_N(_0273_),
    .B(_0272_),
    .X(_0274_));
 sky130_fd_sc_hd__mux2_1 _1832_ (.A0(net314),
    .A1(net18),
    .S(_0274_),
    .X(_0275_));
 sky130_fd_sc_hd__and2_1 _1833_ (.A(net73),
    .B(net315),
    .X(_0060_));
 sky130_fd_sc_hd__mux2_1 _1834_ (.A0(net311),
    .A1(net19),
    .S(_0274_),
    .X(_0276_));
 sky130_fd_sc_hd__and2_1 _1835_ (.A(net73),
    .B(_0276_),
    .X(_0061_));
 sky130_fd_sc_hd__mux2_1 _1836_ (.A0(net302),
    .A1(net20),
    .S(_0274_),
    .X(_0277_));
 sky130_fd_sc_hd__and2_1 _1837_ (.A(net73),
    .B(net303),
    .X(_0062_));
 sky130_fd_sc_hd__mux2_1 _1838_ (.A0(net293),
    .A1(net21),
    .S(_0274_),
    .X(_0278_));
 sky130_fd_sc_hd__and2_1 _1839_ (.A(net73),
    .B(net294),
    .X(_0063_));
 sky130_fd_sc_hd__mux2_1 _1840_ (.A0(net291),
    .A1(net22),
    .S(_0274_),
    .X(_0279_));
 sky130_fd_sc_hd__and2_1 _1841_ (.A(net73),
    .B(net292),
    .X(_0064_));
 sky130_fd_sc_hd__mux2_1 _1842_ (.A0(net295),
    .A1(net23),
    .S(_0274_),
    .X(_0280_));
 sky130_fd_sc_hd__and2_1 _1843_ (.A(net73),
    .B(_0280_),
    .X(_0065_));
 sky130_fd_sc_hd__mux2_1 _1844_ (.A0(net290),
    .A1(net24),
    .S(_0274_),
    .X(_0281_));
 sky130_fd_sc_hd__and2_1 _1845_ (.A(net73),
    .B(_0281_),
    .X(_0066_));
 sky130_fd_sc_hd__mux2_1 _1846_ (.A0(net288),
    .A1(net25),
    .S(_0274_),
    .X(_0282_));
 sky130_fd_sc_hd__and2_1 _1847_ (.A(net73),
    .B(net289),
    .X(_0067_));
 sky130_fd_sc_hd__mux2_1 _1848_ (.A0(net260),
    .A1(net40),
    .S(_0274_),
    .X(_0283_));
 sky130_fd_sc_hd__and2_1 _1849_ (.A(net73),
    .B(_0283_),
    .X(_0068_));
 sky130_fd_sc_hd__mux2_1 _1850_ (.A0(net285),
    .A1(net41),
    .S(_0274_),
    .X(_0284_));
 sky130_fd_sc_hd__and2_1 _1851_ (.A(net73),
    .B(_0284_),
    .X(_0069_));
 sky130_fd_sc_hd__mux2_1 _1852_ (.A0(net274),
    .A1(net42),
    .S(_0274_),
    .X(_0285_));
 sky130_fd_sc_hd__and2_1 _1853_ (.A(net73),
    .B(_0285_),
    .X(_0070_));
 sky130_fd_sc_hd__mux2_1 _1854_ (.A0(net270),
    .A1(net43),
    .S(_0274_),
    .X(_0286_));
 sky130_fd_sc_hd__and2_1 _1855_ (.A(net73),
    .B(net271),
    .X(_0071_));
 sky130_fd_sc_hd__mux2_1 _1856_ (.A0(net266),
    .A1(net44),
    .S(_0274_),
    .X(_0287_));
 sky130_fd_sc_hd__and2_1 _1857_ (.A(net73),
    .B(_0287_),
    .X(_0072_));
 sky130_fd_sc_hd__mux2_1 _1858_ (.A0(net267),
    .A1(net45),
    .S(_0274_),
    .X(_0288_));
 sky130_fd_sc_hd__and2_1 _1859_ (.A(net73),
    .B(_0288_),
    .X(_0073_));
 sky130_fd_sc_hd__mux2_1 _1860_ (.A0(net262),
    .A1(net46),
    .S(_0274_),
    .X(_0289_));
 sky130_fd_sc_hd__and2_1 _1861_ (.A(net73),
    .B(net263),
    .X(_0074_));
 sky130_fd_sc_hd__mux2_1 _1862_ (.A0(net279),
    .A1(net17),
    .S(_0274_),
    .X(_0290_));
 sky130_fd_sc_hd__and2_1 _1863_ (.A(net73),
    .B(_0290_),
    .X(_0075_));
 sky130_fd_sc_hd__and2_1 _1864_ (.A(net74),
    .B(_0599_),
    .X(_0076_));
 sky130_fd_sc_hd__and2_1 _1865_ (.A(net74),
    .B(net309),
    .X(_0077_));
 sky130_fd_sc_hd__and2_1 _1866_ (.A(net75),
    .B(_0585_),
    .X(_0078_));
 sky130_fd_sc_hd__and2_1 _1867_ (.A(net75),
    .B(net313),
    .X(_0079_));
 sky130_fd_sc_hd__and2_1 _1868_ (.A(net75),
    .B(_0570_),
    .X(_0080_));
 sky130_fd_sc_hd__and2_1 _1869_ (.A(net76),
    .B(net307),
    .X(_0081_));
 sky130_fd_sc_hd__and2_1 _1870_ (.A(net76),
    .B(net301),
    .X(_0082_));
 sky130_fd_sc_hd__and2_1 _1871_ (.A(net76),
    .B(_0549_),
    .X(_0083_));
 sky130_fd_sc_hd__a221o_1 _1872_ (.A1(_0436_),
    .A2(_0476_),
    .B1(_0543_),
    .B2(net240),
    .C1(_0507_),
    .X(_0291_));
 sky130_fd_sc_hd__or4b_1 _1873_ (.A(net250),
    .B(net269),
    .C(net238),
    .D_N(\MOS6502.state[3] ),
    .X(_0292_));
 sky130_fd_sc_hd__or3_1 _1874_ (.A(net257),
    .B(net240),
    .C(net198),
    .X(_0293_));
 sky130_fd_sc_hd__o21a_1 _1875_ (.A1(_0292_),
    .A2(_0293_),
    .B1(_0291_),
    .X(_0294_));
 sky130_fd_sc_hd__mux2_1 _1876_ (.A0(_0430_),
    .A1(net259),
    .S(net250),
    .X(_0295_));
 sky130_fd_sc_hd__mux2_1 _1877_ (.A0(_0295_),
    .A1(net275),
    .S(_0293_),
    .X(_0296_));
 sky130_fd_sc_hd__mux2_1 _1878_ (.A0(_0296_),
    .A1(_0599_),
    .S(_0507_),
    .X(_0297_));
 sky130_fd_sc_hd__mux2_1 _1879_ (.A0(net320),
    .A1(_0297_),
    .S(_0294_),
    .X(_0298_));
 sky130_fd_sc_hd__and2_1 _1880_ (.A(net77),
    .B(net321),
    .X(_0084_));
 sky130_fd_sc_hd__or2_2 _1881_ (.A(_0476_),
    .B(_0507_),
    .X(_0299_));
 sky130_fd_sc_hd__nand2_1 _1882_ (.A(_0490_),
    .B(_0495_),
    .Y(_0300_));
 sky130_fd_sc_hd__a2111o_1 _1883_ (.A1(net204),
    .A2(_0300_),
    .B1(_0477_),
    .C1(net250),
    .D1(net257),
    .X(_0301_));
 sky130_fd_sc_hd__o22ai_2 _1884_ (.A1(_0543_),
    .A2(_0299_),
    .B1(_0301_),
    .B2(\MOS6502.bit_ins ),
    .Y(_0302_));
 sky130_fd_sc_hd__and3b_1 _1885_ (.A_N(_0507_),
    .B(\MOS6502.ADD[1] ),
    .C(\MOS6502.plp ),
    .X(_0303_));
 sky130_fd_sc_hd__a21oi_1 _1886_ (.A1(_0507_),
    .A2(_0591_),
    .B1(_0303_),
    .Y(_0304_));
 sky130_fd_sc_hd__o21a_1 _1887_ (.A1(\MOS6502.plp ),
    .A2(_0507_),
    .B1(_0544_),
    .X(_0305_));
 sky130_fd_sc_hd__or4_1 _1888_ (.A(\MOS6502.ADD[2] ),
    .B(\MOS6502.ADD[1] ),
    .C(\MOS6502.ADD[0] ),
    .D(\MOS6502.ADD[7] ),
    .X(_0306_));
 sky130_fd_sc_hd__or4_1 _1889_ (.A(\MOS6502.ADD[5] ),
    .B(\MOS6502.ADD[6] ),
    .C(\MOS6502.ADD[4] ),
    .D(\MOS6502.ADD[3] ),
    .X(_0307_));
 sky130_fd_sc_hd__o32a_1 _1890_ (.A1(_0305_),
    .A2(_0306_),
    .A3(_0307_),
    .B1(_0304_),
    .B2(_0543_),
    .X(_0308_));
 sky130_fd_sc_hd__o21ai_1 _1891_ (.A1(_0302_),
    .A2(_0308_),
    .B1(net14),
    .Y(_0309_));
 sky130_fd_sc_hd__a21o_1 _1892_ (.A1(net231),
    .A2(_0302_),
    .B1(_0309_),
    .X(_0085_));
 sky130_fd_sc_hd__a21oi_1 _1893_ (.A1(net241),
    .A2(_0630_),
    .B1(_0299_),
    .Y(_0310_));
 sky130_fd_sc_hd__a21bo_1 _1894_ (.A1(_0544_),
    .A2(_0310_),
    .B1_N(_0301_),
    .X(_0311_));
 sky130_fd_sc_hd__nor2_1 _1895_ (.A(net55),
    .B(_0543_),
    .Y(_0312_));
 sky130_fd_sc_hd__mux2_1 _1896_ (.A0(net244),
    .A1(_0549_),
    .S(_0312_),
    .X(_0313_));
 sky130_fd_sc_hd__mux2_1 _1897_ (.A0(_0313_),
    .A1(net318),
    .S(_0311_),
    .X(_0314_));
 sky130_fd_sc_hd__and2_1 _1898_ (.A(net14),
    .B(net319),
    .X(_0086_));
 sky130_fd_sc_hd__o32a_1 _1899_ (.A1(_0485_),
    .A2(_0540_),
    .A3(_0299_),
    .B1(_0474_),
    .B2(net250),
    .X(_0315_));
 sky130_fd_sc_hd__o31a_1 _1900_ (.A1(net235),
    .A2(\MOS6502.sei ),
    .A3(_0541_),
    .B1(_0315_),
    .X(_0316_));
 sky130_fd_sc_hd__mux2_1 _1901_ (.A0(_0432_),
    .A1(\MOS6502.ADD[2] ),
    .S(_0541_),
    .X(_0317_));
 sky130_fd_sc_hd__mux2_1 _1902_ (.A0(_0317_),
    .A1(_0585_),
    .S(_0507_),
    .X(_0318_));
 sky130_fd_sc_hd__or3b_1 _1903_ (.A(_0318_),
    .B(_0485_),
    .C_N(_0316_),
    .X(_0319_));
 sky130_fd_sc_hd__o211a_1 _1904_ (.A1(net251),
    .A2(_0316_),
    .B1(_0319_),
    .C1(net77),
    .X(_0087_));
 sky130_fd_sc_hd__o41a_1 _1905_ (.A1(net250),
    .A2(net297),
    .A3(net272),
    .A4(_0477_),
    .B1(_0299_),
    .X(_0320_));
 sky130_fd_sc_hd__mux2_1 _1906_ (.A0(_0431_),
    .A1(net278),
    .S(net250),
    .X(_0321_));
 sky130_fd_sc_hd__mux2_1 _1907_ (.A0(_0321_),
    .A1(net313),
    .S(_0507_),
    .X(_0322_));
 sky130_fd_sc_hd__mux2_1 _1908_ (.A0(net298),
    .A1(_0322_),
    .S(_0320_),
    .X(_0323_));
 sky130_fd_sc_hd__and2_1 _1909_ (.A(net77),
    .B(_0323_),
    .X(_0088_));
 sky130_fd_sc_hd__xnor2_1 _1910_ (.A(net169),
    .B(net175),
    .Y(_0324_));
 sky130_fd_sc_hd__nand2_1 _1911_ (.A(_0907_),
    .B(_0324_),
    .Y(_0325_));
 sky130_fd_sc_hd__nor2_1 _1912_ (.A(net250),
    .B(net228),
    .Y(_0326_));
 sky130_fd_sc_hd__or2_1 _1913_ (.A(_0907_),
    .B(_0324_),
    .X(_0327_));
 sky130_fd_sc_hd__a32o_1 _1914_ (.A1(_0325_),
    .A2(_0326_),
    .A3(_0327_),
    .B1(net277),
    .B2(net250),
    .X(_0328_));
 sky130_fd_sc_hd__a31o_1 _1915_ (.A1(_0434_),
    .A2(net55),
    .A3(_0326_),
    .B1(_0310_),
    .X(_0329_));
 sky130_fd_sc_hd__mux2_1 _1916_ (.A0(net301),
    .A1(_0328_),
    .S(net55),
    .X(_0330_));
 sky130_fd_sc_hd__mux2_1 _1917_ (.A0(_0330_),
    .A1(net316),
    .S(_0329_),
    .X(_0331_));
 sky130_fd_sc_hd__and2_1 _1918_ (.A(net14),
    .B(net317),
    .X(_0089_));
 sky130_fd_sc_hd__and2_1 _1919_ (.A(net79),
    .B(_0835_),
    .X(_0332_));
 sky130_fd_sc_hd__nand2_4 _1920_ (.A(net79),
    .B(_0835_),
    .Y(_0333_));
 sky130_fd_sc_hd__nor2_2 _1921_ (.A(_0429_),
    .B(_0477_),
    .Y(_0334_));
 sky130_fd_sc_hd__nand2_1 _1922_ (.A(net78),
    .B(net55),
    .Y(_0335_));
 sky130_fd_sc_hd__nand2_1 _1923_ (.A(net236),
    .B(net49),
    .Y(_0336_));
 sky130_fd_sc_hd__a21oi_1 _1924_ (.A1(_0333_),
    .A2(_0336_),
    .B1(net72),
    .Y(_0090_));
 sky130_fd_sc_hd__or2_1 _1925_ (.A(\MOS6502.IRHOLD[0] ),
    .B(_0332_),
    .X(_0337_));
 sky130_fd_sc_hd__o211a_1 _1926_ (.A1(net178),
    .A2(_0333_),
    .B1(_0337_),
    .C1(net76),
    .X(_0091_));
 sky130_fd_sc_hd__a31o_1 _1927_ (.A1(net78),
    .A2(\MOS6502.DI[1] ),
    .A3(_0835_),
    .B1(net72),
    .X(_0338_));
 sky130_fd_sc_hd__a21o_1 _1928_ (.A1(net87),
    .A2(_0333_),
    .B1(_0338_),
    .X(_0092_));
 sky130_fd_sc_hd__or2_1 _1929_ (.A(\MOS6502.IRHOLD[2] ),
    .B(_0332_),
    .X(_0339_));
 sky130_fd_sc_hd__o211a_1 _1930_ (.A1(net186),
    .A2(_0333_),
    .B1(_0339_),
    .C1(net76),
    .X(_0093_));
 sky130_fd_sc_hd__a31o_1 _1931_ (.A1(net79),
    .A2(\MOS6502.DI[3] ),
    .A3(_0835_),
    .B1(net72),
    .X(_0340_));
 sky130_fd_sc_hd__a21o_1 _1932_ (.A1(net85),
    .A2(_0333_),
    .B1(_0340_),
    .X(_0094_));
 sky130_fd_sc_hd__or2_1 _1933_ (.A(\MOS6502.IRHOLD[4] ),
    .B(_0332_),
    .X(_0341_));
 sky130_fd_sc_hd__o211a_1 _1934_ (.A1(net180),
    .A2(_0333_),
    .B1(_0341_),
    .C1(net76),
    .X(_0095_));
 sky130_fd_sc_hd__a31o_1 _1935_ (.A1(net79),
    .A2(\MOS6502.DI[5] ),
    .A3(_0835_),
    .B1(net72),
    .X(_0342_));
 sky130_fd_sc_hd__a21o_1 _1936_ (.A1(net111),
    .A2(_0333_),
    .B1(_0342_),
    .X(_0096_));
 sky130_fd_sc_hd__a31o_1 _1937_ (.A1(net79),
    .A2(\MOS6502.DI[6] ),
    .A3(_0835_),
    .B1(_0441_),
    .X(_0343_));
 sky130_fd_sc_hd__a21o_1 _1938_ (.A1(net137),
    .A2(_0333_),
    .B1(_0343_),
    .X(_0097_));
 sky130_fd_sc_hd__a31o_1 _1939_ (.A1(net78),
    .A2(\MOS6502.DI[7] ),
    .A3(_0835_),
    .B1(net72),
    .X(_0344_));
 sky130_fd_sc_hd__a21o_1 _1940_ (.A1(net91),
    .A2(_0333_),
    .B1(_0344_),
    .X(_0098_));
 sky130_fd_sc_hd__and2_1 _1941_ (.A(net77),
    .B(net12),
    .X(_0099_));
 sky130_fd_sc_hd__a21o_1 _1942_ (.A1(net177),
    .A2(_0477_),
    .B1(net72),
    .X(_0100_));
 sky130_fd_sc_hd__nor2_2 _1943_ (.A(_0655_),
    .B(_0657_),
    .Y(_0345_));
 sky130_fd_sc_hd__or2_1 _1944_ (.A(_0655_),
    .B(_0657_),
    .X(_0346_));
 sky130_fd_sc_hd__nand2_2 _1945_ (.A(_0653_),
    .B(_0657_),
    .Y(_0347_));
 sky130_fd_sc_hd__or2_1 _1946_ (.A(_0639_),
    .B(_0691_),
    .X(_0348_));
 sky130_fd_sc_hd__or2_1 _1947_ (.A(_0670_),
    .B(_0348_),
    .X(_0349_));
 sky130_fd_sc_hd__nor2_1 _1948_ (.A(_0347_),
    .B(_0349_),
    .Y(_0350_));
 sky130_fd_sc_hd__a31o_1 _1949_ (.A1(_0651_),
    .A2(_0666_),
    .A3(_0345_),
    .B1(_0350_),
    .X(_0351_));
 sky130_fd_sc_hd__nor2_2 _1950_ (.A(_0647_),
    .B(_0668_),
    .Y(_0352_));
 sky130_fd_sc_hd__inv_2 _1951_ (.A(_0352_),
    .Y(_0353_));
 sky130_fd_sc_hd__o2111a_1 _1952_ (.A1(_0637_),
    .A2(_0669_),
    .B1(_0345_),
    .C1(_0643_),
    .D1(_0650_),
    .X(_0354_));
 sky130_fd_sc_hd__nor2_1 _1953_ (.A(_0650_),
    .B(_0655_),
    .Y(_0355_));
 sky130_fd_sc_hd__nor2_1 _1954_ (.A(_0675_),
    .B(_0355_),
    .Y(_0356_));
 sky130_fd_sc_hd__or4_1 _1955_ (.A(net48),
    .B(_0352_),
    .C(_0354_),
    .D(_0356_),
    .X(_0357_));
 sky130_fd_sc_hd__nand2_1 _1956_ (.A(_0648_),
    .B(_0650_),
    .Y(_0358_));
 sky130_fd_sc_hd__a2bb2o_1 _1957_ (.A1_N(_0346_),
    .A2_N(_0358_),
    .B1(_0655_),
    .B2(_0669_),
    .X(_0359_));
 sky130_fd_sc_hd__a31o_1 _1958_ (.A1(_0640_),
    .A2(_0690_),
    .A3(_0359_),
    .B1(_0357_),
    .X(_0360_));
 sky130_fd_sc_hd__o221a_1 _1959_ (.A1(net204),
    .A2(net50),
    .B1(_0351_),
    .B2(_0360_),
    .C1(net74),
    .X(_0101_));
 sky130_fd_sc_hd__nand2_1 _1960_ (.A(_0651_),
    .B(_0668_),
    .Y(_0361_));
 sky130_fd_sc_hd__o32a_1 _1961_ (.A1(_0346_),
    .A2(_0348_),
    .A3(_0361_),
    .B1(_0677_),
    .B2(_0635_),
    .X(_0362_));
 sky130_fd_sc_hd__a211o_1 _1962_ (.A1(_0638_),
    .A2(_0648_),
    .B1(_0651_),
    .C1(_0646_),
    .X(_0363_));
 sky130_fd_sc_hd__o2bb2a_1 _1963_ (.A1_N(_0352_),
    .A2_N(_0355_),
    .B1(_0363_),
    .B2(_0346_),
    .X(_0364_));
 sky130_fd_sc_hd__nand2_1 _1964_ (.A(_0362_),
    .B(_0364_),
    .Y(_0365_));
 sky130_fd_sc_hd__or2_1 _1965_ (.A(net208),
    .B(net50),
    .X(_0366_));
 sky130_fd_sc_hd__o211a_1 _1966_ (.A1(net49),
    .A2(_0365_),
    .B1(_0366_),
    .C1(net74),
    .X(_0102_));
 sky130_fd_sc_hd__a21oi_1 _1967_ (.A1(_0349_),
    .A2(_0353_),
    .B1(_0347_),
    .Y(_0367_));
 sky130_fd_sc_hd__a311o_1 _1968_ (.A1(_0650_),
    .A2(_0690_),
    .A3(_0345_),
    .B1(_0365_),
    .C1(_0367_),
    .X(_0368_));
 sky130_fd_sc_hd__a21o_1 _1969_ (.A1(net286),
    .A2(net49),
    .B1(net72),
    .X(_0369_));
 sky130_fd_sc_hd__a31o_1 _1970_ (.A1(net50),
    .A2(_0362_),
    .A3(_0368_),
    .B1(_0369_),
    .X(_0103_));
 sky130_fd_sc_hd__mux2_1 _1971_ (.A0(_0678_),
    .A1(_0648_),
    .S(_0657_),
    .X(_0370_));
 sky130_fd_sc_hd__or4_1 _1972_ (.A(_0646_),
    .B(_0650_),
    .C(_0655_),
    .D(_0370_),
    .X(_0371_));
 sky130_fd_sc_hd__or3_1 _1973_ (.A(_0346_),
    .B(_0348_),
    .C(_0358_),
    .X(_0372_));
 sky130_fd_sc_hd__a21oi_1 _1974_ (.A1(_0371_),
    .A2(_0372_),
    .B1(net48),
    .Y(_0373_));
 sky130_fd_sc_hd__a211o_1 _1975_ (.A1(net145),
    .A2(net49),
    .B1(_0373_),
    .C1(net72),
    .X(_0104_));
 sky130_fd_sc_hd__a41o_1 _1976_ (.A1(_0637_),
    .A2(_0643_),
    .A3(_0651_),
    .A4(_0345_),
    .B1(net49),
    .X(_0374_));
 sky130_fd_sc_hd__o31a_1 _1977_ (.A1(_0646_),
    .A2(_0652_),
    .A3(_0347_),
    .B1(_0371_),
    .X(_0375_));
 sky130_fd_sc_hd__or3b_1 _1978_ (.A(_0351_),
    .B(_0374_),
    .C_N(_0375_),
    .X(_0376_));
 sky130_fd_sc_hd__o211a_1 _1979_ (.A1(net163),
    .A2(net50),
    .B1(_0376_),
    .C1(net74),
    .X(_0105_));
 sky130_fd_sc_hd__and4_1 _1980_ (.A(_0637_),
    .B(_0648_),
    .C(_0690_),
    .D(_0345_),
    .X(_0377_));
 sky130_fd_sc_hd__o211a_1 _1981_ (.A1(_0634_),
    .A2(_0668_),
    .B1(_0674_),
    .C1(_0638_),
    .X(_0378_));
 sky130_fd_sc_hd__or2_1 _1982_ (.A(net245),
    .B(net50),
    .X(_0379_));
 sky130_fd_sc_hd__o311a_1 _1983_ (.A1(net49),
    .A2(_0377_),
    .A3(_0378_),
    .B1(_0379_),
    .C1(net76),
    .X(_0106_));
 sky130_fd_sc_hd__and3_1 _1984_ (.A(_0651_),
    .B(_0674_),
    .C(_0345_),
    .X(_0380_));
 sky130_fd_sc_hd__o221a_1 _1985_ (.A1(net215),
    .A2(net50),
    .B1(_0374_),
    .B2(_0380_),
    .C1(net74),
    .X(_0107_));
 sky130_fd_sc_hd__a31o_1 _1986_ (.A1(_0637_),
    .A2(_0690_),
    .A3(_0346_),
    .B1(net48),
    .X(_0381_));
 sky130_fd_sc_hd__o211a_1 _1987_ (.A1(net233),
    .A2(_0334_),
    .B1(_0381_),
    .C1(net77),
    .X(_0108_));
 sky130_fd_sc_hd__a21o_1 _1988_ (.A1(_0650_),
    .A2(_0345_),
    .B1(net48),
    .X(_0382_));
 sky130_fd_sc_hd__o211a_1 _1989_ (.A1(net237),
    .A2(_0334_),
    .B1(_0382_),
    .C1(net75),
    .X(_0109_));
 sky130_fd_sc_hd__nor2_1 _1990_ (.A(net48),
    .B(_0347_),
    .Y(_0383_));
 sky130_fd_sc_hd__a31o_1 _1991_ (.A1(_0637_),
    .A2(_0650_),
    .A3(_0690_),
    .B1(_0352_),
    .X(_0384_));
 sky130_fd_sc_hd__a22o_1 _1992_ (.A1(net229),
    .A2(net48),
    .B1(_0383_),
    .B2(_0384_),
    .X(_0385_));
 sky130_fd_sc_hd__and2_1 _1993_ (.A(net75),
    .B(net230),
    .X(_0110_));
 sky130_fd_sc_hd__nand2_1 _1994_ (.A(net78),
    .B(_0826_),
    .Y(_0386_));
 sky130_fd_sc_hd__nand2_1 _1995_ (.A(_0650_),
    .B(_0657_),
    .Y(_0387_));
 sky130_fd_sc_hd__nor3_1 _1996_ (.A(_0675_),
    .B(_0386_),
    .C(_0387_),
    .Y(_0388_));
 sky130_fd_sc_hd__and2_1 _1997_ (.A(net198),
    .B(_0386_),
    .X(_0389_));
 sky130_fd_sc_hd__o21a_1 _1998_ (.A1(_0388_),
    .A2(_0389_),
    .B1(net74),
    .X(_0111_));
 sky130_fd_sc_hd__a32o_1 _1999_ (.A1(net298),
    .A2(_0655_),
    .A3(_0388_),
    .B1(_0386_),
    .B2(\MOS6502.adc_bcd ),
    .X(_0390_));
 sky130_fd_sc_hd__and2_1 _2000_ (.A(net74),
    .B(net299),
    .X(_0112_));
 sky130_fd_sc_hd__and4_1 _2001_ (.A(_0655_),
    .B(_0679_),
    .C(_0690_),
    .D(net50),
    .X(_0391_));
 sky130_fd_sc_hd__a21oi_1 _2002_ (.A1(net240),
    .A2(net48),
    .B1(_0391_),
    .Y(_0392_));
 sky130_fd_sc_hd__nor2_1 _2003_ (.A(net72),
    .B(_0392_),
    .Y(_0113_));
 sky130_fd_sc_hd__o32a_1 _2004_ (.A1(_0640_),
    .A2(_0646_),
    .A3(_0668_),
    .B1(_0675_),
    .B2(_0650_),
    .X(_0393_));
 sky130_fd_sc_hd__nor2_1 _2005_ (.A(_0347_),
    .B(_0393_),
    .Y(_0394_));
 sky130_fd_sc_hd__or2_1 _2006_ (.A(net257),
    .B(net50),
    .X(_0395_));
 sky130_fd_sc_hd__o211a_1 _2007_ (.A1(net49),
    .A2(_0394_),
    .B1(_0395_),
    .C1(net74),
    .X(_0114_));
 sky130_fd_sc_hd__nor2_1 _2008_ (.A(_0659_),
    .B(_0691_),
    .Y(_0396_));
 sky130_fd_sc_hd__or2_1 _2009_ (.A(net253),
    .B(net50),
    .X(_0397_));
 sky130_fd_sc_hd__o211a_1 _2010_ (.A1(net49),
    .A2(_0396_),
    .B1(_0397_),
    .C1(net74),
    .X(_0115_));
 sky130_fd_sc_hd__a22o_1 _2011_ (.A1(net287),
    .A2(net48),
    .B1(_0391_),
    .B2(_0650_),
    .X(_0398_));
 sky130_fd_sc_hd__and2_1 _2012_ (.A(net75),
    .B(_0398_),
    .X(_0116_));
 sky130_fd_sc_hd__o31a_1 _2013_ (.A1(_0650_),
    .A2(_0654_),
    .A3(_0675_),
    .B1(net50),
    .X(_0399_));
 sky130_fd_sc_hd__a211o_1 _2014_ (.A1(net227),
    .A2(net49),
    .B1(_0399_),
    .C1(net72),
    .X(_0117_));
 sky130_fd_sc_hd__nor4_1 _2015_ (.A(_0638_),
    .B(_0646_),
    .C(_0651_),
    .D(_0687_),
    .Y(_0400_));
 sky130_fd_sc_hd__o311a_1 _2016_ (.A1(_0638_),
    .A2(_0650_),
    .A3(_0691_),
    .B1(_0349_),
    .C1(_0675_),
    .X(_0401_));
 sky130_fd_sc_hd__a31o_1 _2017_ (.A1(_0655_),
    .A2(_0674_),
    .A3(_0387_),
    .B1(_0396_),
    .X(_0402_));
 sky130_fd_sc_hd__a311o_1 _2018_ (.A1(_0651_),
    .A2(_0345_),
    .A3(_0352_),
    .B1(_0400_),
    .C1(_0402_),
    .X(_0403_));
 sky130_fd_sc_hd__nor2_1 _2019_ (.A(_0394_),
    .B(_0403_),
    .Y(_0404_));
 sky130_fd_sc_hd__o21a_1 _2020_ (.A1(_0347_),
    .A2(_0401_),
    .B1(_0404_),
    .X(_0405_));
 sky130_fd_sc_hd__o21a_1 _2021_ (.A1(_0686_),
    .A2(_0691_),
    .B1(_0405_),
    .X(_0406_));
 sky130_fd_sc_hd__o31a_1 _2022_ (.A1(_0686_),
    .A2(_0690_),
    .A3(_0405_),
    .B1(_0334_),
    .X(_0407_));
 sky130_fd_sc_hd__a211o_1 _2023_ (.A1(net167),
    .A2(net49),
    .B1(_0407_),
    .C1(net72),
    .X(_0118_));
 sky130_fd_sc_hd__nand2_1 _2024_ (.A(net50),
    .B(_0405_),
    .Y(_0408_));
 sky130_fd_sc_hd__o211a_1 _2025_ (.A1(net243),
    .A2(net50),
    .B1(_0408_),
    .C1(net74),
    .X(_0119_));
 sky130_fd_sc_hd__o21ai_1 _2026_ (.A1(_0653_),
    .A2(_0406_),
    .B1(net50),
    .Y(_0409_));
 sky130_fd_sc_hd__o211a_1 _2027_ (.A1(net206),
    .A2(net50),
    .B1(_0409_),
    .C1(net74),
    .X(_0120_));
 sky130_fd_sc_hd__or2_1 _2028_ (.A(net241),
    .B(net50),
    .X(_0410_));
 sky130_fd_sc_hd__o211a_1 _2029_ (.A1(net49),
    .A2(_0400_),
    .B1(_0410_),
    .C1(net74),
    .X(_0121_));
 sky130_fd_sc_hd__nor2_1 _2030_ (.A(_0647_),
    .B(_0358_),
    .Y(_0411_));
 sky130_fd_sc_hd__and2_1 _2031_ (.A(_0334_),
    .B(_0411_),
    .X(_0412_));
 sky130_fd_sc_hd__a22o_1 _2032_ (.A1(net228),
    .A2(net49),
    .B1(_0345_),
    .B2(_0412_),
    .X(_0413_));
 sky130_fd_sc_hd__and2_1 _2033_ (.A(net75),
    .B(_0413_),
    .X(_0122_));
 sky130_fd_sc_hd__a22o_1 _2034_ (.A1(net268),
    .A2(net48),
    .B1(_0412_),
    .B2(_0658_),
    .X(_0414_));
 sky130_fd_sc_hd__and2_1 _2035_ (.A(net77),
    .B(_0414_),
    .X(_0123_));
 sky130_fd_sc_hd__nor2_1 _2036_ (.A(_0647_),
    .B(_0361_),
    .Y(_0415_));
 sky130_fd_sc_hd__a21o_1 _2037_ (.A1(_0658_),
    .A2(_0415_),
    .B1(net48),
    .X(_0416_));
 sky130_fd_sc_hd__o211a_1 _2038_ (.A1(net235),
    .A2(net50),
    .B1(_0416_),
    .C1(net77),
    .X(_0124_));
 sky130_fd_sc_hd__a22o_1 _2039_ (.A1(net272),
    .A2(net48),
    .B1(_0383_),
    .B2(_0411_),
    .X(_0417_));
 sky130_fd_sc_hd__and2_1 _2040_ (.A(net75),
    .B(net273),
    .X(_0125_));
 sky130_fd_sc_hd__a22o_1 _2041_ (.A1(net297),
    .A2(net48),
    .B1(_0383_),
    .B2(_0415_),
    .X(_0418_));
 sky130_fd_sc_hd__and2_1 _2042_ (.A(net75),
    .B(_0418_),
    .X(_0126_));
 sky130_fd_sc_hd__nor2_1 _2043_ (.A(_0686_),
    .B(net48),
    .Y(_0419_));
 sky130_fd_sc_hd__a22o_1 _2044_ (.A1(net238),
    .A2(net48),
    .B1(_0411_),
    .B2(_0419_),
    .X(_0420_));
 sky130_fd_sc_hd__and2_1 _2045_ (.A(net77),
    .B(net239),
    .X(_0127_));
 sky130_fd_sc_hd__a22o_1 _2046_ (.A1(net269),
    .A2(net48),
    .B1(_0415_),
    .B2(_0419_),
    .X(_0421_));
 sky130_fd_sc_hd__and2_1 _2047_ (.A(net77),
    .B(_0421_),
    .X(_0128_));
 sky130_fd_sc_hd__a32o_1 _2048_ (.A1(_0651_),
    .A2(_0352_),
    .A3(_0419_),
    .B1(net48),
    .B2(net280),
    .X(_0422_));
 sky130_fd_sc_hd__and2_1 _2049_ (.A(net75),
    .B(net281),
    .X(_0129_));
 sky130_fd_sc_hd__o21ai_1 _2050_ (.A1(_0647_),
    .A2(_0687_),
    .B1(_0334_),
    .Y(_0423_));
 sky130_fd_sc_hd__o211a_1 _2051_ (.A1(net250),
    .A2(_0334_),
    .B1(_0423_),
    .C1(net77),
    .X(_0130_));
 sky130_fd_sc_hd__a22o_1 _2052_ (.A1(net171),
    .A2(net59),
    .B1(_0650_),
    .B2(net63),
    .X(_0131_));
 sky130_fd_sc_hd__a22o_1 _2053_ (.A1(net157),
    .A2(net59),
    .B1(_0657_),
    .B2(net64),
    .X(_0132_));
 sky130_fd_sc_hd__a22o_1 _2054_ (.A1(net165),
    .A2(net59),
    .B1(_0654_),
    .B2(_0620_),
    .X(_0133_));
 sky130_fd_sc_hd__or3b_1 _2055_ (.A(\MOS6502.NMI_edge ),
    .B(net247),
    .C_N(net12),
    .X(_0424_));
 sky130_fd_sc_hd__o21ai_1 _2056_ (.A1(_0428_),
    .A2(_0485_),
    .B1(net248),
    .Y(_0425_));
 sky130_fd_sc_hd__and2_1 _2057_ (.A(net77),
    .B(net249),
    .X(_0134_));
 sky130_fd_sc_hd__a31o_4 _2058_ (.A1(_0490_),
    .A2(_0496_),
    .A3(_0867_),
    .B1(net72),
    .X(_0426_));
 sky130_fd_sc_hd__mux2_1 _2059_ (.A0(net119),
    .A1(_0872_),
    .S(_0426_),
    .X(_0135_));
 sky130_fd_sc_hd__mux2_1 _2060_ (.A0(net97),
    .A1(_0879_),
    .S(_0426_),
    .X(_0136_));
 sky130_fd_sc_hd__mux2_1 _2061_ (.A0(net133),
    .A1(_0886_),
    .S(_0426_),
    .X(_0137_));
 sky130_fd_sc_hd__mux2_1 _2062_ (.A0(net155),
    .A1(_0891_),
    .S(_0426_),
    .X(_0138_));
 sky130_fd_sc_hd__mux2_1 _2063_ (.A0(net147),
    .A1(_0893_),
    .S(_0426_),
    .X(_0139_));
 sky130_fd_sc_hd__mux2_1 _2064_ (.A0(net107),
    .A1(_0899_),
    .S(_0426_),
    .X(_0140_));
 sky130_fd_sc_hd__mux2_1 _2065_ (.A0(net113),
    .A1(_0905_),
    .S(_0426_),
    .X(_0141_));
 sky130_fd_sc_hd__mux2_1 _2066_ (.A0(net129),
    .A1(_0911_),
    .S(_0426_),
    .X(_0142_));
 sky130_fd_sc_hd__a31o_4 _2067_ (.A1(_0491_),
    .A2(_0495_),
    .A3(_0866_),
    .B1(net72),
    .X(_0427_));
 sky130_fd_sc_hd__mux2_1 _2068_ (.A0(net121),
    .A1(_0872_),
    .S(_0427_),
    .X(_0143_));
 sky130_fd_sc_hd__mux2_1 _2069_ (.A0(net141),
    .A1(_0879_),
    .S(_0427_),
    .X(_0144_));
 sky130_fd_sc_hd__mux2_1 _2070_ (.A0(net123),
    .A1(_0886_),
    .S(_0427_),
    .X(_0145_));
 sky130_fd_sc_hd__mux2_1 _2071_ (.A0(net117),
    .A1(_0891_),
    .S(_0427_),
    .X(_0146_));
 sky130_fd_sc_hd__mux2_1 _2072_ (.A0(net95),
    .A1(_0893_),
    .S(_0427_),
    .X(_0147_));
 sky130_fd_sc_hd__mux2_1 _2073_ (.A0(net109),
    .A1(_0899_),
    .S(_0427_),
    .X(_0148_));
 sky130_fd_sc_hd__mux2_1 _2074_ (.A0(net131),
    .A1(_0905_),
    .S(_0427_),
    .X(_0149_));
 sky130_fd_sc_hd__mux2_1 _2075_ (.A0(net101),
    .A1(_0911_),
    .S(_0427_),
    .X(_0150_));
 sky130_fd_sc_hd__dfxtp_1 _2076_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(net170),
    .Q(\MOS6502.ALU.BI7 ));
 sky130_fd_sc_hd__dfxtp_1 _2077_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(net324),
    .Q(\MOS6502.state[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2078_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_0002_),
    .Q(\MOS6502.state[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2079_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_0003_),
    .Q(\MOS6502.state[2] ));
 sky130_fd_sc_hd__dfxtp_2 _2080_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_0004_),
    .Q(\MOS6502.state[3] ));
 sky130_fd_sc_hd__dfxtp_2 _2081_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_0005_),
    .Q(\MOS6502.state[4] ));
 sky130_fd_sc_hd__dfxtp_2 _2082_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_0006_),
    .Q(\MOS6502.state[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2083_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(net150),
    .Q(\MOS6502.AXYS[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2084_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(net94),
    .Q(\MOS6502.AXYS[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2085_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(net160),
    .Q(\MOS6502.AXYS[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2086_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(net128),
    .Q(\MOS6502.AXYS[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2087_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(net136),
    .Q(\MOS6502.AXYS[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _2088_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(net126),
    .Q(\MOS6502.AXYS[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _2089_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(net152),
    .Q(\MOS6502.AXYS[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _2090_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(net106),
    .Q(\MOS6502.AXYS[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _2091_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_0016_),
    .Q(\MOS6502.DI[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2092_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_0017_),
    .Q(\MOS6502.DI[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2093_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_0018_),
    .Q(\MOS6502.DI[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2094_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_0019_),
    .Q(\MOS6502.DI[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2095_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_0020_),
    .Q(\MOS6502.DI[4] ));
 sky130_fd_sc_hd__dfxtp_1 _2096_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_0021_),
    .Q(\MOS6502.DI[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2097_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_0022_),
    .Q(\MOS6502.DI[6] ));
 sky130_fd_sc_hd__dfxtp_1 _2098_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(_0023_),
    .Q(\MOS6502.DI[7] ));
 sky130_fd_sc_hd__dfxtp_1 _2099_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(net162),
    .Q(\MOS6502.AXYS[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2100_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(net140),
    .Q(\MOS6502.AXYS[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2101_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(net144),
    .Q(\MOS6502.AXYS[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2102_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(net154),
    .Q(\MOS6502.AXYS[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2103_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(net100),
    .Q(\MOS6502.AXYS[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _2104_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(net116),
    .Q(\MOS6502.AXYS[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _2105_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(net104),
    .Q(\MOS6502.AXYS[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _2106_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(net90),
    .Q(\MOS6502.AXYS[1][7] ));
 sky130_fd_sc_hd__dfxtp_2 _2107_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(net193),
    .Q(\MOS6502.backwards ));
 sky130_fd_sc_hd__dfxtp_2 _2108_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(net276),
    .Q(\MOS6502.ALU.CO ));
 sky130_fd_sc_hd__dfxtp_1 _2109_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(net174),
    .Q(\MOS6502.ALU.HC ));
 sky130_fd_sc_hd__dfxtp_2 _2110_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_0035_),
    .Q(\MOS6502.ADD[0] ));
 sky130_fd_sc_hd__dfxtp_2 _2111_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_0036_),
    .Q(\MOS6502.ADD[1] ));
 sky130_fd_sc_hd__dfxtp_4 _2112_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_0037_),
    .Q(\MOS6502.ADD[2] ));
 sky130_fd_sc_hd__dfxtp_2 _2113_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_0038_),
    .Q(\MOS6502.ADD[3] ));
 sky130_fd_sc_hd__dfxtp_2 _2114_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(net256),
    .Q(\MOS6502.ADD[4] ));
 sky130_fd_sc_hd__dfxtp_2 _2115_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(net265),
    .Q(\MOS6502.ADD[5] ));
 sky130_fd_sc_hd__dfxtp_2 _2116_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_0041_),
    .Q(\MOS6502.ADD[6] ));
 sky130_fd_sc_hd__dfxtp_2 _2117_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_0042_),
    .Q(\MOS6502.ADD[7] ));
 sky130_fd_sc_hd__dfxtp_1 _2118_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(net176),
    .Q(\MOS6502.ALU.AI7 ));
 sky130_fd_sc_hd__dfxtp_1 _2119_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(net224),
    .Q(\MOS6502.PC[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2120_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(net220),
    .Q(\MOS6502.PC[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2121_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(net218),
    .Q(\MOS6502.PC[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2122_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(net214),
    .Q(\MOS6502.PC[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2123_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(net222),
    .Q(\MOS6502.PC[4] ));
 sky130_fd_sc_hd__dfxtp_1 _2124_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(net226),
    .Q(\MOS6502.PC[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2125_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(net212),
    .Q(\MOS6502.PC[6] ));
 sky130_fd_sc_hd__dfxtp_1 _2126_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(net210),
    .Q(\MOS6502.PC[7] ));
 sky130_fd_sc_hd__dfxtp_1 _2127_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(net185),
    .Q(\MOS6502.PC[8] ));
 sky130_fd_sc_hd__dfxtp_1 _2128_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(net183),
    .Q(\MOS6502.PC[9] ));
 sky130_fd_sc_hd__dfxtp_1 _2129_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(net189),
    .Q(\MOS6502.PC[10] ));
 sky130_fd_sc_hd__dfxtp_1 _2130_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(net195),
    .Q(\MOS6502.PC[11] ));
 sky130_fd_sc_hd__dfxtp_1 _2131_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(net191),
    .Q(\MOS6502.PC[12] ));
 sky130_fd_sc_hd__dfxtp_1 _2132_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(net197),
    .Q(\MOS6502.PC[13] ));
 sky130_fd_sc_hd__dfxtp_1 _2133_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(net203),
    .Q(\MOS6502.PC[14] ));
 sky130_fd_sc_hd__dfxtp_1 _2134_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(net201),
    .Q(\MOS6502.PC[15] ));
 sky130_fd_sc_hd__dfxtp_1 _2135_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_0060_),
    .Q(\MOS6502.ABH[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2136_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_0061_),
    .Q(\MOS6502.ABH[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2137_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_0062_),
    .Q(\MOS6502.ABH[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2138_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_0063_),
    .Q(\MOS6502.ABH[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2139_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_0064_),
    .Q(\MOS6502.ABH[4] ));
 sky130_fd_sc_hd__dfxtp_1 _2140_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_0065_),
    .Q(\MOS6502.ABH[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2141_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_0066_),
    .Q(\MOS6502.ABH[6] ));
 sky130_fd_sc_hd__dfxtp_1 _2142_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_0067_),
    .Q(\MOS6502.ABH[7] ));
 sky130_fd_sc_hd__dfxtp_1 _2143_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_0068_),
    .Q(\MOS6502.ABL[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2144_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_0069_),
    .Q(\MOS6502.ABL[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2145_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_0070_),
    .Q(\MOS6502.ABL[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2146_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_0071_),
    .Q(\MOS6502.ABL[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2147_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_0072_),
    .Q(\MOS6502.ABL[4] ));
 sky130_fd_sc_hd__dfxtp_1 _2148_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_0073_),
    .Q(\MOS6502.ABL[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2149_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_0074_),
    .Q(\MOS6502.ABL[6] ));
 sky130_fd_sc_hd__dfxtp_1 _2150_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_0075_),
    .Q(\MOS6502.ABL[7] ));
 sky130_fd_sc_hd__dfxtp_1 _2151_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(net199),
    .Q(\MOS6502.adj_bcd ));
 sky130_fd_sc_hd__dfxtp_1 _2152_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_0076_),
    .Q(\MOS6502.DIHOLD[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2153_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_0077_),
    .Q(\MOS6502.DIHOLD[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2154_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_0078_),
    .Q(\MOS6502.DIHOLD[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2155_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_0079_),
    .Q(\MOS6502.DIHOLD[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2156_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(_0080_),
    .Q(\MOS6502.DIHOLD[4] ));
 sky130_fd_sc_hd__dfxtp_1 _2157_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_0081_),
    .Q(\MOS6502.DIHOLD[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2158_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(_0082_),
    .Q(\MOS6502.DIHOLD[6] ));
 sky130_fd_sc_hd__dfxtp_1 _2159_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_0083_),
    .Q(\MOS6502.DIHOLD[7] ));
 sky130_fd_sc_hd__dfxtp_4 _2160_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_0084_),
    .Q(net16));
 sky130_fd_sc_hd__dfxtp_2 _2161_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(net232),
    .Q(net27));
 sky130_fd_sc_hd__dfxtp_2 _2162_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_0086_),
    .Q(net39));
 sky130_fd_sc_hd__dfxtp_2 _2163_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(net252),
    .Q(net37));
 sky130_fd_sc_hd__dfxtp_2 _2164_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_0088_),
    .Q(net36));
 sky130_fd_sc_hd__dfxtp_2 _2165_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_0089_),
    .Q(net38));
 sky130_fd_sc_hd__dfxtp_2 _2166_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_0090_),
    .Q(\MOS6502.IRHOLD_valid ));
 sky130_fd_sc_hd__dfxtp_1 _2167_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(net179),
    .Q(\MOS6502.IRHOLD[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2168_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(net88),
    .Q(\MOS6502.IRHOLD[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2169_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(net187),
    .Q(\MOS6502.IRHOLD[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2170_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(net86),
    .Q(\MOS6502.IRHOLD[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2171_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(net181),
    .Q(\MOS6502.IRHOLD[4] ));
 sky130_fd_sc_hd__dfxtp_1 _2172_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(net112),
    .Q(\MOS6502.IRHOLD[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2173_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(net138),
    .Q(\MOS6502.IRHOLD[6] ));
 sky130_fd_sc_hd__dfxtp_1 _2174_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(net92),
    .Q(\MOS6502.IRHOLD[7] ));
 sky130_fd_sc_hd__dfxtp_1 _2175_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_0099_),
    .Q(\MOS6502.NMI_1 ));
 sky130_fd_sc_hd__dfxtp_1 _2176_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(_0100_),
    .Q(\MOS6502.res ));
 sky130_fd_sc_hd__dfxtp_1 _2177_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(net205),
    .Q(\MOS6502.load_reg ));
 sky130_fd_sc_hd__dfxtp_1 _2178_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(_0102_),
    .Q(\MOS6502.dst_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2179_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(_0103_),
    .Q(\MOS6502.dst_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2180_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(net146),
    .Q(\MOS6502.src_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2181_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(net164),
    .Q(\MOS6502.src_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2182_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(net246),
    .Q(\MOS6502.index_y ));
 sky130_fd_sc_hd__dfxtp_1 _2183_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(net216),
    .Q(\MOS6502.store ));
 sky130_fd_sc_hd__dfxtp_1 _2184_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(net234),
    .Q(\MOS6502.write_back ));
 sky130_fd_sc_hd__dfxtp_1 _2185_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_0109_),
    .Q(\MOS6502.load_only ));
 sky130_fd_sc_hd__dfxtp_1 _2186_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_0110_),
    .Q(\MOS6502.inc ));
 sky130_fd_sc_hd__dfxtp_1 _2187_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(_0111_),
    .Q(\MOS6502.adc_sbc ));
 sky130_fd_sc_hd__dfxtp_1 _2188_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(_0112_),
    .Q(\MOS6502.adc_bcd ));
 sky130_fd_sc_hd__dfxtp_1 _2189_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_0113_),
    .Q(\MOS6502.shift ));
 sky130_fd_sc_hd__dfxtp_1 _2190_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(net258),
    .Q(\MOS6502.compare ));
 sky130_fd_sc_hd__dfxtp_1 _2191_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(net254),
    .Q(\MOS6502.shift_right ));
 sky130_fd_sc_hd__dfxtp_1 _2192_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_0116_),
    .Q(\MOS6502.rotate ));
 sky130_fd_sc_hd__dfxtp_1 _2193_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_0117_),
    .Q(\MOS6502.op[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2194_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(net168),
    .Q(\MOS6502.op[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2195_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_0119_),
    .Q(\MOS6502.op[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2196_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(net207),
    .Q(\MOS6502.op[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2197_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(net242),
    .Q(\MOS6502.bit_ins ));
 sky130_fd_sc_hd__dfxtp_1 _2198_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_0122_),
    .Q(\MOS6502.clv ));
 sky130_fd_sc_hd__dfxtp_1 _2199_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_0123_),
    .Q(\MOS6502.sei ));
 sky130_fd_sc_hd__dfxtp_1 _2200_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_0124_),
    .Q(\MOS6502.cli ));
 sky130_fd_sc_hd__dfxtp_1 _2201_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_0125_),
    .Q(\MOS6502.sed ));
 sky130_fd_sc_hd__dfxtp_1 _2202_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_0126_),
    .Q(\MOS6502.cld ));
 sky130_fd_sc_hd__dfxtp_1 _2203_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_0127_),
    .Q(\MOS6502.sec ));
 sky130_fd_sc_hd__dfxtp_1 _2204_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_0128_),
    .Q(\MOS6502.clc ));
 sky130_fd_sc_hd__dfxtp_2 _2205_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_0129_),
    .Q(\MOS6502.php ));
 sky130_fd_sc_hd__dfxtp_1 _2206_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_0130_),
    .Q(\MOS6502.plp ));
 sky130_fd_sc_hd__dfxtp_1 _2207_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(net172),
    .Q(\MOS6502.cond_code[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2208_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(net158),
    .Q(\MOS6502.cond_code[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2209_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(net166),
    .Q(\MOS6502.cond_code[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2210_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_0134_),
    .Q(\MOS6502.NMI_edge ));
 sky130_fd_sc_hd__dfxtp_1 _2211_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(net120),
    .Q(\MOS6502.AXYS[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2212_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(net98),
    .Q(\MOS6502.AXYS[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2213_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(net134),
    .Q(\MOS6502.AXYS[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2214_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(net156),
    .Q(\MOS6502.AXYS[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2215_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(net148),
    .Q(\MOS6502.AXYS[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _2216_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(net108),
    .Q(\MOS6502.AXYS[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _2217_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(net114),
    .Q(\MOS6502.AXYS[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _2218_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(net130),
    .Q(\MOS6502.AXYS[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _2219_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(net122),
    .Q(\MOS6502.AXYS[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2220_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(net142),
    .Q(\MOS6502.AXYS[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2221_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(net124),
    .Q(\MOS6502.AXYS[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2222_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(net118),
    .Q(\MOS6502.AXYS[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2223_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(net96),
    .Q(\MOS6502.AXYS[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _2224_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(net110),
    .Q(\MOS6502.AXYS[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _2225_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(net132),
    .Q(\MOS6502.AXYS[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _2226_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(net102),
    .Q(\MOS6502.AXYS[3][7] ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_wb_clk_i (.A(wb_clk_i),
    .X(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_0_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_10_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_11_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_12_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_13_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_14_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_15_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_1_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_2_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_3_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_4_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_5_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_6_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_7_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_8_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_9_0_wb_clk_i));
 sky130_fd_sc_hd__buf_4 fanout48 (.A(net49),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_4 fanout49 (.A(_0335_),
    .X(net49));
 sky130_fd_sc_hd__buf_4 fanout50 (.A(_0334_),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_8 fanout52 (.A(_0632_),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_8 fanout53 (.A(_0527_),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_8 fanout54 (.A(_0509_),
    .X(net54));
 sky130_fd_sc_hd__buf_6 fanout55 (.A(_0476_),
    .X(net55));
 sky130_fd_sc_hd__buf_4 fanout56 (.A(net57),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_4 fanout57 (.A(net59),
    .X(net57));
 sky130_fd_sc_hd__buf_4 fanout58 (.A(net59),
    .X(net58));
 sky130_fd_sc_hd__buf_2 fanout59 (.A(_0628_),
    .X(net59));
 sky130_fd_sc_hd__buf_4 fanout60 (.A(_0628_),
    .X(net60));
 sky130_fd_sc_hd__buf_4 fanout61 (.A(net62),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_4 fanout62 (.A(net63),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_4 fanout63 (.A(net64),
    .X(net63));
 sky130_fd_sc_hd__buf_4 fanout64 (.A(_0620_),
    .X(net64));
 sky130_fd_sc_hd__buf_8 fanout65 (.A(_0462_),
    .X(net65));
 sky130_fd_sc_hd__buf_6 fanout66 (.A(_0448_),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_8 fanout67 (.A(_0444_),
    .X(net67));
 sky130_fd_sc_hd__buf_4 fanout68 (.A(\MOS6502.state[3] ),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_4 fanout69 (.A(\MOS6502.state[2] ),
    .X(net69));
 sky130_fd_sc_hd__buf_4 fanout70 (.A(\MOS6502.state[1] ),
    .X(net70));
 sky130_fd_sc_hd__buf_4 fanout71 (.A(\MOS6502.state[0] ),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_8 fanout72 (.A(_0441_),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_4 fanout73 (.A(net14),
    .X(net73));
 sky130_fd_sc_hd__buf_4 fanout74 (.A(net76),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_4 fanout75 (.A(net76),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_4 fanout76 (.A(net77),
    .X(net76));
 sky130_fd_sc_hd__buf_4 fanout77 (.A(net14),
    .X(net77));
 sky130_fd_sc_hd__buf_6 fanout78 (.A(net79),
    .X(net78));
 sky130_fd_sc_hd__buf_6 fanout79 (.A(net13),
    .X(net79));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\MOS6502.IRHOLD[3] ),
    .X(net85));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(_0009_),
    .X(net94));
 sky130_fd_sc_hd__buf_1 hold100 (.A(\MOS6502.PC[8] ),
    .X(net184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(_0052_),
    .X(net185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(\MOS6502.DI[2] ),
    .X(net186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(_0093_),
    .X(net187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(\MOS6502.PC[10] ),
    .X(net188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(_0054_),
    .X(net189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(\MOS6502.PC[12] ),
    .X(net190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(_0056_),
    .X(net191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(\MOS6502.DI[7] ),
    .X(net192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(_0032_),
    .X(net193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\MOS6502.AXYS[3][4] ),
    .X(net95));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(\MOS6502.PC[11] ),
    .X(net194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(_0055_),
    .X(net195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(\MOS6502.PC[13] ),
    .X(net196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(_0057_),
    .X(net197));
 sky130_fd_sc_hd__buf_1 hold114 (.A(\MOS6502.adc_sbc ),
    .X(net198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(_0000_),
    .X(net199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(\MOS6502.PC[15] ),
    .X(net200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(_0059_),
    .X(net201));
 sky130_fd_sc_hd__buf_1 hold118 (.A(\MOS6502.PC[14] ),
    .X(net202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(_0058_),
    .X(net203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(_0147_),
    .X(net96));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(\MOS6502.load_reg ),
    .X(net204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(_0101_),
    .X(net205));
 sky130_fd_sc_hd__buf_1 hold122 (.A(\MOS6502.op[3] ),
    .X(net206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(_0120_),
    .X(net207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(\MOS6502.dst_reg[0] ),
    .X(net208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(\MOS6502.PC[7] ),
    .X(net209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(_0051_),
    .X(net210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(\MOS6502.PC[6] ),
    .X(net211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(_0050_),
    .X(net212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(\MOS6502.PC[3] ),
    .X(net213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\MOS6502.AXYS[0][1] ),
    .X(net97));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(_0047_),
    .X(net214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(\MOS6502.store ),
    .X(net215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(_0107_),
    .X(net216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(\MOS6502.PC[2] ),
    .X(net217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(_0046_),
    .X(net218));
 sky130_fd_sc_hd__buf_1 hold135 (.A(\MOS6502.PC[1] ),
    .X(net219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(_0045_),
    .X(net220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(\MOS6502.PC[4] ),
    .X(net221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(_0048_),
    .X(net222));
 sky130_fd_sc_hd__buf_1 hold139 (.A(\MOS6502.PC[0] ),
    .X(net223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(_0136_),
    .X(net98));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(_0044_),
    .X(net224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(\MOS6502.PC[5] ),
    .X(net225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(_0049_),
    .X(net226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(\MOS6502.op[0] ),
    .X(net227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(\MOS6502.clv ),
    .X(net228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(\MOS6502.inc ),
    .X(net229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(_0385_),
    .X(net230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(net27),
    .X(net231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(_0085_),
    .X(net232));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold149 (.A(\MOS6502.write_back ),
    .X(net233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\MOS6502.AXYS[1][4] ),
    .X(net99));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(_0108_),
    .X(net234));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold151 (.A(net327),
    .X(net235));
 sky130_fd_sc_hd__buf_1 hold152 (.A(net329),
    .X(net236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(\MOS6502.load_only ),
    .X(net237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(\MOS6502.sec ),
    .X(net238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(_0420_),
    .X(net239));
 sky130_fd_sc_hd__buf_1 hold156 (.A(net328),
    .X(net240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(\MOS6502.bit_ins ),
    .X(net241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(_0121_),
    .X(net242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(\MOS6502.op[2] ),
    .X(net243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(_0028_),
    .X(net100));
 sky130_fd_sc_hd__buf_2 hold160 (.A(\MOS6502.ADD[7] ),
    .X(net244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(\MOS6502.index_y ),
    .X(net245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(_0106_),
    .X(net246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(\MOS6502.NMI_1 ),
    .X(net247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(_0424_),
    .X(net248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(_0425_),
    .X(net249));
 sky130_fd_sc_hd__clkbuf_4 hold166 (.A(\MOS6502.plp ),
    .X(net250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(net37),
    .X(net251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(_0087_),
    .X(net252));
 sky130_fd_sc_hd__buf_1 hold169 (.A(\MOS6502.shift_right ),
    .X(net253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\MOS6502.AXYS[3][7] ),
    .X(net101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(_0115_),
    .X(net254));
 sky130_fd_sc_hd__buf_1 hold171 (.A(\MOS6502.ADD[4] ),
    .X(net255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(_0039_),
    .X(net256));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold173 (.A(\MOS6502.compare ),
    .X(net257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(_0114_),
    .X(net258));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold175 (.A(\MOS6502.ADD[0] ),
    .X(net259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(\MOS6502.ABL[0] ),
    .X(net260));
 sky130_fd_sc_hd__buf_1 hold177 (.A(\MOS6502.ADD[1] ),
    .X(net261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(\MOS6502.ABL[6] ),
    .X(net262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(_0289_),
    .X(net263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(_0150_),
    .X(net102));
 sky130_fd_sc_hd__buf_1 hold180 (.A(\MOS6502.ADD[5] ),
    .X(net264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(_0040_),
    .X(net265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(\MOS6502.ABL[4] ),
    .X(net266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(\MOS6502.ABL[5] ),
    .X(net267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(\MOS6502.sei ),
    .X(net268));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold185 (.A(\MOS6502.clc ),
    .X(net269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(\MOS6502.ABL[3] ),
    .X(net270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(_0286_),
    .X(net271));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold188 (.A(\MOS6502.sed ),
    .X(net272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(_0417_),
    .X(net273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\MOS6502.AXYS[1][6] ),
    .X(net103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(\MOS6502.ABL[2] ),
    .X(net274));
 sky130_fd_sc_hd__clkbuf_2 hold191 (.A(\MOS6502.ALU.CO ),
    .X(net275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(_0033_),
    .X(net276));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold193 (.A(\MOS6502.ADD[6] ),
    .X(net277));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold194 (.A(\MOS6502.ADD[3] ),
    .X(net278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(\MOS6502.ABL[7] ),
    .X(net279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(\MOS6502.php ),
    .X(net280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold197 (.A(_0422_),
    .X(net281));
 sky130_fd_sc_hd__buf_1 hold198 (.A(\MOS6502.state[5] ),
    .X(net282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(_0460_),
    .X(net283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(_0094_),
    .X(net86));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(_0030_),
    .X(net104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(\MOS6502.ADD[2] ),
    .X(net284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(\MOS6502.ABL[1] ),
    .X(net285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(\MOS6502.dst_reg[1] ),
    .X(net286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(\MOS6502.rotate ),
    .X(net287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(\MOS6502.ABH[7] ),
    .X(net288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(_0282_),
    .X(net289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(\MOS6502.ABH[6] ),
    .X(net290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(\MOS6502.ABH[4] ),
    .X(net291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(_0279_),
    .X(net292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold209 (.A(\MOS6502.ABH[3] ),
    .X(net293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\MOS6502.AXYS[2][7] ),
    .X(net105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold210 (.A(_0278_),
    .X(net294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(\MOS6502.ABH[5] ),
    .X(net295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(\MOS6502.DIHOLD[4] ),
    .X(net296));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold213 (.A(\MOS6502.cld ),
    .X(net297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold214 (.A(net36),
    .X(net298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(_0390_),
    .X(net299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(\MOS6502.DIHOLD[6] ),
    .X(net300));
 sky130_fd_sc_hd__buf_1 hold217 (.A(_0558_),
    .X(net301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold218 (.A(\MOS6502.ABH[2] ),
    .X(net302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold219 (.A(_0277_),
    .X(net303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(_0015_),
    .X(net106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(\MOS6502.DIHOLD[0] ),
    .X(net304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold221 (.A(\MOS6502.DIHOLD[2] ),
    .X(net305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold222 (.A(\MOS6502.DIHOLD[5] ),
    .X(net306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold223 (.A(_0564_),
    .X(net307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(\MOS6502.DIHOLD[1] ),
    .X(net308));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold225 (.A(_0591_),
    .X(net309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold226 (.A(\MOS6502.DIHOLD[7] ),
    .X(net310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold227 (.A(\MOS6502.ABH[1] ),
    .X(net311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold228 (.A(\MOS6502.DIHOLD[3] ),
    .X(net312));
 sky130_fd_sc_hd__buf_1 hold229 (.A(_0577_),
    .X(net313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\MOS6502.AXYS[0][5] ),
    .X(net107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold230 (.A(\MOS6502.ABH[0] ),
    .X(net314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold231 (.A(_0275_),
    .X(net315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold232 (.A(net38),
    .X(net316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold233 (.A(_0331_),
    .X(net317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold234 (.A(net39),
    .X(net318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold235 (.A(_0314_),
    .X(net319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold236 (.A(net16),
    .X(net320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold237 (.A(_0298_),
    .X(net321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(\MOS6502.state[5] ),
    .X(net322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold239 (.A(\MOS6502.state[0] ),
    .X(net323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(_0140_),
    .X(net108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold240 (.A(_0001_),
    .X(net324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(\MOS6502.IRHOLD[4] ),
    .X(net325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold242 (.A(\MOS6502.res ),
    .X(net326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold243 (.A(\MOS6502.cli ),
    .X(net327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold244 (.A(\MOS6502.shift ),
    .X(net328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold245 (.A(\MOS6502.IRHOLD_valid ),
    .X(net329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\MOS6502.AXYS[3][5] ),
    .X(net109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(_0148_),
    .X(net110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\MOS6502.IRHOLD[5] ),
    .X(net111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(_0096_),
    .X(net112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\MOS6502.AXYS[0][6] ),
    .X(net113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\MOS6502.IRHOLD[1] ),
    .X(net87));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(_0141_),
    .X(net114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\MOS6502.AXYS[1][5] ),
    .X(net115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(_0029_),
    .X(net116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\MOS6502.AXYS[3][3] ),
    .X(net117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(_0146_),
    .X(net118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\MOS6502.AXYS[0][0] ),
    .X(net119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(_0135_),
    .X(net120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\MOS6502.AXYS[3][0] ),
    .X(net121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(_0143_),
    .X(net122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\MOS6502.AXYS[3][2] ),
    .X(net123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(_0092_),
    .X(net88));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(_0145_),
    .X(net124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\MOS6502.AXYS[2][5] ),
    .X(net125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(_0013_),
    .X(net126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\MOS6502.AXYS[2][3] ),
    .X(net127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(_0011_),
    .X(net128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\MOS6502.AXYS[0][7] ),
    .X(net129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(_0142_),
    .X(net130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\MOS6502.AXYS[3][6] ),
    .X(net131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(_0149_),
    .X(net132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\MOS6502.AXYS[0][2] ),
    .X(net133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\MOS6502.AXYS[1][7] ),
    .X(net89));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(_0137_),
    .X(net134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(\MOS6502.AXYS[2][4] ),
    .X(net135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(_0012_),
    .X(net136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\MOS6502.IRHOLD[6] ),
    .X(net137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(_0097_),
    .X(net138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(\MOS6502.AXYS[1][1] ),
    .X(net139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(_0025_),
    .X(net140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(\MOS6502.AXYS[3][1] ),
    .X(net141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(_0144_),
    .X(net142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(\MOS6502.AXYS[1][2] ),
    .X(net143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(_0031_),
    .X(net90));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(_0026_),
    .X(net144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(\MOS6502.src_reg[0] ),
    .X(net145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(_0104_),
    .X(net146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(\MOS6502.AXYS[0][4] ),
    .X(net147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(_0139_),
    .X(net148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(\MOS6502.AXYS[2][0] ),
    .X(net149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(_0008_),
    .X(net150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(\MOS6502.AXYS[2][6] ),
    .X(net151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(_0014_),
    .X(net152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(\MOS6502.AXYS[1][3] ),
    .X(net153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\MOS6502.IRHOLD[7] ),
    .X(net91));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(_0027_),
    .X(net154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(\MOS6502.AXYS[0][3] ),
    .X(net155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(_0138_),
    .X(net156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(\MOS6502.cond_code[1] ),
    .X(net157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(_0132_),
    .X(net158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(\MOS6502.AXYS[2][2] ),
    .X(net159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(_0010_),
    .X(net160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(\MOS6502.AXYS[1][0] ),
    .X(net161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(_0024_),
    .X(net162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(\MOS6502.src_reg[1] ),
    .X(net163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(_0098_),
    .X(net92));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(_0105_),
    .X(net164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(\MOS6502.cond_code[2] ),
    .X(net165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(_0133_),
    .X(net166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(\MOS6502.op[1] ),
    .X(net167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(_0118_),
    .X(net168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(\MOS6502.ALU.BI7 ),
    .X(net169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(_0007_),
    .X(net170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(\MOS6502.cond_code[0] ),
    .X(net171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(_0131_),
    .X(net172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(\MOS6502.ALU.HC ),
    .X(net173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\MOS6502.AXYS[2][1] ),
    .X(net93));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(_0034_),
    .X(net174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(\MOS6502.ALU.AI7 ),
    .X(net175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(_0043_),
    .X(net176));
 sky130_fd_sc_hd__buf_1 hold93 (.A(net326),
    .X(net177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(\MOS6502.DI[0] ),
    .X(net178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(_0091_),
    .X(net179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(\MOS6502.DI[4] ),
    .X(net180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(_0095_),
    .X(net181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(\MOS6502.PC[9] ),
    .X(net182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(_0053_),
    .X(net183));
 sky130_fd_sc_hd__buf_1 input1 (.A(custom_settings[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(io_in[26]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_2 input11 (.A(io_in[28]),
    .X(net11));
 sky130_fd_sc_hd__buf_1 input12 (.A(io_in[29]),
    .X(net12));
 sky130_fd_sc_hd__buf_1 input13 (.A(io_in[30]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_4 input14 (.A(rst_n),
    .X(net14));
 sky130_fd_sc_hd__buf_1 input2 (.A(custom_settings[1]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(io_in[19]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(io_in[20]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(io_in[21]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(io_in[22]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(io_in[23]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(io_in[24]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(io_in[25]),
    .X(net9));
 sky130_fd_sc_hd__buf_4 max_cap47 (.A(_0552_),
    .X(net47));
 sky130_fd_sc_hd__buf_12 output15 (.A(net15),
    .X(io_oeb));
 sky130_fd_sc_hd__buf_12 output16 (.A(net16),
    .X(io_out[0]));
 sky130_fd_sc_hd__buf_12 output17 (.A(net17),
    .X(io_out[10]));
 sky130_fd_sc_hd__buf_12 output18 (.A(net18),
    .X(io_out[11]));
 sky130_fd_sc_hd__buf_12 output19 (.A(net19),
    .X(io_out[12]));
 sky130_fd_sc_hd__buf_12 output20 (.A(net20),
    .X(io_out[13]));
 sky130_fd_sc_hd__buf_12 output21 (.A(net21),
    .X(io_out[14]));
 sky130_fd_sc_hd__buf_12 output22 (.A(net22),
    .X(io_out[15]));
 sky130_fd_sc_hd__buf_12 output23 (.A(net23),
    .X(io_out[16]));
 sky130_fd_sc_hd__buf_12 output24 (.A(net24),
    .X(io_out[17]));
 sky130_fd_sc_hd__buf_12 output25 (.A(net25),
    .X(io_out[18]));
 sky130_fd_sc_hd__buf_12 output26 (.A(net26),
    .X(io_out[19]));
 sky130_fd_sc_hd__buf_12 output27 (.A(net27),
    .X(io_out[1]));
 sky130_fd_sc_hd__buf_12 output28 (.A(net28),
    .X(io_out[20]));
 sky130_fd_sc_hd__buf_12 output29 (.A(net29),
    .X(io_out[21]));
 sky130_fd_sc_hd__buf_12 output30 (.A(net30),
    .X(io_out[22]));
 sky130_fd_sc_hd__buf_12 output31 (.A(net31),
    .X(io_out[23]));
 sky130_fd_sc_hd__buf_12 output32 (.A(net32),
    .X(io_out[24]));
 sky130_fd_sc_hd__buf_12 output33 (.A(net33),
    .X(io_out[25]));
 sky130_fd_sc_hd__buf_12 output34 (.A(net34),
    .X(io_out[26]));
 sky130_fd_sc_hd__buf_1 output35 (.A(net35),
    .X(io_out[27]));
 sky130_fd_sc_hd__buf_12 output36 (.A(net36),
    .X(io_out[2]));
 sky130_fd_sc_hd__buf_12 output37 (.A(net37),
    .X(io_out[31]));
 sky130_fd_sc_hd__buf_12 output38 (.A(net38),
    .X(io_out[32]));
 sky130_fd_sc_hd__buf_12 output39 (.A(net39),
    .X(io_out[33]));
 sky130_fd_sc_hd__buf_12 output40 (.A(net40),
    .X(io_out[3]));
 sky130_fd_sc_hd__buf_12 output41 (.A(net41),
    .X(io_out[4]));
 sky130_fd_sc_hd__buf_12 output42 (.A(net42),
    .X(io_out[5]));
 sky130_fd_sc_hd__buf_12 output43 (.A(net43),
    .X(io_out[6]));
 sky130_fd_sc_hd__buf_12 output44 (.A(net44),
    .X(io_out[7]));
 sky130_fd_sc_hd__buf_12 output45 (.A(net45),
    .X(io_out[8]));
 sky130_fd_sc_hd__buf_12 output46 (.A(net46),
    .X(io_out[9]));
 sky130_fd_sc_hd__clkbuf_2 wire51 (.A(_0478_),
    .X(net51));
 sky130_fd_sc_hd__conb_1 wrapped_6502_80 (.LO(net80));
 sky130_fd_sc_hd__conb_1 wrapped_6502_81 (.LO(net81));
 sky130_fd_sc_hd__conb_1 wrapped_6502_82 (.LO(net82));
 sky130_fd_sc_hd__conb_1 wrapped_6502_83 (.LO(net83));
 sky130_fd_sc_hd__conb_1 wrapped_6502_84 (.LO(net84));
 assign io_out[28] = net80;
 assign io_out[29] = net81;
 assign io_out[30] = net82;
 assign io_out[34] = net83;
 assign io_out[35] = net84;
endmodule

