magic
tech sky130B
magscale 1 2
timestamp 1717545214
<< obsli1 >>
rect 1104 2159 438840 167569
<< obsm1 >>
rect 1104 76 439378 169992
<< metal2 >>
rect 5354 169200 5410 170000
rect 6366 169200 6422 170000
rect 7378 169200 7434 170000
rect 8390 169200 8446 170000
rect 9402 169200 9458 170000
rect 10414 169200 10470 170000
rect 11426 169200 11482 170000
rect 12438 169200 12494 170000
rect 13450 169200 13506 170000
rect 14462 169200 14518 170000
rect 15474 169200 15530 170000
rect 16486 169200 16542 170000
rect 17498 169200 17554 170000
rect 18510 169200 18566 170000
rect 19522 169200 19578 170000
rect 20534 169200 20590 170000
rect 21546 169200 21602 170000
rect 22558 169200 22614 170000
rect 23570 169200 23626 170000
rect 24582 169200 24638 170000
rect 25594 169200 25650 170000
rect 26606 169200 26662 170000
rect 27618 169200 27674 170000
rect 28630 169200 28686 170000
rect 29642 169200 29698 170000
rect 30654 169200 30710 170000
rect 31666 169200 31722 170000
rect 32678 169200 32734 170000
rect 33690 169200 33746 170000
rect 34702 169200 34758 170000
rect 35714 169200 35770 170000
rect 36726 169200 36782 170000
rect 37738 169200 37794 170000
rect 38750 169200 38806 170000
rect 39762 169200 39818 170000
rect 40774 169200 40830 170000
rect 41786 169200 41842 170000
rect 42798 169200 42854 170000
rect 43810 169200 43866 170000
rect 44822 169200 44878 170000
rect 45834 169200 45890 170000
rect 46846 169200 46902 170000
rect 47858 169200 47914 170000
rect 48870 169200 48926 170000
rect 49882 169200 49938 170000
rect 50894 169200 50950 170000
rect 51906 169200 51962 170000
rect 52918 169200 52974 170000
rect 53930 169200 53986 170000
rect 54942 169200 54998 170000
rect 55954 169200 56010 170000
rect 56966 169200 57022 170000
rect 57978 169200 58034 170000
rect 58990 169200 59046 170000
rect 60002 169200 60058 170000
rect 61014 169200 61070 170000
rect 62026 169200 62082 170000
rect 63038 169200 63094 170000
rect 64050 169200 64106 170000
rect 65062 169200 65118 170000
rect 66074 169200 66130 170000
rect 67086 169200 67142 170000
rect 68098 169200 68154 170000
rect 69110 169200 69166 170000
rect 70122 169200 70178 170000
rect 71134 169200 71190 170000
rect 72146 169200 72202 170000
rect 73158 169200 73214 170000
rect 74170 169200 74226 170000
rect 75182 169200 75238 170000
rect 76194 169200 76250 170000
rect 77206 169200 77262 170000
rect 78218 169200 78274 170000
rect 79230 169200 79286 170000
rect 80242 169200 80298 170000
rect 81254 169200 81310 170000
rect 82266 169200 82322 170000
rect 83278 169200 83334 170000
rect 84290 169200 84346 170000
rect 85302 169200 85358 170000
rect 86314 169200 86370 170000
rect 87326 169200 87382 170000
rect 88338 169200 88394 170000
rect 89350 169200 89406 170000
rect 90362 169200 90418 170000
rect 91374 169200 91430 170000
rect 92386 169200 92442 170000
rect 93398 169200 93454 170000
rect 94410 169200 94466 170000
rect 95422 169200 95478 170000
rect 96434 169200 96490 170000
rect 97446 169200 97502 170000
rect 98458 169200 98514 170000
rect 99470 169200 99526 170000
rect 100482 169200 100538 170000
rect 101494 169200 101550 170000
rect 102506 169200 102562 170000
rect 103518 169200 103574 170000
rect 104530 169200 104586 170000
rect 105542 169200 105598 170000
rect 106554 169200 106610 170000
rect 107566 169200 107622 170000
rect 108578 169200 108634 170000
rect 109590 169200 109646 170000
rect 110602 169200 110658 170000
rect 111614 169200 111670 170000
rect 112626 169200 112682 170000
rect 113638 169200 113694 170000
rect 114650 169200 114706 170000
rect 115662 169200 115718 170000
rect 116674 169200 116730 170000
rect 117686 169200 117742 170000
rect 118698 169200 118754 170000
rect 119710 169200 119766 170000
rect 120722 169200 120778 170000
rect 121734 169200 121790 170000
rect 122746 169200 122802 170000
rect 123758 169200 123814 170000
rect 124770 169200 124826 170000
rect 125782 169200 125838 170000
rect 126794 169200 126850 170000
rect 127806 169200 127862 170000
rect 128818 169200 128874 170000
rect 129830 169200 129886 170000
rect 130842 169200 130898 170000
rect 131854 169200 131910 170000
rect 132866 169200 132922 170000
rect 133878 169200 133934 170000
rect 134890 169200 134946 170000
rect 135902 169200 135958 170000
rect 136914 169200 136970 170000
rect 137926 169200 137982 170000
rect 138938 169200 138994 170000
rect 139950 169200 140006 170000
rect 140962 169200 141018 170000
rect 141974 169200 142030 170000
rect 142986 169200 143042 170000
rect 143998 169200 144054 170000
rect 145010 169200 145066 170000
rect 146022 169200 146078 170000
rect 147034 169200 147090 170000
rect 148046 169200 148102 170000
rect 149058 169200 149114 170000
rect 150070 169200 150126 170000
rect 151082 169200 151138 170000
rect 152094 169200 152150 170000
rect 153106 169200 153162 170000
rect 154118 169200 154174 170000
rect 155130 169200 155186 170000
rect 156142 169200 156198 170000
rect 157154 169200 157210 170000
rect 158166 169200 158222 170000
rect 159178 169200 159234 170000
rect 160190 169200 160246 170000
rect 161202 169200 161258 170000
rect 162214 169200 162270 170000
rect 163226 169200 163282 170000
rect 164238 169200 164294 170000
rect 165250 169200 165306 170000
rect 166262 169200 166318 170000
rect 167274 169200 167330 170000
rect 168286 169200 168342 170000
rect 169298 169200 169354 170000
rect 170310 169200 170366 170000
rect 171322 169200 171378 170000
rect 172334 169200 172390 170000
rect 173346 169200 173402 170000
rect 174358 169200 174414 170000
rect 175370 169200 175426 170000
rect 176382 169200 176438 170000
rect 177394 169200 177450 170000
rect 178406 169200 178462 170000
rect 179418 169200 179474 170000
rect 180430 169200 180486 170000
rect 181442 169200 181498 170000
rect 182454 169200 182510 170000
rect 183466 169200 183522 170000
rect 184478 169200 184534 170000
rect 185490 169200 185546 170000
rect 186502 169200 186558 170000
rect 187514 169200 187570 170000
rect 188526 169200 188582 170000
rect 189538 169200 189594 170000
rect 190550 169200 190606 170000
rect 191562 169200 191618 170000
rect 192574 169200 192630 170000
rect 193586 169200 193642 170000
rect 194598 169200 194654 170000
rect 195610 169200 195666 170000
rect 196622 169200 196678 170000
rect 197634 169200 197690 170000
rect 198646 169200 198702 170000
rect 199658 169200 199714 170000
rect 200670 169200 200726 170000
rect 201682 169200 201738 170000
rect 202694 169200 202750 170000
rect 203706 169200 203762 170000
rect 204718 169200 204774 170000
rect 205730 169200 205786 170000
rect 206742 169200 206798 170000
rect 207754 169200 207810 170000
rect 208766 169200 208822 170000
rect 209778 169200 209834 170000
rect 210790 169200 210846 170000
rect 211802 169200 211858 170000
rect 212814 169200 212870 170000
rect 213826 169200 213882 170000
rect 214838 169200 214894 170000
rect 215850 169200 215906 170000
rect 216862 169200 216918 170000
rect 217874 169200 217930 170000
rect 218886 169200 218942 170000
rect 219898 169200 219954 170000
rect 220910 169200 220966 170000
rect 221922 169200 221978 170000
rect 222934 169200 222990 170000
rect 223946 169200 224002 170000
rect 224958 169200 225014 170000
rect 225970 169200 226026 170000
rect 226982 169200 227038 170000
rect 227994 169200 228050 170000
rect 229006 169200 229062 170000
rect 230018 169200 230074 170000
rect 231030 169200 231086 170000
rect 232042 169200 232098 170000
rect 233054 169200 233110 170000
rect 234066 169200 234122 170000
rect 235078 169200 235134 170000
rect 236090 169200 236146 170000
rect 237102 169200 237158 170000
rect 238114 169200 238170 170000
rect 239126 169200 239182 170000
rect 240138 169200 240194 170000
rect 241150 169200 241206 170000
rect 242162 169200 242218 170000
rect 243174 169200 243230 170000
rect 244186 169200 244242 170000
rect 245198 169200 245254 170000
rect 246210 169200 246266 170000
rect 247222 169200 247278 170000
rect 248234 169200 248290 170000
rect 249246 169200 249302 170000
rect 250258 169200 250314 170000
rect 251270 169200 251326 170000
rect 252282 169200 252338 170000
rect 253294 169200 253350 170000
rect 254306 169200 254362 170000
rect 255318 169200 255374 170000
rect 256330 169200 256386 170000
rect 257342 169200 257398 170000
rect 258354 169200 258410 170000
rect 259366 169200 259422 170000
rect 260378 169200 260434 170000
rect 261390 169200 261446 170000
rect 262402 169200 262458 170000
rect 263414 169200 263470 170000
rect 264426 169200 264482 170000
rect 265438 169200 265494 170000
rect 266450 169200 266506 170000
rect 267462 169200 267518 170000
rect 268474 169200 268530 170000
rect 269486 169200 269542 170000
rect 270498 169200 270554 170000
rect 271510 169200 271566 170000
rect 272522 169200 272578 170000
rect 273534 169200 273590 170000
rect 274546 169200 274602 170000
rect 275558 169200 275614 170000
rect 276570 169200 276626 170000
rect 277582 169200 277638 170000
rect 278594 169200 278650 170000
rect 279606 169200 279662 170000
rect 280618 169200 280674 170000
rect 281630 169200 281686 170000
rect 282642 169200 282698 170000
rect 283654 169200 283710 170000
rect 284666 169200 284722 170000
rect 285678 169200 285734 170000
rect 286690 169200 286746 170000
rect 287702 169200 287758 170000
rect 288714 169200 288770 170000
rect 289726 169200 289782 170000
rect 290738 169200 290794 170000
rect 291750 169200 291806 170000
rect 292762 169200 292818 170000
rect 293774 169200 293830 170000
rect 294786 169200 294842 170000
rect 295798 169200 295854 170000
rect 296810 169200 296866 170000
rect 297822 169200 297878 170000
rect 298834 169200 298890 170000
rect 299846 169200 299902 170000
rect 300858 169200 300914 170000
rect 301870 169200 301926 170000
rect 302882 169200 302938 170000
rect 303894 169200 303950 170000
rect 304906 169200 304962 170000
rect 305918 169200 305974 170000
rect 306930 169200 306986 170000
rect 307942 169200 307998 170000
rect 308954 169200 309010 170000
rect 309966 169200 310022 170000
rect 310978 169200 311034 170000
rect 311990 169200 312046 170000
rect 313002 169200 313058 170000
rect 314014 169200 314070 170000
rect 315026 169200 315082 170000
rect 316038 169200 316094 170000
rect 317050 169200 317106 170000
rect 318062 169200 318118 170000
rect 319074 169200 319130 170000
rect 320086 169200 320142 170000
rect 321098 169200 321154 170000
rect 322110 169200 322166 170000
rect 323122 169200 323178 170000
rect 324134 169200 324190 170000
rect 325146 169200 325202 170000
rect 326158 169200 326214 170000
rect 327170 169200 327226 170000
rect 328182 169200 328238 170000
rect 329194 169200 329250 170000
rect 330206 169200 330262 170000
rect 331218 169200 331274 170000
rect 332230 169200 332286 170000
rect 333242 169200 333298 170000
rect 334254 169200 334310 170000
rect 335266 169200 335322 170000
rect 336278 169200 336334 170000
rect 337290 169200 337346 170000
rect 338302 169200 338358 170000
rect 339314 169200 339370 170000
rect 340326 169200 340382 170000
rect 341338 169200 341394 170000
rect 342350 169200 342406 170000
rect 343362 169200 343418 170000
rect 344374 169200 344430 170000
rect 345386 169200 345442 170000
rect 346398 169200 346454 170000
rect 347410 169200 347466 170000
rect 348422 169200 348478 170000
rect 349434 169200 349490 170000
rect 350446 169200 350502 170000
rect 351458 169200 351514 170000
rect 352470 169200 352526 170000
rect 353482 169200 353538 170000
rect 354494 169200 354550 170000
rect 355506 169200 355562 170000
rect 356518 169200 356574 170000
rect 357530 169200 357586 170000
rect 358542 169200 358598 170000
rect 359554 169200 359610 170000
rect 360566 169200 360622 170000
rect 361578 169200 361634 170000
rect 362590 169200 362646 170000
rect 363602 169200 363658 170000
rect 364614 169200 364670 170000
rect 365626 169200 365682 170000
rect 366638 169200 366694 170000
rect 367650 169200 367706 170000
rect 368662 169200 368718 170000
rect 369674 169200 369730 170000
rect 370686 169200 370742 170000
rect 371698 169200 371754 170000
rect 372710 169200 372766 170000
rect 373722 169200 373778 170000
rect 374734 169200 374790 170000
rect 375746 169200 375802 170000
rect 376758 169200 376814 170000
rect 377770 169200 377826 170000
rect 378782 169200 378838 170000
rect 379794 169200 379850 170000
rect 380806 169200 380862 170000
rect 381818 169200 381874 170000
rect 382830 169200 382886 170000
rect 383842 169200 383898 170000
rect 384854 169200 384910 170000
rect 385866 169200 385922 170000
rect 386878 169200 386934 170000
rect 387890 169200 387946 170000
rect 388902 169200 388958 170000
rect 389914 169200 389970 170000
rect 390926 169200 390982 170000
rect 391938 169200 391994 170000
rect 392950 169200 393006 170000
rect 393962 169200 394018 170000
rect 394974 169200 395030 170000
rect 395986 169200 396042 170000
rect 396998 169200 397054 170000
rect 398010 169200 398066 170000
rect 399022 169200 399078 170000
rect 400034 169200 400090 170000
rect 401046 169200 401102 170000
rect 402058 169200 402114 170000
rect 403070 169200 403126 170000
rect 404082 169200 404138 170000
rect 405094 169200 405150 170000
rect 406106 169200 406162 170000
rect 407118 169200 407174 170000
rect 408130 169200 408186 170000
rect 409142 169200 409198 170000
rect 410154 169200 410210 170000
rect 411166 169200 411222 170000
rect 412178 169200 412234 170000
rect 413190 169200 413246 170000
rect 414202 169200 414258 170000
rect 415214 169200 415270 170000
rect 416226 169200 416282 170000
rect 417238 169200 417294 170000
rect 418250 169200 418306 170000
rect 419262 169200 419318 170000
rect 420274 169200 420330 170000
rect 421286 169200 421342 170000
rect 422298 169200 422354 170000
rect 423310 169200 423366 170000
rect 424322 169200 424378 170000
rect 425334 169200 425390 170000
rect 426346 169200 426402 170000
rect 427358 169200 427414 170000
rect 428370 169200 428426 170000
rect 429382 169200 429438 170000
rect 430394 169200 430450 170000
rect 431406 169200 431462 170000
rect 432418 169200 432474 170000
rect 433430 169200 433486 170000
rect 434442 169200 434498 170000
rect 8390 0 8446 800
rect 10138 0 10194 800
rect 11886 0 11942 800
rect 13634 0 13690 800
rect 15382 0 15438 800
rect 17130 0 17186 800
rect 18878 0 18934 800
rect 20626 0 20682 800
rect 22374 0 22430 800
rect 24122 0 24178 800
rect 25870 0 25926 800
rect 27618 0 27674 800
rect 29366 0 29422 800
rect 31114 0 31170 800
rect 32862 0 32918 800
rect 34610 0 34666 800
rect 36358 0 36414 800
rect 38106 0 38162 800
rect 39854 0 39910 800
rect 41602 0 41658 800
rect 43350 0 43406 800
rect 45098 0 45154 800
rect 46846 0 46902 800
rect 48594 0 48650 800
rect 50342 0 50398 800
rect 52090 0 52146 800
rect 53838 0 53894 800
rect 55586 0 55642 800
rect 57334 0 57390 800
rect 59082 0 59138 800
rect 60830 0 60886 800
rect 62578 0 62634 800
rect 64326 0 64382 800
rect 66074 0 66130 800
rect 67822 0 67878 800
rect 69570 0 69626 800
rect 71318 0 71374 800
rect 73066 0 73122 800
rect 74814 0 74870 800
rect 76562 0 76618 800
rect 78310 0 78366 800
rect 80058 0 80114 800
rect 81806 0 81862 800
rect 83554 0 83610 800
rect 85302 0 85358 800
rect 87050 0 87106 800
rect 88798 0 88854 800
rect 90546 0 90602 800
rect 92294 0 92350 800
rect 94042 0 94098 800
rect 95790 0 95846 800
rect 97538 0 97594 800
rect 99286 0 99342 800
rect 101034 0 101090 800
rect 102782 0 102838 800
rect 104530 0 104586 800
rect 106278 0 106334 800
rect 108026 0 108082 800
rect 109774 0 109830 800
rect 111522 0 111578 800
rect 113270 0 113326 800
rect 115018 0 115074 800
rect 116766 0 116822 800
rect 118514 0 118570 800
rect 120262 0 120318 800
rect 122010 0 122066 800
rect 123758 0 123814 800
rect 125506 0 125562 800
rect 127254 0 127310 800
rect 129002 0 129058 800
rect 130750 0 130806 800
rect 132498 0 132554 800
rect 134246 0 134302 800
rect 135994 0 136050 800
rect 137742 0 137798 800
rect 139490 0 139546 800
rect 141238 0 141294 800
rect 142986 0 143042 800
rect 144734 0 144790 800
rect 146482 0 146538 800
rect 148230 0 148286 800
rect 149978 0 150034 800
rect 151726 0 151782 800
rect 153474 0 153530 800
rect 155222 0 155278 800
rect 156970 0 157026 800
rect 158718 0 158774 800
rect 160466 0 160522 800
rect 162214 0 162270 800
rect 163962 0 164018 800
rect 165710 0 165766 800
rect 167458 0 167514 800
rect 169206 0 169262 800
rect 170954 0 171010 800
rect 172702 0 172758 800
rect 174450 0 174506 800
rect 176198 0 176254 800
rect 177946 0 178002 800
rect 179694 0 179750 800
rect 181442 0 181498 800
rect 183190 0 183246 800
rect 184938 0 184994 800
rect 186686 0 186742 800
rect 188434 0 188490 800
rect 190182 0 190238 800
rect 191930 0 191986 800
rect 193678 0 193734 800
rect 195426 0 195482 800
rect 197174 0 197230 800
rect 198922 0 198978 800
rect 200670 0 200726 800
rect 202418 0 202474 800
rect 204166 0 204222 800
rect 205914 0 205970 800
rect 207662 0 207718 800
rect 209410 0 209466 800
rect 211158 0 211214 800
rect 212906 0 212962 800
rect 214654 0 214710 800
rect 216402 0 216458 800
rect 218150 0 218206 800
rect 219898 0 219954 800
rect 221646 0 221702 800
rect 223394 0 223450 800
rect 225142 0 225198 800
rect 226890 0 226946 800
rect 228638 0 228694 800
rect 230386 0 230442 800
rect 232134 0 232190 800
rect 233882 0 233938 800
rect 235630 0 235686 800
rect 237378 0 237434 800
rect 239126 0 239182 800
rect 240874 0 240930 800
rect 242622 0 242678 800
rect 244370 0 244426 800
rect 246118 0 246174 800
rect 247866 0 247922 800
rect 249614 0 249670 800
rect 251362 0 251418 800
rect 253110 0 253166 800
rect 254858 0 254914 800
rect 256606 0 256662 800
rect 258354 0 258410 800
rect 260102 0 260158 800
rect 261850 0 261906 800
rect 263598 0 263654 800
rect 265346 0 265402 800
rect 267094 0 267150 800
rect 268842 0 268898 800
rect 270590 0 270646 800
rect 272338 0 272394 800
rect 274086 0 274142 800
rect 275834 0 275890 800
rect 277582 0 277638 800
rect 279330 0 279386 800
rect 281078 0 281134 800
rect 282826 0 282882 800
rect 284574 0 284630 800
rect 286322 0 286378 800
rect 288070 0 288126 800
rect 289818 0 289874 800
rect 291566 0 291622 800
rect 293314 0 293370 800
rect 295062 0 295118 800
rect 296810 0 296866 800
rect 298558 0 298614 800
rect 300306 0 300362 800
rect 302054 0 302110 800
rect 303802 0 303858 800
rect 305550 0 305606 800
rect 307298 0 307354 800
rect 309046 0 309102 800
rect 310794 0 310850 800
rect 312542 0 312598 800
rect 314290 0 314346 800
rect 316038 0 316094 800
rect 317786 0 317842 800
rect 319534 0 319590 800
rect 321282 0 321338 800
rect 323030 0 323086 800
rect 324778 0 324834 800
rect 326526 0 326582 800
rect 328274 0 328330 800
rect 330022 0 330078 800
rect 331770 0 331826 800
rect 333518 0 333574 800
rect 335266 0 335322 800
rect 337014 0 337070 800
rect 338762 0 338818 800
rect 340510 0 340566 800
rect 342258 0 342314 800
rect 344006 0 344062 800
rect 345754 0 345810 800
rect 347502 0 347558 800
rect 349250 0 349306 800
rect 350998 0 351054 800
rect 352746 0 352802 800
rect 354494 0 354550 800
rect 356242 0 356298 800
rect 357990 0 358046 800
rect 359738 0 359794 800
rect 361486 0 361542 800
rect 363234 0 363290 800
rect 364982 0 365038 800
rect 366730 0 366786 800
rect 368478 0 368534 800
rect 370226 0 370282 800
rect 371974 0 372030 800
rect 373722 0 373778 800
rect 375470 0 375526 800
rect 377218 0 377274 800
rect 378966 0 379022 800
rect 380714 0 380770 800
rect 382462 0 382518 800
rect 384210 0 384266 800
rect 385958 0 386014 800
rect 387706 0 387762 800
rect 389454 0 389510 800
rect 391202 0 391258 800
rect 392950 0 393006 800
rect 394698 0 394754 800
rect 396446 0 396502 800
rect 398194 0 398250 800
rect 399942 0 399998 800
rect 401690 0 401746 800
rect 403438 0 403494 800
rect 405186 0 405242 800
rect 406934 0 406990 800
rect 408682 0 408738 800
rect 410430 0 410486 800
rect 412178 0 412234 800
rect 413926 0 413982 800
rect 415674 0 415730 800
rect 417422 0 417478 800
rect 419170 0 419226 800
rect 420918 0 420974 800
rect 422666 0 422722 800
rect 424414 0 424470 800
rect 426162 0 426218 800
rect 427910 0 427966 800
rect 429658 0 429714 800
rect 431406 0 431462 800
<< obsm2 >>
rect 1214 169144 5298 169998
rect 5466 169144 6310 169998
rect 6478 169144 7322 169998
rect 7490 169144 8334 169998
rect 8502 169144 9346 169998
rect 9514 169144 10358 169998
rect 10526 169144 11370 169998
rect 11538 169144 12382 169998
rect 12550 169144 13394 169998
rect 13562 169144 14406 169998
rect 14574 169144 15418 169998
rect 15586 169144 16430 169998
rect 16598 169144 17442 169998
rect 17610 169144 18454 169998
rect 18622 169144 19466 169998
rect 19634 169144 20478 169998
rect 20646 169144 21490 169998
rect 21658 169144 22502 169998
rect 22670 169144 23514 169998
rect 23682 169144 24526 169998
rect 24694 169144 25538 169998
rect 25706 169144 26550 169998
rect 26718 169144 27562 169998
rect 27730 169144 28574 169998
rect 28742 169144 29586 169998
rect 29754 169144 30598 169998
rect 30766 169144 31610 169998
rect 31778 169144 32622 169998
rect 32790 169144 33634 169998
rect 33802 169144 34646 169998
rect 34814 169144 35658 169998
rect 35826 169144 36670 169998
rect 36838 169144 37682 169998
rect 37850 169144 38694 169998
rect 38862 169144 39706 169998
rect 39874 169144 40718 169998
rect 40886 169144 41730 169998
rect 41898 169144 42742 169998
rect 42910 169144 43754 169998
rect 43922 169144 44766 169998
rect 44934 169144 45778 169998
rect 45946 169144 46790 169998
rect 46958 169144 47802 169998
rect 47970 169144 48814 169998
rect 48982 169144 49826 169998
rect 49994 169144 50838 169998
rect 51006 169144 51850 169998
rect 52018 169144 52862 169998
rect 53030 169144 53874 169998
rect 54042 169144 54886 169998
rect 55054 169144 55898 169998
rect 56066 169144 56910 169998
rect 57078 169144 57922 169998
rect 58090 169144 58934 169998
rect 59102 169144 59946 169998
rect 60114 169144 60958 169998
rect 61126 169144 61970 169998
rect 62138 169144 62982 169998
rect 63150 169144 63994 169998
rect 64162 169144 65006 169998
rect 65174 169144 66018 169998
rect 66186 169144 67030 169998
rect 67198 169144 68042 169998
rect 68210 169144 69054 169998
rect 69222 169144 70066 169998
rect 70234 169144 71078 169998
rect 71246 169144 72090 169998
rect 72258 169144 73102 169998
rect 73270 169144 74114 169998
rect 74282 169144 75126 169998
rect 75294 169144 76138 169998
rect 76306 169144 77150 169998
rect 77318 169144 78162 169998
rect 78330 169144 79174 169998
rect 79342 169144 80186 169998
rect 80354 169144 81198 169998
rect 81366 169144 82210 169998
rect 82378 169144 83222 169998
rect 83390 169144 84234 169998
rect 84402 169144 85246 169998
rect 85414 169144 86258 169998
rect 86426 169144 87270 169998
rect 87438 169144 88282 169998
rect 88450 169144 89294 169998
rect 89462 169144 90306 169998
rect 90474 169144 91318 169998
rect 91486 169144 92330 169998
rect 92498 169144 93342 169998
rect 93510 169144 94354 169998
rect 94522 169144 95366 169998
rect 95534 169144 96378 169998
rect 96546 169144 97390 169998
rect 97558 169144 98402 169998
rect 98570 169144 99414 169998
rect 99582 169144 100426 169998
rect 100594 169144 101438 169998
rect 101606 169144 102450 169998
rect 102618 169144 103462 169998
rect 103630 169144 104474 169998
rect 104642 169144 105486 169998
rect 105654 169144 106498 169998
rect 106666 169144 107510 169998
rect 107678 169144 108522 169998
rect 108690 169144 109534 169998
rect 109702 169144 110546 169998
rect 110714 169144 111558 169998
rect 111726 169144 112570 169998
rect 112738 169144 113582 169998
rect 113750 169144 114594 169998
rect 114762 169144 115606 169998
rect 115774 169144 116618 169998
rect 116786 169144 117630 169998
rect 117798 169144 118642 169998
rect 118810 169144 119654 169998
rect 119822 169144 120666 169998
rect 120834 169144 121678 169998
rect 121846 169144 122690 169998
rect 122858 169144 123702 169998
rect 123870 169144 124714 169998
rect 124882 169144 125726 169998
rect 125894 169144 126738 169998
rect 126906 169144 127750 169998
rect 127918 169144 128762 169998
rect 128930 169144 129774 169998
rect 129942 169144 130786 169998
rect 130954 169144 131798 169998
rect 131966 169144 132810 169998
rect 132978 169144 133822 169998
rect 133990 169144 134834 169998
rect 135002 169144 135846 169998
rect 136014 169144 136858 169998
rect 137026 169144 137870 169998
rect 138038 169144 138882 169998
rect 139050 169144 139894 169998
rect 140062 169144 140906 169998
rect 141074 169144 141918 169998
rect 142086 169144 142930 169998
rect 143098 169144 143942 169998
rect 144110 169144 144954 169998
rect 145122 169144 145966 169998
rect 146134 169144 146978 169998
rect 147146 169144 147990 169998
rect 148158 169144 149002 169998
rect 149170 169144 150014 169998
rect 150182 169144 151026 169998
rect 151194 169144 152038 169998
rect 152206 169144 153050 169998
rect 153218 169144 154062 169998
rect 154230 169144 155074 169998
rect 155242 169144 156086 169998
rect 156254 169144 157098 169998
rect 157266 169144 158110 169998
rect 158278 169144 159122 169998
rect 159290 169144 160134 169998
rect 160302 169144 161146 169998
rect 161314 169144 162158 169998
rect 162326 169144 163170 169998
rect 163338 169144 164182 169998
rect 164350 169144 165194 169998
rect 165362 169144 166206 169998
rect 166374 169144 167218 169998
rect 167386 169144 168230 169998
rect 168398 169144 169242 169998
rect 169410 169144 170254 169998
rect 170422 169144 171266 169998
rect 171434 169144 172278 169998
rect 172446 169144 173290 169998
rect 173458 169144 174302 169998
rect 174470 169144 175314 169998
rect 175482 169144 176326 169998
rect 176494 169144 177338 169998
rect 177506 169144 178350 169998
rect 178518 169144 179362 169998
rect 179530 169144 180374 169998
rect 180542 169144 181386 169998
rect 181554 169144 182398 169998
rect 182566 169144 183410 169998
rect 183578 169144 184422 169998
rect 184590 169144 185434 169998
rect 185602 169144 186446 169998
rect 186614 169144 187458 169998
rect 187626 169144 188470 169998
rect 188638 169144 189482 169998
rect 189650 169144 190494 169998
rect 190662 169144 191506 169998
rect 191674 169144 192518 169998
rect 192686 169144 193530 169998
rect 193698 169144 194542 169998
rect 194710 169144 195554 169998
rect 195722 169144 196566 169998
rect 196734 169144 197578 169998
rect 197746 169144 198590 169998
rect 198758 169144 199602 169998
rect 199770 169144 200614 169998
rect 200782 169144 201626 169998
rect 201794 169144 202638 169998
rect 202806 169144 203650 169998
rect 203818 169144 204662 169998
rect 204830 169144 205674 169998
rect 205842 169144 206686 169998
rect 206854 169144 207698 169998
rect 207866 169144 208710 169998
rect 208878 169144 209722 169998
rect 209890 169144 210734 169998
rect 210902 169144 211746 169998
rect 211914 169144 212758 169998
rect 212926 169144 213770 169998
rect 213938 169144 214782 169998
rect 214950 169144 215794 169998
rect 215962 169144 216806 169998
rect 216974 169144 217818 169998
rect 217986 169144 218830 169998
rect 218998 169144 219842 169998
rect 220010 169144 220854 169998
rect 221022 169144 221866 169998
rect 222034 169144 222878 169998
rect 223046 169144 223890 169998
rect 224058 169144 224902 169998
rect 225070 169144 225914 169998
rect 226082 169144 226926 169998
rect 227094 169144 227938 169998
rect 228106 169144 228950 169998
rect 229118 169144 229962 169998
rect 230130 169144 230974 169998
rect 231142 169144 231986 169998
rect 232154 169144 232998 169998
rect 233166 169144 234010 169998
rect 234178 169144 235022 169998
rect 235190 169144 236034 169998
rect 236202 169144 237046 169998
rect 237214 169144 238058 169998
rect 238226 169144 239070 169998
rect 239238 169144 240082 169998
rect 240250 169144 241094 169998
rect 241262 169144 242106 169998
rect 242274 169144 243118 169998
rect 243286 169144 244130 169998
rect 244298 169144 245142 169998
rect 245310 169144 246154 169998
rect 246322 169144 247166 169998
rect 247334 169144 248178 169998
rect 248346 169144 249190 169998
rect 249358 169144 250202 169998
rect 250370 169144 251214 169998
rect 251382 169144 252226 169998
rect 252394 169144 253238 169998
rect 253406 169144 254250 169998
rect 254418 169144 255262 169998
rect 255430 169144 256274 169998
rect 256442 169144 257286 169998
rect 257454 169144 258298 169998
rect 258466 169144 259310 169998
rect 259478 169144 260322 169998
rect 260490 169144 261334 169998
rect 261502 169144 262346 169998
rect 262514 169144 263358 169998
rect 263526 169144 264370 169998
rect 264538 169144 265382 169998
rect 265550 169144 266394 169998
rect 266562 169144 267406 169998
rect 267574 169144 268418 169998
rect 268586 169144 269430 169998
rect 269598 169144 270442 169998
rect 270610 169144 271454 169998
rect 271622 169144 272466 169998
rect 272634 169144 273478 169998
rect 273646 169144 274490 169998
rect 274658 169144 275502 169998
rect 275670 169144 276514 169998
rect 276682 169144 277526 169998
rect 277694 169144 278538 169998
rect 278706 169144 279550 169998
rect 279718 169144 280562 169998
rect 280730 169144 281574 169998
rect 281742 169144 282586 169998
rect 282754 169144 283598 169998
rect 283766 169144 284610 169998
rect 284778 169144 285622 169998
rect 285790 169144 286634 169998
rect 286802 169144 287646 169998
rect 287814 169144 288658 169998
rect 288826 169144 289670 169998
rect 289838 169144 290682 169998
rect 290850 169144 291694 169998
rect 291862 169144 292706 169998
rect 292874 169144 293718 169998
rect 293886 169144 294730 169998
rect 294898 169144 295742 169998
rect 295910 169144 296754 169998
rect 296922 169144 297766 169998
rect 297934 169144 298778 169998
rect 298946 169144 299790 169998
rect 299958 169144 300802 169998
rect 300970 169144 301814 169998
rect 301982 169144 302826 169998
rect 302994 169144 303838 169998
rect 304006 169144 304850 169998
rect 305018 169144 305862 169998
rect 306030 169144 306874 169998
rect 307042 169144 307886 169998
rect 308054 169144 308898 169998
rect 309066 169144 309910 169998
rect 310078 169144 310922 169998
rect 311090 169144 311934 169998
rect 312102 169144 312946 169998
rect 313114 169144 313958 169998
rect 314126 169144 314970 169998
rect 315138 169144 315982 169998
rect 316150 169144 316994 169998
rect 317162 169144 318006 169998
rect 318174 169144 319018 169998
rect 319186 169144 320030 169998
rect 320198 169144 321042 169998
rect 321210 169144 322054 169998
rect 322222 169144 323066 169998
rect 323234 169144 324078 169998
rect 324246 169144 325090 169998
rect 325258 169144 326102 169998
rect 326270 169144 327114 169998
rect 327282 169144 328126 169998
rect 328294 169144 329138 169998
rect 329306 169144 330150 169998
rect 330318 169144 331162 169998
rect 331330 169144 332174 169998
rect 332342 169144 333186 169998
rect 333354 169144 334198 169998
rect 334366 169144 335210 169998
rect 335378 169144 336222 169998
rect 336390 169144 337234 169998
rect 337402 169144 338246 169998
rect 338414 169144 339258 169998
rect 339426 169144 340270 169998
rect 340438 169144 341282 169998
rect 341450 169144 342294 169998
rect 342462 169144 343306 169998
rect 343474 169144 344318 169998
rect 344486 169144 345330 169998
rect 345498 169144 346342 169998
rect 346510 169144 347354 169998
rect 347522 169144 348366 169998
rect 348534 169144 349378 169998
rect 349546 169144 350390 169998
rect 350558 169144 351402 169998
rect 351570 169144 352414 169998
rect 352582 169144 353426 169998
rect 353594 169144 354438 169998
rect 354606 169144 355450 169998
rect 355618 169144 356462 169998
rect 356630 169144 357474 169998
rect 357642 169144 358486 169998
rect 358654 169144 359498 169998
rect 359666 169144 360510 169998
rect 360678 169144 361522 169998
rect 361690 169144 362534 169998
rect 362702 169144 363546 169998
rect 363714 169144 364558 169998
rect 364726 169144 365570 169998
rect 365738 169144 366582 169998
rect 366750 169144 367594 169998
rect 367762 169144 368606 169998
rect 368774 169144 369618 169998
rect 369786 169144 370630 169998
rect 370798 169144 371642 169998
rect 371810 169144 372654 169998
rect 372822 169144 373666 169998
rect 373834 169144 374678 169998
rect 374846 169144 375690 169998
rect 375858 169144 376702 169998
rect 376870 169144 377714 169998
rect 377882 169144 378726 169998
rect 378894 169144 379738 169998
rect 379906 169144 380750 169998
rect 380918 169144 381762 169998
rect 381930 169144 382774 169998
rect 382942 169144 383786 169998
rect 383954 169144 384798 169998
rect 384966 169144 385810 169998
rect 385978 169144 386822 169998
rect 386990 169144 387834 169998
rect 388002 169144 388846 169998
rect 389014 169144 389858 169998
rect 390026 169144 390870 169998
rect 391038 169144 391882 169998
rect 392050 169144 392894 169998
rect 393062 169144 393906 169998
rect 394074 169144 394918 169998
rect 395086 169144 395930 169998
rect 396098 169144 396942 169998
rect 397110 169144 397954 169998
rect 398122 169144 398966 169998
rect 399134 169144 399978 169998
rect 400146 169144 400990 169998
rect 401158 169144 402002 169998
rect 402170 169144 403014 169998
rect 403182 169144 404026 169998
rect 404194 169144 405038 169998
rect 405206 169144 406050 169998
rect 406218 169144 407062 169998
rect 407230 169144 408074 169998
rect 408242 169144 409086 169998
rect 409254 169144 410098 169998
rect 410266 169144 411110 169998
rect 411278 169144 412122 169998
rect 412290 169144 413134 169998
rect 413302 169144 414146 169998
rect 414314 169144 415158 169998
rect 415326 169144 416170 169998
rect 416338 169144 417182 169998
rect 417350 169144 418194 169998
rect 418362 169144 419206 169998
rect 419374 169144 420218 169998
rect 420386 169144 421230 169998
rect 421398 169144 422242 169998
rect 422410 169144 423254 169998
rect 423422 169144 424266 169998
rect 424434 169144 425278 169998
rect 425446 169144 426290 169998
rect 426458 169144 427302 169998
rect 427470 169144 428314 169998
rect 428482 169144 429326 169998
rect 429494 169144 430338 169998
rect 430506 169144 431350 169998
rect 431518 169144 432362 169998
rect 432530 169144 433374 169998
rect 433542 169144 434386 169998
rect 434554 169144 439372 169998
rect 1214 856 439372 169144
rect 1214 31 8334 856
rect 8502 31 10082 856
rect 10250 31 11830 856
rect 11998 31 13578 856
rect 13746 31 15326 856
rect 15494 31 17074 856
rect 17242 31 18822 856
rect 18990 31 20570 856
rect 20738 31 22318 856
rect 22486 31 24066 856
rect 24234 31 25814 856
rect 25982 31 27562 856
rect 27730 31 29310 856
rect 29478 31 31058 856
rect 31226 31 32806 856
rect 32974 31 34554 856
rect 34722 31 36302 856
rect 36470 31 38050 856
rect 38218 31 39798 856
rect 39966 31 41546 856
rect 41714 31 43294 856
rect 43462 31 45042 856
rect 45210 31 46790 856
rect 46958 31 48538 856
rect 48706 31 50286 856
rect 50454 31 52034 856
rect 52202 31 53782 856
rect 53950 31 55530 856
rect 55698 31 57278 856
rect 57446 31 59026 856
rect 59194 31 60774 856
rect 60942 31 62522 856
rect 62690 31 64270 856
rect 64438 31 66018 856
rect 66186 31 67766 856
rect 67934 31 69514 856
rect 69682 31 71262 856
rect 71430 31 73010 856
rect 73178 31 74758 856
rect 74926 31 76506 856
rect 76674 31 78254 856
rect 78422 31 80002 856
rect 80170 31 81750 856
rect 81918 31 83498 856
rect 83666 31 85246 856
rect 85414 31 86994 856
rect 87162 31 88742 856
rect 88910 31 90490 856
rect 90658 31 92238 856
rect 92406 31 93986 856
rect 94154 31 95734 856
rect 95902 31 97482 856
rect 97650 31 99230 856
rect 99398 31 100978 856
rect 101146 31 102726 856
rect 102894 31 104474 856
rect 104642 31 106222 856
rect 106390 31 107970 856
rect 108138 31 109718 856
rect 109886 31 111466 856
rect 111634 31 113214 856
rect 113382 31 114962 856
rect 115130 31 116710 856
rect 116878 31 118458 856
rect 118626 31 120206 856
rect 120374 31 121954 856
rect 122122 31 123702 856
rect 123870 31 125450 856
rect 125618 31 127198 856
rect 127366 31 128946 856
rect 129114 31 130694 856
rect 130862 31 132442 856
rect 132610 31 134190 856
rect 134358 31 135938 856
rect 136106 31 137686 856
rect 137854 31 139434 856
rect 139602 31 141182 856
rect 141350 31 142930 856
rect 143098 31 144678 856
rect 144846 31 146426 856
rect 146594 31 148174 856
rect 148342 31 149922 856
rect 150090 31 151670 856
rect 151838 31 153418 856
rect 153586 31 155166 856
rect 155334 31 156914 856
rect 157082 31 158662 856
rect 158830 31 160410 856
rect 160578 31 162158 856
rect 162326 31 163906 856
rect 164074 31 165654 856
rect 165822 31 167402 856
rect 167570 31 169150 856
rect 169318 31 170898 856
rect 171066 31 172646 856
rect 172814 31 174394 856
rect 174562 31 176142 856
rect 176310 31 177890 856
rect 178058 31 179638 856
rect 179806 31 181386 856
rect 181554 31 183134 856
rect 183302 31 184882 856
rect 185050 31 186630 856
rect 186798 31 188378 856
rect 188546 31 190126 856
rect 190294 31 191874 856
rect 192042 31 193622 856
rect 193790 31 195370 856
rect 195538 31 197118 856
rect 197286 31 198866 856
rect 199034 31 200614 856
rect 200782 31 202362 856
rect 202530 31 204110 856
rect 204278 31 205858 856
rect 206026 31 207606 856
rect 207774 31 209354 856
rect 209522 31 211102 856
rect 211270 31 212850 856
rect 213018 31 214598 856
rect 214766 31 216346 856
rect 216514 31 218094 856
rect 218262 31 219842 856
rect 220010 31 221590 856
rect 221758 31 223338 856
rect 223506 31 225086 856
rect 225254 31 226834 856
rect 227002 31 228582 856
rect 228750 31 230330 856
rect 230498 31 232078 856
rect 232246 31 233826 856
rect 233994 31 235574 856
rect 235742 31 237322 856
rect 237490 31 239070 856
rect 239238 31 240818 856
rect 240986 31 242566 856
rect 242734 31 244314 856
rect 244482 31 246062 856
rect 246230 31 247810 856
rect 247978 31 249558 856
rect 249726 31 251306 856
rect 251474 31 253054 856
rect 253222 31 254802 856
rect 254970 31 256550 856
rect 256718 31 258298 856
rect 258466 31 260046 856
rect 260214 31 261794 856
rect 261962 31 263542 856
rect 263710 31 265290 856
rect 265458 31 267038 856
rect 267206 31 268786 856
rect 268954 31 270534 856
rect 270702 31 272282 856
rect 272450 31 274030 856
rect 274198 31 275778 856
rect 275946 31 277526 856
rect 277694 31 279274 856
rect 279442 31 281022 856
rect 281190 31 282770 856
rect 282938 31 284518 856
rect 284686 31 286266 856
rect 286434 31 288014 856
rect 288182 31 289762 856
rect 289930 31 291510 856
rect 291678 31 293258 856
rect 293426 31 295006 856
rect 295174 31 296754 856
rect 296922 31 298502 856
rect 298670 31 300250 856
rect 300418 31 301998 856
rect 302166 31 303746 856
rect 303914 31 305494 856
rect 305662 31 307242 856
rect 307410 31 308990 856
rect 309158 31 310738 856
rect 310906 31 312486 856
rect 312654 31 314234 856
rect 314402 31 315982 856
rect 316150 31 317730 856
rect 317898 31 319478 856
rect 319646 31 321226 856
rect 321394 31 322974 856
rect 323142 31 324722 856
rect 324890 31 326470 856
rect 326638 31 328218 856
rect 328386 31 329966 856
rect 330134 31 331714 856
rect 331882 31 333462 856
rect 333630 31 335210 856
rect 335378 31 336958 856
rect 337126 31 338706 856
rect 338874 31 340454 856
rect 340622 31 342202 856
rect 342370 31 343950 856
rect 344118 31 345698 856
rect 345866 31 347446 856
rect 347614 31 349194 856
rect 349362 31 350942 856
rect 351110 31 352690 856
rect 352858 31 354438 856
rect 354606 31 356186 856
rect 356354 31 357934 856
rect 358102 31 359682 856
rect 359850 31 361430 856
rect 361598 31 363178 856
rect 363346 31 364926 856
rect 365094 31 366674 856
rect 366842 31 368422 856
rect 368590 31 370170 856
rect 370338 31 371918 856
rect 372086 31 373666 856
rect 373834 31 375414 856
rect 375582 31 377162 856
rect 377330 31 378910 856
rect 379078 31 380658 856
rect 380826 31 382406 856
rect 382574 31 384154 856
rect 384322 31 385902 856
rect 386070 31 387650 856
rect 387818 31 389398 856
rect 389566 31 391146 856
rect 391314 31 392894 856
rect 393062 31 394642 856
rect 394810 31 396390 856
rect 396558 31 398138 856
rect 398306 31 399886 856
rect 400054 31 401634 856
rect 401802 31 403382 856
rect 403550 31 405130 856
rect 405298 31 406878 856
rect 407046 31 408626 856
rect 408794 31 410374 856
rect 410542 31 412122 856
rect 412290 31 413870 856
rect 414038 31 415618 856
rect 415786 31 417366 856
rect 417534 31 419114 856
rect 419282 31 420862 856
rect 421030 31 422610 856
rect 422778 31 424358 856
rect 424526 31 426106 856
rect 426274 31 427854 856
rect 428022 31 429602 856
rect 429770 31 431350 856
rect 431518 31 439372 856
<< metal3 >>
rect 439200 150968 440000 151088
rect 439200 150424 440000 150544
rect 0 149880 800 150000
rect 439200 149880 440000 150000
rect 0 149336 800 149456
rect 439200 149336 440000 149456
rect 0 148792 800 148912
rect 439200 148792 440000 148912
rect 0 148248 800 148368
rect 439200 148248 440000 148368
rect 0 147704 800 147824
rect 439200 147704 440000 147824
rect 0 147160 800 147280
rect 439200 147160 440000 147280
rect 0 146616 800 146736
rect 439200 146616 440000 146736
rect 0 146072 800 146192
rect 439200 146072 440000 146192
rect 0 145528 800 145648
rect 439200 145528 440000 145648
rect 0 144984 800 145104
rect 439200 144984 440000 145104
rect 0 144440 800 144560
rect 439200 144440 440000 144560
rect 0 143896 800 144016
rect 439200 143896 440000 144016
rect 0 143352 800 143472
rect 439200 143352 440000 143472
rect 0 142808 800 142928
rect 439200 142808 440000 142928
rect 0 142264 800 142384
rect 439200 142264 440000 142384
rect 0 141720 800 141840
rect 439200 141720 440000 141840
rect 0 141176 800 141296
rect 439200 141176 440000 141296
rect 0 140632 800 140752
rect 439200 140632 440000 140752
rect 0 140088 800 140208
rect 439200 140088 440000 140208
rect 0 139544 800 139664
rect 439200 139544 440000 139664
rect 0 139000 800 139120
rect 439200 139000 440000 139120
rect 0 138456 800 138576
rect 439200 138456 440000 138576
rect 0 137912 800 138032
rect 439200 137912 440000 138032
rect 0 137368 800 137488
rect 439200 137368 440000 137488
rect 0 136824 800 136944
rect 439200 136824 440000 136944
rect 0 136280 800 136400
rect 439200 136280 440000 136400
rect 0 135736 800 135856
rect 439200 135736 440000 135856
rect 0 135192 800 135312
rect 439200 135192 440000 135312
rect 0 134648 800 134768
rect 439200 134648 440000 134768
rect 0 134104 800 134224
rect 439200 134104 440000 134224
rect 0 133560 800 133680
rect 439200 133560 440000 133680
rect 0 133016 800 133136
rect 439200 133016 440000 133136
rect 0 132472 800 132592
rect 439200 132472 440000 132592
rect 0 131928 800 132048
rect 439200 131928 440000 132048
rect 0 131384 800 131504
rect 439200 131384 440000 131504
rect 0 130840 800 130960
rect 439200 130840 440000 130960
rect 0 130296 800 130416
rect 439200 130296 440000 130416
rect 0 129752 800 129872
rect 439200 129752 440000 129872
rect 0 129208 800 129328
rect 439200 129208 440000 129328
rect 0 128664 800 128784
rect 439200 128664 440000 128784
rect 0 128120 800 128240
rect 439200 128120 440000 128240
rect 0 127576 800 127696
rect 439200 127576 440000 127696
rect 0 127032 800 127152
rect 439200 127032 440000 127152
rect 0 126488 800 126608
rect 439200 126488 440000 126608
rect 0 125944 800 126064
rect 439200 125944 440000 126064
rect 0 125400 800 125520
rect 439200 125400 440000 125520
rect 0 124856 800 124976
rect 439200 124856 440000 124976
rect 0 124312 800 124432
rect 439200 124312 440000 124432
rect 0 123768 800 123888
rect 439200 123768 440000 123888
rect 0 123224 800 123344
rect 439200 123224 440000 123344
rect 0 122680 800 122800
rect 439200 122680 440000 122800
rect 0 122136 800 122256
rect 439200 122136 440000 122256
rect 0 121592 800 121712
rect 439200 121592 440000 121712
rect 0 121048 800 121168
rect 439200 121048 440000 121168
rect 0 120504 800 120624
rect 439200 120504 440000 120624
rect 0 119960 800 120080
rect 439200 119960 440000 120080
rect 0 119416 800 119536
rect 439200 119416 440000 119536
rect 0 118872 800 118992
rect 439200 118872 440000 118992
rect 0 118328 800 118448
rect 439200 118328 440000 118448
rect 0 117784 800 117904
rect 439200 117784 440000 117904
rect 0 117240 800 117360
rect 439200 117240 440000 117360
rect 0 116696 800 116816
rect 439200 116696 440000 116816
rect 0 116152 800 116272
rect 439200 116152 440000 116272
rect 0 115608 800 115728
rect 439200 115608 440000 115728
rect 0 115064 800 115184
rect 439200 115064 440000 115184
rect 0 114520 800 114640
rect 439200 114520 440000 114640
rect 0 113976 800 114096
rect 439200 113976 440000 114096
rect 0 113432 800 113552
rect 439200 113432 440000 113552
rect 0 112888 800 113008
rect 439200 112888 440000 113008
rect 0 112344 800 112464
rect 439200 112344 440000 112464
rect 0 111800 800 111920
rect 439200 111800 440000 111920
rect 0 111256 800 111376
rect 439200 111256 440000 111376
rect 0 110712 800 110832
rect 439200 110712 440000 110832
rect 0 110168 800 110288
rect 439200 110168 440000 110288
rect 0 109624 800 109744
rect 439200 109624 440000 109744
rect 0 109080 800 109200
rect 439200 109080 440000 109200
rect 0 108536 800 108656
rect 439200 108536 440000 108656
rect 0 107992 800 108112
rect 439200 107992 440000 108112
rect 0 107448 800 107568
rect 439200 107448 440000 107568
rect 0 106904 800 107024
rect 439200 106904 440000 107024
rect 0 106360 800 106480
rect 439200 106360 440000 106480
rect 0 105816 800 105936
rect 439200 105816 440000 105936
rect 0 105272 800 105392
rect 439200 105272 440000 105392
rect 0 104728 800 104848
rect 439200 104728 440000 104848
rect 0 104184 800 104304
rect 439200 104184 440000 104304
rect 0 103640 800 103760
rect 439200 103640 440000 103760
rect 0 103096 800 103216
rect 439200 103096 440000 103216
rect 0 102552 800 102672
rect 439200 102552 440000 102672
rect 0 102008 800 102128
rect 439200 102008 440000 102128
rect 0 101464 800 101584
rect 439200 101464 440000 101584
rect 0 100920 800 101040
rect 439200 100920 440000 101040
rect 0 100376 800 100496
rect 439200 100376 440000 100496
rect 0 99832 800 99952
rect 439200 99832 440000 99952
rect 0 99288 800 99408
rect 439200 99288 440000 99408
rect 0 98744 800 98864
rect 439200 98744 440000 98864
rect 0 98200 800 98320
rect 439200 98200 440000 98320
rect 0 97656 800 97776
rect 439200 97656 440000 97776
rect 0 97112 800 97232
rect 439200 97112 440000 97232
rect 0 96568 800 96688
rect 439200 96568 440000 96688
rect 0 96024 800 96144
rect 439200 96024 440000 96144
rect 0 95480 800 95600
rect 439200 95480 440000 95600
rect 0 94936 800 95056
rect 439200 94936 440000 95056
rect 0 94392 800 94512
rect 439200 94392 440000 94512
rect 0 93848 800 93968
rect 439200 93848 440000 93968
rect 0 93304 800 93424
rect 439200 93304 440000 93424
rect 0 92760 800 92880
rect 439200 92760 440000 92880
rect 0 92216 800 92336
rect 439200 92216 440000 92336
rect 0 91672 800 91792
rect 439200 91672 440000 91792
rect 0 91128 800 91248
rect 439200 91128 440000 91248
rect 0 90584 800 90704
rect 439200 90584 440000 90704
rect 0 90040 800 90160
rect 439200 90040 440000 90160
rect 0 89496 800 89616
rect 439200 89496 440000 89616
rect 0 88952 800 89072
rect 439200 88952 440000 89072
rect 0 88408 800 88528
rect 439200 88408 440000 88528
rect 0 87864 800 87984
rect 439200 87864 440000 87984
rect 0 87320 800 87440
rect 439200 87320 440000 87440
rect 0 86776 800 86896
rect 439200 86776 440000 86896
rect 0 86232 800 86352
rect 439200 86232 440000 86352
rect 0 85688 800 85808
rect 439200 85688 440000 85808
rect 0 85144 800 85264
rect 439200 85144 440000 85264
rect 0 84600 800 84720
rect 439200 84600 440000 84720
rect 0 84056 800 84176
rect 439200 84056 440000 84176
rect 0 83512 800 83632
rect 439200 83512 440000 83632
rect 0 82968 800 83088
rect 439200 82968 440000 83088
rect 0 82424 800 82544
rect 439200 82424 440000 82544
rect 0 81880 800 82000
rect 439200 81880 440000 82000
rect 0 81336 800 81456
rect 439200 81336 440000 81456
rect 0 80792 800 80912
rect 439200 80792 440000 80912
rect 0 80248 800 80368
rect 439200 80248 440000 80368
rect 0 79704 800 79824
rect 439200 79704 440000 79824
rect 0 79160 800 79280
rect 439200 79160 440000 79280
rect 0 78616 800 78736
rect 439200 78616 440000 78736
rect 0 78072 800 78192
rect 439200 78072 440000 78192
rect 0 77528 800 77648
rect 439200 77528 440000 77648
rect 0 76984 800 77104
rect 439200 76984 440000 77104
rect 0 76440 800 76560
rect 439200 76440 440000 76560
rect 0 75896 800 76016
rect 439200 75896 440000 76016
rect 0 75352 800 75472
rect 439200 75352 440000 75472
rect 0 74808 800 74928
rect 439200 74808 440000 74928
rect 0 74264 800 74384
rect 439200 74264 440000 74384
rect 0 73720 800 73840
rect 439200 73720 440000 73840
rect 0 73176 800 73296
rect 439200 73176 440000 73296
rect 0 72632 800 72752
rect 439200 72632 440000 72752
rect 0 72088 800 72208
rect 439200 72088 440000 72208
rect 0 71544 800 71664
rect 439200 71544 440000 71664
rect 0 71000 800 71120
rect 439200 71000 440000 71120
rect 0 70456 800 70576
rect 439200 70456 440000 70576
rect 0 69912 800 70032
rect 439200 69912 440000 70032
rect 0 69368 800 69488
rect 439200 69368 440000 69488
rect 0 68824 800 68944
rect 439200 68824 440000 68944
rect 0 68280 800 68400
rect 439200 68280 440000 68400
rect 0 67736 800 67856
rect 439200 67736 440000 67856
rect 0 67192 800 67312
rect 439200 67192 440000 67312
rect 0 66648 800 66768
rect 439200 66648 440000 66768
rect 0 66104 800 66224
rect 439200 66104 440000 66224
rect 0 65560 800 65680
rect 439200 65560 440000 65680
rect 0 65016 800 65136
rect 439200 65016 440000 65136
rect 0 64472 800 64592
rect 439200 64472 440000 64592
rect 0 63928 800 64048
rect 439200 63928 440000 64048
rect 0 63384 800 63504
rect 439200 63384 440000 63504
rect 0 62840 800 62960
rect 439200 62840 440000 62960
rect 0 62296 800 62416
rect 439200 62296 440000 62416
rect 0 61752 800 61872
rect 439200 61752 440000 61872
rect 0 61208 800 61328
rect 439200 61208 440000 61328
rect 0 60664 800 60784
rect 439200 60664 440000 60784
rect 0 60120 800 60240
rect 439200 60120 440000 60240
rect 0 59576 800 59696
rect 439200 59576 440000 59696
rect 0 59032 800 59152
rect 439200 59032 440000 59152
rect 0 58488 800 58608
rect 439200 58488 440000 58608
rect 0 57944 800 58064
rect 439200 57944 440000 58064
rect 0 57400 800 57520
rect 439200 57400 440000 57520
rect 0 56856 800 56976
rect 439200 56856 440000 56976
rect 0 56312 800 56432
rect 439200 56312 440000 56432
rect 0 55768 800 55888
rect 439200 55768 440000 55888
rect 0 55224 800 55344
rect 439200 55224 440000 55344
rect 0 54680 800 54800
rect 439200 54680 440000 54800
rect 0 54136 800 54256
rect 439200 54136 440000 54256
rect 0 53592 800 53712
rect 439200 53592 440000 53712
rect 0 53048 800 53168
rect 439200 53048 440000 53168
rect 0 52504 800 52624
rect 439200 52504 440000 52624
rect 0 51960 800 52080
rect 439200 51960 440000 52080
rect 0 51416 800 51536
rect 439200 51416 440000 51536
rect 0 50872 800 50992
rect 439200 50872 440000 50992
rect 0 50328 800 50448
rect 439200 50328 440000 50448
rect 0 49784 800 49904
rect 439200 49784 440000 49904
rect 0 49240 800 49360
rect 439200 49240 440000 49360
rect 0 48696 800 48816
rect 439200 48696 440000 48816
rect 0 48152 800 48272
rect 439200 48152 440000 48272
rect 0 47608 800 47728
rect 439200 47608 440000 47728
rect 0 47064 800 47184
rect 439200 47064 440000 47184
rect 0 46520 800 46640
rect 439200 46520 440000 46640
rect 0 45976 800 46096
rect 439200 45976 440000 46096
rect 0 45432 800 45552
rect 439200 45432 440000 45552
rect 0 44888 800 45008
rect 439200 44888 440000 45008
rect 0 44344 800 44464
rect 439200 44344 440000 44464
rect 0 43800 800 43920
rect 439200 43800 440000 43920
rect 0 43256 800 43376
rect 439200 43256 440000 43376
rect 0 42712 800 42832
rect 439200 42712 440000 42832
rect 0 42168 800 42288
rect 439200 42168 440000 42288
rect 0 41624 800 41744
rect 439200 41624 440000 41744
rect 0 41080 800 41200
rect 439200 41080 440000 41200
rect 0 40536 800 40656
rect 439200 40536 440000 40656
rect 0 39992 800 40112
rect 439200 39992 440000 40112
rect 0 39448 800 39568
rect 439200 39448 440000 39568
rect 0 38904 800 39024
rect 439200 38904 440000 39024
rect 0 38360 800 38480
rect 439200 38360 440000 38480
rect 0 37816 800 37936
rect 439200 37816 440000 37936
rect 0 37272 800 37392
rect 439200 37272 440000 37392
rect 0 36728 800 36848
rect 439200 36728 440000 36848
rect 0 36184 800 36304
rect 439200 36184 440000 36304
rect 0 35640 800 35760
rect 439200 35640 440000 35760
rect 0 35096 800 35216
rect 439200 35096 440000 35216
rect 0 34552 800 34672
rect 439200 34552 440000 34672
rect 0 34008 800 34128
rect 439200 34008 440000 34128
rect 0 33464 800 33584
rect 439200 33464 440000 33584
rect 0 32920 800 33040
rect 439200 32920 440000 33040
rect 0 32376 800 32496
rect 439200 32376 440000 32496
rect 0 31832 800 31952
rect 439200 31832 440000 31952
rect 0 31288 800 31408
rect 439200 31288 440000 31408
rect 0 30744 800 30864
rect 439200 30744 440000 30864
rect 0 30200 800 30320
rect 439200 30200 440000 30320
rect 0 29656 800 29776
rect 439200 29656 440000 29776
rect 0 29112 800 29232
rect 439200 29112 440000 29232
rect 0 28568 800 28688
rect 439200 28568 440000 28688
rect 0 28024 800 28144
rect 439200 28024 440000 28144
rect 0 27480 800 27600
rect 439200 27480 440000 27600
rect 0 26936 800 27056
rect 439200 26936 440000 27056
rect 0 26392 800 26512
rect 439200 26392 440000 26512
rect 0 25848 800 25968
rect 439200 25848 440000 25968
rect 0 25304 800 25424
rect 439200 25304 440000 25424
rect 0 24760 800 24880
rect 439200 24760 440000 24880
rect 0 24216 800 24336
rect 439200 24216 440000 24336
rect 0 23672 800 23792
rect 439200 23672 440000 23792
rect 0 23128 800 23248
rect 439200 23128 440000 23248
rect 0 22584 800 22704
rect 439200 22584 440000 22704
rect 0 22040 800 22160
rect 439200 22040 440000 22160
rect 0 21496 800 21616
rect 439200 21496 440000 21616
rect 0 20952 800 21072
rect 439200 20952 440000 21072
rect 0 20408 800 20528
rect 439200 20408 440000 20528
rect 0 19864 800 19984
rect 439200 19864 440000 19984
rect 439200 19320 440000 19440
rect 439200 18776 440000 18896
<< obsm3 >>
rect 800 151168 439200 169285
rect 800 150888 439120 151168
rect 800 150624 439200 150888
rect 800 150344 439120 150624
rect 800 150080 439200 150344
rect 880 149800 439120 150080
rect 800 149536 439200 149800
rect 880 149256 439120 149536
rect 800 148992 439200 149256
rect 880 148712 439120 148992
rect 800 148448 439200 148712
rect 880 148168 439120 148448
rect 800 147904 439200 148168
rect 880 147624 439120 147904
rect 800 147360 439200 147624
rect 880 147080 439120 147360
rect 800 146816 439200 147080
rect 880 146536 439120 146816
rect 800 146272 439200 146536
rect 880 145992 439120 146272
rect 800 145728 439200 145992
rect 880 145448 439120 145728
rect 800 145184 439200 145448
rect 880 144904 439120 145184
rect 800 144640 439200 144904
rect 880 144360 439120 144640
rect 800 144096 439200 144360
rect 880 143816 439120 144096
rect 800 143552 439200 143816
rect 880 143272 439120 143552
rect 800 143008 439200 143272
rect 880 142728 439120 143008
rect 800 142464 439200 142728
rect 880 142184 439120 142464
rect 800 141920 439200 142184
rect 880 141640 439120 141920
rect 800 141376 439200 141640
rect 880 141096 439120 141376
rect 800 140832 439200 141096
rect 880 140552 439120 140832
rect 800 140288 439200 140552
rect 880 140008 439120 140288
rect 800 139744 439200 140008
rect 880 139464 439120 139744
rect 800 139200 439200 139464
rect 880 138920 439120 139200
rect 800 138656 439200 138920
rect 880 138376 439120 138656
rect 800 138112 439200 138376
rect 880 137832 439120 138112
rect 800 137568 439200 137832
rect 880 137288 439120 137568
rect 800 137024 439200 137288
rect 880 136744 439120 137024
rect 800 136480 439200 136744
rect 880 136200 439120 136480
rect 800 135936 439200 136200
rect 880 135656 439120 135936
rect 800 135392 439200 135656
rect 880 135112 439120 135392
rect 800 134848 439200 135112
rect 880 134568 439120 134848
rect 800 134304 439200 134568
rect 880 134024 439120 134304
rect 800 133760 439200 134024
rect 880 133480 439120 133760
rect 800 133216 439200 133480
rect 880 132936 439120 133216
rect 800 132672 439200 132936
rect 880 132392 439120 132672
rect 800 132128 439200 132392
rect 880 131848 439120 132128
rect 800 131584 439200 131848
rect 880 131304 439120 131584
rect 800 131040 439200 131304
rect 880 130760 439120 131040
rect 800 130496 439200 130760
rect 880 130216 439120 130496
rect 800 129952 439200 130216
rect 880 129672 439120 129952
rect 800 129408 439200 129672
rect 880 129128 439120 129408
rect 800 128864 439200 129128
rect 880 128584 439120 128864
rect 800 128320 439200 128584
rect 880 128040 439120 128320
rect 800 127776 439200 128040
rect 880 127496 439120 127776
rect 800 127232 439200 127496
rect 880 126952 439120 127232
rect 800 126688 439200 126952
rect 880 126408 439120 126688
rect 800 126144 439200 126408
rect 880 125864 439120 126144
rect 800 125600 439200 125864
rect 880 125320 439120 125600
rect 800 125056 439200 125320
rect 880 124776 439120 125056
rect 800 124512 439200 124776
rect 880 124232 439120 124512
rect 800 123968 439200 124232
rect 880 123688 439120 123968
rect 800 123424 439200 123688
rect 880 123144 439120 123424
rect 800 122880 439200 123144
rect 880 122600 439120 122880
rect 800 122336 439200 122600
rect 880 122056 439120 122336
rect 800 121792 439200 122056
rect 880 121512 439120 121792
rect 800 121248 439200 121512
rect 880 120968 439120 121248
rect 800 120704 439200 120968
rect 880 120424 439120 120704
rect 800 120160 439200 120424
rect 880 119880 439120 120160
rect 800 119616 439200 119880
rect 880 119336 439120 119616
rect 800 119072 439200 119336
rect 880 118792 439120 119072
rect 800 118528 439200 118792
rect 880 118248 439120 118528
rect 800 117984 439200 118248
rect 880 117704 439120 117984
rect 800 117440 439200 117704
rect 880 117160 439120 117440
rect 800 116896 439200 117160
rect 880 116616 439120 116896
rect 800 116352 439200 116616
rect 880 116072 439120 116352
rect 800 115808 439200 116072
rect 880 115528 439120 115808
rect 800 115264 439200 115528
rect 880 114984 439120 115264
rect 800 114720 439200 114984
rect 880 114440 439120 114720
rect 800 114176 439200 114440
rect 880 113896 439120 114176
rect 800 113632 439200 113896
rect 880 113352 439120 113632
rect 800 113088 439200 113352
rect 880 112808 439120 113088
rect 800 112544 439200 112808
rect 880 112264 439120 112544
rect 800 112000 439200 112264
rect 880 111720 439120 112000
rect 800 111456 439200 111720
rect 880 111176 439120 111456
rect 800 110912 439200 111176
rect 880 110632 439120 110912
rect 800 110368 439200 110632
rect 880 110088 439120 110368
rect 800 109824 439200 110088
rect 880 109544 439120 109824
rect 800 109280 439200 109544
rect 880 109000 439120 109280
rect 800 108736 439200 109000
rect 880 108456 439120 108736
rect 800 108192 439200 108456
rect 880 107912 439120 108192
rect 800 107648 439200 107912
rect 880 107368 439120 107648
rect 800 107104 439200 107368
rect 880 106824 439120 107104
rect 800 106560 439200 106824
rect 880 106280 439120 106560
rect 800 106016 439200 106280
rect 880 105736 439120 106016
rect 800 105472 439200 105736
rect 880 105192 439120 105472
rect 800 104928 439200 105192
rect 880 104648 439120 104928
rect 800 104384 439200 104648
rect 880 104104 439120 104384
rect 800 103840 439200 104104
rect 880 103560 439120 103840
rect 800 103296 439200 103560
rect 880 103016 439120 103296
rect 800 102752 439200 103016
rect 880 102472 439120 102752
rect 800 102208 439200 102472
rect 880 101928 439120 102208
rect 800 101664 439200 101928
rect 880 101384 439120 101664
rect 800 101120 439200 101384
rect 880 100840 439120 101120
rect 800 100576 439200 100840
rect 880 100296 439120 100576
rect 800 100032 439200 100296
rect 880 99752 439120 100032
rect 800 99488 439200 99752
rect 880 99208 439120 99488
rect 800 98944 439200 99208
rect 880 98664 439120 98944
rect 800 98400 439200 98664
rect 880 98120 439120 98400
rect 800 97856 439200 98120
rect 880 97576 439120 97856
rect 800 97312 439200 97576
rect 880 97032 439120 97312
rect 800 96768 439200 97032
rect 880 96488 439120 96768
rect 800 96224 439200 96488
rect 880 95944 439120 96224
rect 800 95680 439200 95944
rect 880 95400 439120 95680
rect 800 95136 439200 95400
rect 880 94856 439120 95136
rect 800 94592 439200 94856
rect 880 94312 439120 94592
rect 800 94048 439200 94312
rect 880 93768 439120 94048
rect 800 93504 439200 93768
rect 880 93224 439120 93504
rect 800 92960 439200 93224
rect 880 92680 439120 92960
rect 800 92416 439200 92680
rect 880 92136 439120 92416
rect 800 91872 439200 92136
rect 880 91592 439120 91872
rect 800 91328 439200 91592
rect 880 91048 439120 91328
rect 800 90784 439200 91048
rect 880 90504 439120 90784
rect 800 90240 439200 90504
rect 880 89960 439120 90240
rect 800 89696 439200 89960
rect 880 89416 439120 89696
rect 800 89152 439200 89416
rect 880 88872 439120 89152
rect 800 88608 439200 88872
rect 880 88328 439120 88608
rect 800 88064 439200 88328
rect 880 87784 439120 88064
rect 800 87520 439200 87784
rect 880 87240 439120 87520
rect 800 86976 439200 87240
rect 880 86696 439120 86976
rect 800 86432 439200 86696
rect 880 86152 439120 86432
rect 800 85888 439200 86152
rect 880 85608 439120 85888
rect 800 85344 439200 85608
rect 880 85064 439120 85344
rect 800 84800 439200 85064
rect 880 84520 439120 84800
rect 800 84256 439200 84520
rect 880 83976 439120 84256
rect 800 83712 439200 83976
rect 880 83432 439120 83712
rect 800 83168 439200 83432
rect 880 82888 439120 83168
rect 800 82624 439200 82888
rect 880 82344 439120 82624
rect 800 82080 439200 82344
rect 880 81800 439120 82080
rect 800 81536 439200 81800
rect 880 81256 439120 81536
rect 800 80992 439200 81256
rect 880 80712 439120 80992
rect 800 80448 439200 80712
rect 880 80168 439120 80448
rect 800 79904 439200 80168
rect 880 79624 439120 79904
rect 800 79360 439200 79624
rect 880 79080 439120 79360
rect 800 78816 439200 79080
rect 880 78536 439120 78816
rect 800 78272 439200 78536
rect 880 77992 439120 78272
rect 800 77728 439200 77992
rect 880 77448 439120 77728
rect 800 77184 439200 77448
rect 880 76904 439120 77184
rect 800 76640 439200 76904
rect 880 76360 439120 76640
rect 800 76096 439200 76360
rect 880 75816 439120 76096
rect 800 75552 439200 75816
rect 880 75272 439120 75552
rect 800 75008 439200 75272
rect 880 74728 439120 75008
rect 800 74464 439200 74728
rect 880 74184 439120 74464
rect 800 73920 439200 74184
rect 880 73640 439120 73920
rect 800 73376 439200 73640
rect 880 73096 439120 73376
rect 800 72832 439200 73096
rect 880 72552 439120 72832
rect 800 72288 439200 72552
rect 880 72008 439120 72288
rect 800 71744 439200 72008
rect 880 71464 439120 71744
rect 800 71200 439200 71464
rect 880 70920 439120 71200
rect 800 70656 439200 70920
rect 880 70376 439120 70656
rect 800 70112 439200 70376
rect 880 69832 439120 70112
rect 800 69568 439200 69832
rect 880 69288 439120 69568
rect 800 69024 439200 69288
rect 880 68744 439120 69024
rect 800 68480 439200 68744
rect 880 68200 439120 68480
rect 800 67936 439200 68200
rect 880 67656 439120 67936
rect 800 67392 439200 67656
rect 880 67112 439120 67392
rect 800 66848 439200 67112
rect 880 66568 439120 66848
rect 800 66304 439200 66568
rect 880 66024 439120 66304
rect 800 65760 439200 66024
rect 880 65480 439120 65760
rect 800 65216 439200 65480
rect 880 64936 439120 65216
rect 800 64672 439200 64936
rect 880 64392 439120 64672
rect 800 64128 439200 64392
rect 880 63848 439120 64128
rect 800 63584 439200 63848
rect 880 63304 439120 63584
rect 800 63040 439200 63304
rect 880 62760 439120 63040
rect 800 62496 439200 62760
rect 880 62216 439120 62496
rect 800 61952 439200 62216
rect 880 61672 439120 61952
rect 800 61408 439200 61672
rect 880 61128 439120 61408
rect 800 60864 439200 61128
rect 880 60584 439120 60864
rect 800 60320 439200 60584
rect 880 60040 439120 60320
rect 800 59776 439200 60040
rect 880 59496 439120 59776
rect 800 59232 439200 59496
rect 880 58952 439120 59232
rect 800 58688 439200 58952
rect 880 58408 439120 58688
rect 800 58144 439200 58408
rect 880 57864 439120 58144
rect 800 57600 439200 57864
rect 880 57320 439120 57600
rect 800 57056 439200 57320
rect 880 56776 439120 57056
rect 800 56512 439200 56776
rect 880 56232 439120 56512
rect 800 55968 439200 56232
rect 880 55688 439120 55968
rect 800 55424 439200 55688
rect 880 55144 439120 55424
rect 800 54880 439200 55144
rect 880 54600 439120 54880
rect 800 54336 439200 54600
rect 880 54056 439120 54336
rect 800 53792 439200 54056
rect 880 53512 439120 53792
rect 800 53248 439200 53512
rect 880 52968 439120 53248
rect 800 52704 439200 52968
rect 880 52424 439120 52704
rect 800 52160 439200 52424
rect 880 51880 439120 52160
rect 800 51616 439200 51880
rect 880 51336 439120 51616
rect 800 51072 439200 51336
rect 880 50792 439120 51072
rect 800 50528 439200 50792
rect 880 50248 439120 50528
rect 800 49984 439200 50248
rect 880 49704 439120 49984
rect 800 49440 439200 49704
rect 880 49160 439120 49440
rect 800 48896 439200 49160
rect 880 48616 439120 48896
rect 800 48352 439200 48616
rect 880 48072 439120 48352
rect 800 47808 439200 48072
rect 880 47528 439120 47808
rect 800 47264 439200 47528
rect 880 46984 439120 47264
rect 800 46720 439200 46984
rect 880 46440 439120 46720
rect 800 46176 439200 46440
rect 880 45896 439120 46176
rect 800 45632 439200 45896
rect 880 45352 439120 45632
rect 800 45088 439200 45352
rect 880 44808 439120 45088
rect 800 44544 439200 44808
rect 880 44264 439120 44544
rect 800 44000 439200 44264
rect 880 43720 439120 44000
rect 800 43456 439200 43720
rect 880 43176 439120 43456
rect 800 42912 439200 43176
rect 880 42632 439120 42912
rect 800 42368 439200 42632
rect 880 42088 439120 42368
rect 800 41824 439200 42088
rect 880 41544 439120 41824
rect 800 41280 439200 41544
rect 880 41000 439120 41280
rect 800 40736 439200 41000
rect 880 40456 439120 40736
rect 800 40192 439200 40456
rect 880 39912 439120 40192
rect 800 39648 439200 39912
rect 880 39368 439120 39648
rect 800 39104 439200 39368
rect 880 38824 439120 39104
rect 800 38560 439200 38824
rect 880 38280 439120 38560
rect 800 38016 439200 38280
rect 880 37736 439120 38016
rect 800 37472 439200 37736
rect 880 37192 439120 37472
rect 800 36928 439200 37192
rect 880 36648 439120 36928
rect 800 36384 439200 36648
rect 880 36104 439120 36384
rect 800 35840 439200 36104
rect 880 35560 439120 35840
rect 800 35296 439200 35560
rect 880 35016 439120 35296
rect 800 34752 439200 35016
rect 880 34472 439120 34752
rect 800 34208 439200 34472
rect 880 33928 439120 34208
rect 800 33664 439200 33928
rect 880 33384 439120 33664
rect 800 33120 439200 33384
rect 880 32840 439120 33120
rect 800 32576 439200 32840
rect 880 32296 439120 32576
rect 800 32032 439200 32296
rect 880 31752 439120 32032
rect 800 31488 439200 31752
rect 880 31208 439120 31488
rect 800 30944 439200 31208
rect 880 30664 439120 30944
rect 800 30400 439200 30664
rect 880 30120 439120 30400
rect 800 29856 439200 30120
rect 880 29576 439120 29856
rect 800 29312 439200 29576
rect 880 29032 439120 29312
rect 800 28768 439200 29032
rect 880 28488 439120 28768
rect 800 28224 439200 28488
rect 880 27944 439120 28224
rect 800 27680 439200 27944
rect 880 27400 439120 27680
rect 800 27136 439200 27400
rect 880 26856 439120 27136
rect 800 26592 439200 26856
rect 880 26312 439120 26592
rect 800 26048 439200 26312
rect 880 25768 439120 26048
rect 800 25504 439200 25768
rect 880 25224 439120 25504
rect 800 24960 439200 25224
rect 880 24680 439120 24960
rect 800 24416 439200 24680
rect 880 24136 439120 24416
rect 800 23872 439200 24136
rect 880 23592 439120 23872
rect 800 23328 439200 23592
rect 880 23048 439120 23328
rect 800 22784 439200 23048
rect 880 22504 439120 22784
rect 800 22240 439200 22504
rect 880 21960 439120 22240
rect 800 21696 439200 21960
rect 880 21416 439120 21696
rect 800 21152 439200 21416
rect 880 20872 439120 21152
rect 800 20608 439200 20872
rect 880 20328 439120 20608
rect 800 20064 439200 20328
rect 880 19784 439120 20064
rect 800 19520 439200 19784
rect 800 19240 439120 19520
rect 800 18976 439200 19240
rect 800 18696 439120 18976
rect 800 35 439200 18696
<< metal4 >>
rect 4208 2128 4528 167600
rect 19568 2128 19888 167600
rect 34928 2128 35248 167600
rect 50288 2128 50608 167600
rect 65648 2128 65968 167600
rect 81008 2128 81328 167600
rect 96368 2128 96688 167600
rect 111728 2128 112048 167600
rect 127088 2128 127408 167600
rect 142448 2128 142768 167600
rect 157808 2128 158128 167600
rect 173168 2128 173488 167600
rect 188528 2128 188848 167600
rect 203888 2128 204208 167600
rect 219248 2128 219568 167600
rect 234608 2128 234928 167600
rect 249968 2128 250288 167600
rect 265328 2128 265648 167600
rect 280688 2128 281008 167600
rect 296048 2128 296368 167600
rect 311408 2128 311728 167600
rect 326768 2128 327088 167600
rect 342128 2128 342448 167600
rect 357488 2128 357808 167600
rect 372848 2128 373168 167600
rect 388208 2128 388528 167600
rect 403568 2128 403888 167600
rect 418928 2128 419248 167600
rect 434288 2128 434608 167600
<< obsm4 >>
rect 3371 167680 436941 169149
rect 3371 2048 4128 167680
rect 4608 2048 19488 167680
rect 19968 2048 34848 167680
rect 35328 2048 50208 167680
rect 50688 2048 65568 167680
rect 66048 2048 80928 167680
rect 81408 2048 96288 167680
rect 96768 2048 111648 167680
rect 112128 2048 127008 167680
rect 127488 2048 142368 167680
rect 142848 2048 157728 167680
rect 158208 2048 173088 167680
rect 173568 2048 188448 167680
rect 188928 2048 203808 167680
rect 204288 2048 219168 167680
rect 219648 2048 234528 167680
rect 235008 2048 249888 167680
rect 250368 2048 265248 167680
rect 265728 2048 280608 167680
rect 281088 2048 295968 167680
rect 296448 2048 311328 167680
rect 311808 2048 326688 167680
rect 327168 2048 342048 167680
rect 342528 2048 357408 167680
rect 357888 2048 372768 167680
rect 373248 2048 388128 167680
rect 388608 2048 403488 167680
rect 403968 2048 418848 167680
rect 419328 2048 434208 167680
rect 434688 2048 436941 167680
rect 3371 35 436941 2048
<< labels >>
rlabel metal2 s 5354 169200 5410 170000 6 cache_PC[0]
port 1 nsew signal output
rlabel metal2 s 15474 169200 15530 170000 6 cache_PC[10]
port 2 nsew signal output
rlabel metal2 s 16486 169200 16542 170000 6 cache_PC[11]
port 3 nsew signal output
rlabel metal2 s 17498 169200 17554 170000 6 cache_PC[12]
port 4 nsew signal output
rlabel metal2 s 18510 169200 18566 170000 6 cache_PC[13]
port 5 nsew signal output
rlabel metal2 s 19522 169200 19578 170000 6 cache_PC[14]
port 6 nsew signal output
rlabel metal2 s 20534 169200 20590 170000 6 cache_PC[15]
port 7 nsew signal output
rlabel metal2 s 21546 169200 21602 170000 6 cache_PC[16]
port 8 nsew signal output
rlabel metal2 s 22558 169200 22614 170000 6 cache_PC[17]
port 9 nsew signal output
rlabel metal2 s 23570 169200 23626 170000 6 cache_PC[18]
port 10 nsew signal output
rlabel metal2 s 24582 169200 24638 170000 6 cache_PC[19]
port 11 nsew signal output
rlabel metal2 s 6366 169200 6422 170000 6 cache_PC[1]
port 12 nsew signal output
rlabel metal2 s 25594 169200 25650 170000 6 cache_PC[20]
port 13 nsew signal output
rlabel metal2 s 26606 169200 26662 170000 6 cache_PC[21]
port 14 nsew signal output
rlabel metal2 s 27618 169200 27674 170000 6 cache_PC[22]
port 15 nsew signal output
rlabel metal2 s 28630 169200 28686 170000 6 cache_PC[23]
port 16 nsew signal output
rlabel metal2 s 29642 169200 29698 170000 6 cache_PC[24]
port 17 nsew signal output
rlabel metal2 s 30654 169200 30710 170000 6 cache_PC[25]
port 18 nsew signal output
rlabel metal2 s 31666 169200 31722 170000 6 cache_PC[26]
port 19 nsew signal output
rlabel metal2 s 32678 169200 32734 170000 6 cache_PC[27]
port 20 nsew signal output
rlabel metal2 s 7378 169200 7434 170000 6 cache_PC[2]
port 21 nsew signal output
rlabel metal2 s 8390 169200 8446 170000 6 cache_PC[3]
port 22 nsew signal output
rlabel metal2 s 9402 169200 9458 170000 6 cache_PC[4]
port 23 nsew signal output
rlabel metal2 s 10414 169200 10470 170000 6 cache_PC[5]
port 24 nsew signal output
rlabel metal2 s 11426 169200 11482 170000 6 cache_PC[6]
port 25 nsew signal output
rlabel metal2 s 12438 169200 12494 170000 6 cache_PC[7]
port 26 nsew signal output
rlabel metal2 s 13450 169200 13506 170000 6 cache_PC[8]
port 27 nsew signal output
rlabel metal2 s 14462 169200 14518 170000 6 cache_PC[9]
port 28 nsew signal output
rlabel metal2 s 33690 169200 33746 170000 6 cache_entry[0]
port 29 nsew signal input
rlabel metal2 s 134890 169200 134946 170000 6 cache_entry[100]
port 30 nsew signal input
rlabel metal2 s 135902 169200 135958 170000 6 cache_entry[101]
port 31 nsew signal input
rlabel metal2 s 136914 169200 136970 170000 6 cache_entry[102]
port 32 nsew signal input
rlabel metal2 s 137926 169200 137982 170000 6 cache_entry[103]
port 33 nsew signal input
rlabel metal2 s 138938 169200 138994 170000 6 cache_entry[104]
port 34 nsew signal input
rlabel metal2 s 139950 169200 140006 170000 6 cache_entry[105]
port 35 nsew signal input
rlabel metal2 s 140962 169200 141018 170000 6 cache_entry[106]
port 36 nsew signal input
rlabel metal2 s 141974 169200 142030 170000 6 cache_entry[107]
port 37 nsew signal input
rlabel metal2 s 142986 169200 143042 170000 6 cache_entry[108]
port 38 nsew signal input
rlabel metal2 s 143998 169200 144054 170000 6 cache_entry[109]
port 39 nsew signal input
rlabel metal2 s 43810 169200 43866 170000 6 cache_entry[10]
port 40 nsew signal input
rlabel metal2 s 145010 169200 145066 170000 6 cache_entry[110]
port 41 nsew signal input
rlabel metal2 s 146022 169200 146078 170000 6 cache_entry[111]
port 42 nsew signal input
rlabel metal2 s 147034 169200 147090 170000 6 cache_entry[112]
port 43 nsew signal input
rlabel metal2 s 148046 169200 148102 170000 6 cache_entry[113]
port 44 nsew signal input
rlabel metal2 s 149058 169200 149114 170000 6 cache_entry[114]
port 45 nsew signal input
rlabel metal2 s 150070 169200 150126 170000 6 cache_entry[115]
port 46 nsew signal input
rlabel metal2 s 151082 169200 151138 170000 6 cache_entry[116]
port 47 nsew signal input
rlabel metal2 s 152094 169200 152150 170000 6 cache_entry[117]
port 48 nsew signal input
rlabel metal2 s 153106 169200 153162 170000 6 cache_entry[118]
port 49 nsew signal input
rlabel metal2 s 154118 169200 154174 170000 6 cache_entry[119]
port 50 nsew signal input
rlabel metal2 s 44822 169200 44878 170000 6 cache_entry[11]
port 51 nsew signal input
rlabel metal2 s 155130 169200 155186 170000 6 cache_entry[120]
port 52 nsew signal input
rlabel metal2 s 156142 169200 156198 170000 6 cache_entry[121]
port 53 nsew signal input
rlabel metal2 s 157154 169200 157210 170000 6 cache_entry[122]
port 54 nsew signal input
rlabel metal2 s 158166 169200 158222 170000 6 cache_entry[123]
port 55 nsew signal input
rlabel metal2 s 159178 169200 159234 170000 6 cache_entry[124]
port 56 nsew signal input
rlabel metal2 s 160190 169200 160246 170000 6 cache_entry[125]
port 57 nsew signal input
rlabel metal2 s 161202 169200 161258 170000 6 cache_entry[126]
port 58 nsew signal input
rlabel metal2 s 162214 169200 162270 170000 6 cache_entry[127]
port 59 nsew signal input
rlabel metal2 s 45834 169200 45890 170000 6 cache_entry[12]
port 60 nsew signal input
rlabel metal2 s 46846 169200 46902 170000 6 cache_entry[13]
port 61 nsew signal input
rlabel metal2 s 47858 169200 47914 170000 6 cache_entry[14]
port 62 nsew signal input
rlabel metal2 s 48870 169200 48926 170000 6 cache_entry[15]
port 63 nsew signal input
rlabel metal2 s 49882 169200 49938 170000 6 cache_entry[16]
port 64 nsew signal input
rlabel metal2 s 50894 169200 50950 170000 6 cache_entry[17]
port 65 nsew signal input
rlabel metal2 s 51906 169200 51962 170000 6 cache_entry[18]
port 66 nsew signal input
rlabel metal2 s 52918 169200 52974 170000 6 cache_entry[19]
port 67 nsew signal input
rlabel metal2 s 34702 169200 34758 170000 6 cache_entry[1]
port 68 nsew signal input
rlabel metal2 s 53930 169200 53986 170000 6 cache_entry[20]
port 69 nsew signal input
rlabel metal2 s 54942 169200 54998 170000 6 cache_entry[21]
port 70 nsew signal input
rlabel metal2 s 55954 169200 56010 170000 6 cache_entry[22]
port 71 nsew signal input
rlabel metal2 s 56966 169200 57022 170000 6 cache_entry[23]
port 72 nsew signal input
rlabel metal2 s 57978 169200 58034 170000 6 cache_entry[24]
port 73 nsew signal input
rlabel metal2 s 58990 169200 59046 170000 6 cache_entry[25]
port 74 nsew signal input
rlabel metal2 s 60002 169200 60058 170000 6 cache_entry[26]
port 75 nsew signal input
rlabel metal2 s 61014 169200 61070 170000 6 cache_entry[27]
port 76 nsew signal input
rlabel metal2 s 62026 169200 62082 170000 6 cache_entry[28]
port 77 nsew signal input
rlabel metal2 s 63038 169200 63094 170000 6 cache_entry[29]
port 78 nsew signal input
rlabel metal2 s 35714 169200 35770 170000 6 cache_entry[2]
port 79 nsew signal input
rlabel metal2 s 64050 169200 64106 170000 6 cache_entry[30]
port 80 nsew signal input
rlabel metal2 s 65062 169200 65118 170000 6 cache_entry[31]
port 81 nsew signal input
rlabel metal2 s 66074 169200 66130 170000 6 cache_entry[32]
port 82 nsew signal input
rlabel metal2 s 67086 169200 67142 170000 6 cache_entry[33]
port 83 nsew signal input
rlabel metal2 s 68098 169200 68154 170000 6 cache_entry[34]
port 84 nsew signal input
rlabel metal2 s 69110 169200 69166 170000 6 cache_entry[35]
port 85 nsew signal input
rlabel metal2 s 70122 169200 70178 170000 6 cache_entry[36]
port 86 nsew signal input
rlabel metal2 s 71134 169200 71190 170000 6 cache_entry[37]
port 87 nsew signal input
rlabel metal2 s 72146 169200 72202 170000 6 cache_entry[38]
port 88 nsew signal input
rlabel metal2 s 73158 169200 73214 170000 6 cache_entry[39]
port 89 nsew signal input
rlabel metal2 s 36726 169200 36782 170000 6 cache_entry[3]
port 90 nsew signal input
rlabel metal2 s 74170 169200 74226 170000 6 cache_entry[40]
port 91 nsew signal input
rlabel metal2 s 75182 169200 75238 170000 6 cache_entry[41]
port 92 nsew signal input
rlabel metal2 s 76194 169200 76250 170000 6 cache_entry[42]
port 93 nsew signal input
rlabel metal2 s 77206 169200 77262 170000 6 cache_entry[43]
port 94 nsew signal input
rlabel metal2 s 78218 169200 78274 170000 6 cache_entry[44]
port 95 nsew signal input
rlabel metal2 s 79230 169200 79286 170000 6 cache_entry[45]
port 96 nsew signal input
rlabel metal2 s 80242 169200 80298 170000 6 cache_entry[46]
port 97 nsew signal input
rlabel metal2 s 81254 169200 81310 170000 6 cache_entry[47]
port 98 nsew signal input
rlabel metal2 s 82266 169200 82322 170000 6 cache_entry[48]
port 99 nsew signal input
rlabel metal2 s 83278 169200 83334 170000 6 cache_entry[49]
port 100 nsew signal input
rlabel metal2 s 37738 169200 37794 170000 6 cache_entry[4]
port 101 nsew signal input
rlabel metal2 s 84290 169200 84346 170000 6 cache_entry[50]
port 102 nsew signal input
rlabel metal2 s 85302 169200 85358 170000 6 cache_entry[51]
port 103 nsew signal input
rlabel metal2 s 86314 169200 86370 170000 6 cache_entry[52]
port 104 nsew signal input
rlabel metal2 s 87326 169200 87382 170000 6 cache_entry[53]
port 105 nsew signal input
rlabel metal2 s 88338 169200 88394 170000 6 cache_entry[54]
port 106 nsew signal input
rlabel metal2 s 89350 169200 89406 170000 6 cache_entry[55]
port 107 nsew signal input
rlabel metal2 s 90362 169200 90418 170000 6 cache_entry[56]
port 108 nsew signal input
rlabel metal2 s 91374 169200 91430 170000 6 cache_entry[57]
port 109 nsew signal input
rlabel metal2 s 92386 169200 92442 170000 6 cache_entry[58]
port 110 nsew signal input
rlabel metal2 s 93398 169200 93454 170000 6 cache_entry[59]
port 111 nsew signal input
rlabel metal2 s 38750 169200 38806 170000 6 cache_entry[5]
port 112 nsew signal input
rlabel metal2 s 94410 169200 94466 170000 6 cache_entry[60]
port 113 nsew signal input
rlabel metal2 s 95422 169200 95478 170000 6 cache_entry[61]
port 114 nsew signal input
rlabel metal2 s 96434 169200 96490 170000 6 cache_entry[62]
port 115 nsew signal input
rlabel metal2 s 97446 169200 97502 170000 6 cache_entry[63]
port 116 nsew signal input
rlabel metal2 s 98458 169200 98514 170000 6 cache_entry[64]
port 117 nsew signal input
rlabel metal2 s 99470 169200 99526 170000 6 cache_entry[65]
port 118 nsew signal input
rlabel metal2 s 100482 169200 100538 170000 6 cache_entry[66]
port 119 nsew signal input
rlabel metal2 s 101494 169200 101550 170000 6 cache_entry[67]
port 120 nsew signal input
rlabel metal2 s 102506 169200 102562 170000 6 cache_entry[68]
port 121 nsew signal input
rlabel metal2 s 103518 169200 103574 170000 6 cache_entry[69]
port 122 nsew signal input
rlabel metal2 s 39762 169200 39818 170000 6 cache_entry[6]
port 123 nsew signal input
rlabel metal2 s 104530 169200 104586 170000 6 cache_entry[70]
port 124 nsew signal input
rlabel metal2 s 105542 169200 105598 170000 6 cache_entry[71]
port 125 nsew signal input
rlabel metal2 s 106554 169200 106610 170000 6 cache_entry[72]
port 126 nsew signal input
rlabel metal2 s 107566 169200 107622 170000 6 cache_entry[73]
port 127 nsew signal input
rlabel metal2 s 108578 169200 108634 170000 6 cache_entry[74]
port 128 nsew signal input
rlabel metal2 s 109590 169200 109646 170000 6 cache_entry[75]
port 129 nsew signal input
rlabel metal2 s 110602 169200 110658 170000 6 cache_entry[76]
port 130 nsew signal input
rlabel metal2 s 111614 169200 111670 170000 6 cache_entry[77]
port 131 nsew signal input
rlabel metal2 s 112626 169200 112682 170000 6 cache_entry[78]
port 132 nsew signal input
rlabel metal2 s 113638 169200 113694 170000 6 cache_entry[79]
port 133 nsew signal input
rlabel metal2 s 40774 169200 40830 170000 6 cache_entry[7]
port 134 nsew signal input
rlabel metal2 s 114650 169200 114706 170000 6 cache_entry[80]
port 135 nsew signal input
rlabel metal2 s 115662 169200 115718 170000 6 cache_entry[81]
port 136 nsew signal input
rlabel metal2 s 116674 169200 116730 170000 6 cache_entry[82]
port 137 nsew signal input
rlabel metal2 s 117686 169200 117742 170000 6 cache_entry[83]
port 138 nsew signal input
rlabel metal2 s 118698 169200 118754 170000 6 cache_entry[84]
port 139 nsew signal input
rlabel metal2 s 119710 169200 119766 170000 6 cache_entry[85]
port 140 nsew signal input
rlabel metal2 s 120722 169200 120778 170000 6 cache_entry[86]
port 141 nsew signal input
rlabel metal2 s 121734 169200 121790 170000 6 cache_entry[87]
port 142 nsew signal input
rlabel metal2 s 122746 169200 122802 170000 6 cache_entry[88]
port 143 nsew signal input
rlabel metal2 s 123758 169200 123814 170000 6 cache_entry[89]
port 144 nsew signal input
rlabel metal2 s 41786 169200 41842 170000 6 cache_entry[8]
port 145 nsew signal input
rlabel metal2 s 124770 169200 124826 170000 6 cache_entry[90]
port 146 nsew signal input
rlabel metal2 s 125782 169200 125838 170000 6 cache_entry[91]
port 147 nsew signal input
rlabel metal2 s 126794 169200 126850 170000 6 cache_entry[92]
port 148 nsew signal input
rlabel metal2 s 127806 169200 127862 170000 6 cache_entry[93]
port 149 nsew signal input
rlabel metal2 s 128818 169200 128874 170000 6 cache_entry[94]
port 150 nsew signal input
rlabel metal2 s 129830 169200 129886 170000 6 cache_entry[95]
port 151 nsew signal input
rlabel metal2 s 130842 169200 130898 170000 6 cache_entry[96]
port 152 nsew signal input
rlabel metal2 s 131854 169200 131910 170000 6 cache_entry[97]
port 153 nsew signal input
rlabel metal2 s 132866 169200 132922 170000 6 cache_entry[98]
port 154 nsew signal input
rlabel metal2 s 133878 169200 133934 170000 6 cache_entry[99]
port 155 nsew signal input
rlabel metal2 s 42798 169200 42854 170000 6 cache_entry[9]
port 156 nsew signal input
rlabel metal3 s 439200 20408 440000 20528 6 cache_entry_valid
port 157 nsew signal output
rlabel metal3 s 439200 18776 440000 18896 6 cache_hit
port 158 nsew signal input
rlabel metal3 s 439200 19320 440000 19440 6 cache_invalidate
port 159 nsew signal output
rlabel metal2 s 8390 0 8446 800 6 cache_new_entry[0]
port 160 nsew signal output
rlabel metal2 s 183190 0 183246 800 6 cache_new_entry[100]
port 161 nsew signal output
rlabel metal2 s 184938 0 184994 800 6 cache_new_entry[101]
port 162 nsew signal output
rlabel metal2 s 186686 0 186742 800 6 cache_new_entry[102]
port 163 nsew signal output
rlabel metal2 s 188434 0 188490 800 6 cache_new_entry[103]
port 164 nsew signal output
rlabel metal2 s 190182 0 190238 800 6 cache_new_entry[104]
port 165 nsew signal output
rlabel metal2 s 191930 0 191986 800 6 cache_new_entry[105]
port 166 nsew signal output
rlabel metal2 s 193678 0 193734 800 6 cache_new_entry[106]
port 167 nsew signal output
rlabel metal2 s 195426 0 195482 800 6 cache_new_entry[107]
port 168 nsew signal output
rlabel metal2 s 197174 0 197230 800 6 cache_new_entry[108]
port 169 nsew signal output
rlabel metal2 s 198922 0 198978 800 6 cache_new_entry[109]
port 170 nsew signal output
rlabel metal2 s 25870 0 25926 800 6 cache_new_entry[10]
port 171 nsew signal output
rlabel metal2 s 200670 0 200726 800 6 cache_new_entry[110]
port 172 nsew signal output
rlabel metal2 s 202418 0 202474 800 6 cache_new_entry[111]
port 173 nsew signal output
rlabel metal2 s 204166 0 204222 800 6 cache_new_entry[112]
port 174 nsew signal output
rlabel metal2 s 205914 0 205970 800 6 cache_new_entry[113]
port 175 nsew signal output
rlabel metal2 s 207662 0 207718 800 6 cache_new_entry[114]
port 176 nsew signal output
rlabel metal2 s 209410 0 209466 800 6 cache_new_entry[115]
port 177 nsew signal output
rlabel metal2 s 211158 0 211214 800 6 cache_new_entry[116]
port 178 nsew signal output
rlabel metal2 s 212906 0 212962 800 6 cache_new_entry[117]
port 179 nsew signal output
rlabel metal2 s 214654 0 214710 800 6 cache_new_entry[118]
port 180 nsew signal output
rlabel metal2 s 216402 0 216458 800 6 cache_new_entry[119]
port 181 nsew signal output
rlabel metal2 s 27618 0 27674 800 6 cache_new_entry[11]
port 182 nsew signal output
rlabel metal2 s 218150 0 218206 800 6 cache_new_entry[120]
port 183 nsew signal output
rlabel metal2 s 219898 0 219954 800 6 cache_new_entry[121]
port 184 nsew signal output
rlabel metal2 s 221646 0 221702 800 6 cache_new_entry[122]
port 185 nsew signal output
rlabel metal2 s 223394 0 223450 800 6 cache_new_entry[123]
port 186 nsew signal output
rlabel metal2 s 225142 0 225198 800 6 cache_new_entry[124]
port 187 nsew signal output
rlabel metal2 s 226890 0 226946 800 6 cache_new_entry[125]
port 188 nsew signal output
rlabel metal2 s 228638 0 228694 800 6 cache_new_entry[126]
port 189 nsew signal output
rlabel metal2 s 230386 0 230442 800 6 cache_new_entry[127]
port 190 nsew signal output
rlabel metal2 s 29366 0 29422 800 6 cache_new_entry[12]
port 191 nsew signal output
rlabel metal2 s 31114 0 31170 800 6 cache_new_entry[13]
port 192 nsew signal output
rlabel metal2 s 32862 0 32918 800 6 cache_new_entry[14]
port 193 nsew signal output
rlabel metal2 s 34610 0 34666 800 6 cache_new_entry[15]
port 194 nsew signal output
rlabel metal2 s 36358 0 36414 800 6 cache_new_entry[16]
port 195 nsew signal output
rlabel metal2 s 38106 0 38162 800 6 cache_new_entry[17]
port 196 nsew signal output
rlabel metal2 s 39854 0 39910 800 6 cache_new_entry[18]
port 197 nsew signal output
rlabel metal2 s 41602 0 41658 800 6 cache_new_entry[19]
port 198 nsew signal output
rlabel metal2 s 10138 0 10194 800 6 cache_new_entry[1]
port 199 nsew signal output
rlabel metal2 s 43350 0 43406 800 6 cache_new_entry[20]
port 200 nsew signal output
rlabel metal2 s 45098 0 45154 800 6 cache_new_entry[21]
port 201 nsew signal output
rlabel metal2 s 46846 0 46902 800 6 cache_new_entry[22]
port 202 nsew signal output
rlabel metal2 s 48594 0 48650 800 6 cache_new_entry[23]
port 203 nsew signal output
rlabel metal2 s 50342 0 50398 800 6 cache_new_entry[24]
port 204 nsew signal output
rlabel metal2 s 52090 0 52146 800 6 cache_new_entry[25]
port 205 nsew signal output
rlabel metal2 s 53838 0 53894 800 6 cache_new_entry[26]
port 206 nsew signal output
rlabel metal2 s 55586 0 55642 800 6 cache_new_entry[27]
port 207 nsew signal output
rlabel metal2 s 57334 0 57390 800 6 cache_new_entry[28]
port 208 nsew signal output
rlabel metal2 s 59082 0 59138 800 6 cache_new_entry[29]
port 209 nsew signal output
rlabel metal2 s 11886 0 11942 800 6 cache_new_entry[2]
port 210 nsew signal output
rlabel metal2 s 60830 0 60886 800 6 cache_new_entry[30]
port 211 nsew signal output
rlabel metal2 s 62578 0 62634 800 6 cache_new_entry[31]
port 212 nsew signal output
rlabel metal2 s 64326 0 64382 800 6 cache_new_entry[32]
port 213 nsew signal output
rlabel metal2 s 66074 0 66130 800 6 cache_new_entry[33]
port 214 nsew signal output
rlabel metal2 s 67822 0 67878 800 6 cache_new_entry[34]
port 215 nsew signal output
rlabel metal2 s 69570 0 69626 800 6 cache_new_entry[35]
port 216 nsew signal output
rlabel metal2 s 71318 0 71374 800 6 cache_new_entry[36]
port 217 nsew signal output
rlabel metal2 s 73066 0 73122 800 6 cache_new_entry[37]
port 218 nsew signal output
rlabel metal2 s 74814 0 74870 800 6 cache_new_entry[38]
port 219 nsew signal output
rlabel metal2 s 76562 0 76618 800 6 cache_new_entry[39]
port 220 nsew signal output
rlabel metal2 s 13634 0 13690 800 6 cache_new_entry[3]
port 221 nsew signal output
rlabel metal2 s 78310 0 78366 800 6 cache_new_entry[40]
port 222 nsew signal output
rlabel metal2 s 80058 0 80114 800 6 cache_new_entry[41]
port 223 nsew signal output
rlabel metal2 s 81806 0 81862 800 6 cache_new_entry[42]
port 224 nsew signal output
rlabel metal2 s 83554 0 83610 800 6 cache_new_entry[43]
port 225 nsew signal output
rlabel metal2 s 85302 0 85358 800 6 cache_new_entry[44]
port 226 nsew signal output
rlabel metal2 s 87050 0 87106 800 6 cache_new_entry[45]
port 227 nsew signal output
rlabel metal2 s 88798 0 88854 800 6 cache_new_entry[46]
port 228 nsew signal output
rlabel metal2 s 90546 0 90602 800 6 cache_new_entry[47]
port 229 nsew signal output
rlabel metal2 s 92294 0 92350 800 6 cache_new_entry[48]
port 230 nsew signal output
rlabel metal2 s 94042 0 94098 800 6 cache_new_entry[49]
port 231 nsew signal output
rlabel metal2 s 15382 0 15438 800 6 cache_new_entry[4]
port 232 nsew signal output
rlabel metal2 s 95790 0 95846 800 6 cache_new_entry[50]
port 233 nsew signal output
rlabel metal2 s 97538 0 97594 800 6 cache_new_entry[51]
port 234 nsew signal output
rlabel metal2 s 99286 0 99342 800 6 cache_new_entry[52]
port 235 nsew signal output
rlabel metal2 s 101034 0 101090 800 6 cache_new_entry[53]
port 236 nsew signal output
rlabel metal2 s 102782 0 102838 800 6 cache_new_entry[54]
port 237 nsew signal output
rlabel metal2 s 104530 0 104586 800 6 cache_new_entry[55]
port 238 nsew signal output
rlabel metal2 s 106278 0 106334 800 6 cache_new_entry[56]
port 239 nsew signal output
rlabel metal2 s 108026 0 108082 800 6 cache_new_entry[57]
port 240 nsew signal output
rlabel metal2 s 109774 0 109830 800 6 cache_new_entry[58]
port 241 nsew signal output
rlabel metal2 s 111522 0 111578 800 6 cache_new_entry[59]
port 242 nsew signal output
rlabel metal2 s 17130 0 17186 800 6 cache_new_entry[5]
port 243 nsew signal output
rlabel metal2 s 113270 0 113326 800 6 cache_new_entry[60]
port 244 nsew signal output
rlabel metal2 s 115018 0 115074 800 6 cache_new_entry[61]
port 245 nsew signal output
rlabel metal2 s 116766 0 116822 800 6 cache_new_entry[62]
port 246 nsew signal output
rlabel metal2 s 118514 0 118570 800 6 cache_new_entry[63]
port 247 nsew signal output
rlabel metal2 s 120262 0 120318 800 6 cache_new_entry[64]
port 248 nsew signal output
rlabel metal2 s 122010 0 122066 800 6 cache_new_entry[65]
port 249 nsew signal output
rlabel metal2 s 123758 0 123814 800 6 cache_new_entry[66]
port 250 nsew signal output
rlabel metal2 s 125506 0 125562 800 6 cache_new_entry[67]
port 251 nsew signal output
rlabel metal2 s 127254 0 127310 800 6 cache_new_entry[68]
port 252 nsew signal output
rlabel metal2 s 129002 0 129058 800 6 cache_new_entry[69]
port 253 nsew signal output
rlabel metal2 s 18878 0 18934 800 6 cache_new_entry[6]
port 254 nsew signal output
rlabel metal2 s 130750 0 130806 800 6 cache_new_entry[70]
port 255 nsew signal output
rlabel metal2 s 132498 0 132554 800 6 cache_new_entry[71]
port 256 nsew signal output
rlabel metal2 s 134246 0 134302 800 6 cache_new_entry[72]
port 257 nsew signal output
rlabel metal2 s 135994 0 136050 800 6 cache_new_entry[73]
port 258 nsew signal output
rlabel metal2 s 137742 0 137798 800 6 cache_new_entry[74]
port 259 nsew signal output
rlabel metal2 s 139490 0 139546 800 6 cache_new_entry[75]
port 260 nsew signal output
rlabel metal2 s 141238 0 141294 800 6 cache_new_entry[76]
port 261 nsew signal output
rlabel metal2 s 142986 0 143042 800 6 cache_new_entry[77]
port 262 nsew signal output
rlabel metal2 s 144734 0 144790 800 6 cache_new_entry[78]
port 263 nsew signal output
rlabel metal2 s 146482 0 146538 800 6 cache_new_entry[79]
port 264 nsew signal output
rlabel metal2 s 20626 0 20682 800 6 cache_new_entry[7]
port 265 nsew signal output
rlabel metal2 s 148230 0 148286 800 6 cache_new_entry[80]
port 266 nsew signal output
rlabel metal2 s 149978 0 150034 800 6 cache_new_entry[81]
port 267 nsew signal output
rlabel metal2 s 151726 0 151782 800 6 cache_new_entry[82]
port 268 nsew signal output
rlabel metal2 s 153474 0 153530 800 6 cache_new_entry[83]
port 269 nsew signal output
rlabel metal2 s 155222 0 155278 800 6 cache_new_entry[84]
port 270 nsew signal output
rlabel metal2 s 156970 0 157026 800 6 cache_new_entry[85]
port 271 nsew signal output
rlabel metal2 s 158718 0 158774 800 6 cache_new_entry[86]
port 272 nsew signal output
rlabel metal2 s 160466 0 160522 800 6 cache_new_entry[87]
port 273 nsew signal output
rlabel metal2 s 162214 0 162270 800 6 cache_new_entry[88]
port 274 nsew signal output
rlabel metal2 s 163962 0 164018 800 6 cache_new_entry[89]
port 275 nsew signal output
rlabel metal2 s 22374 0 22430 800 6 cache_new_entry[8]
port 276 nsew signal output
rlabel metal2 s 165710 0 165766 800 6 cache_new_entry[90]
port 277 nsew signal output
rlabel metal2 s 167458 0 167514 800 6 cache_new_entry[91]
port 278 nsew signal output
rlabel metal2 s 169206 0 169262 800 6 cache_new_entry[92]
port 279 nsew signal output
rlabel metal2 s 170954 0 171010 800 6 cache_new_entry[93]
port 280 nsew signal output
rlabel metal2 s 172702 0 172758 800 6 cache_new_entry[94]
port 281 nsew signal output
rlabel metal2 s 174450 0 174506 800 6 cache_new_entry[95]
port 282 nsew signal output
rlabel metal2 s 176198 0 176254 800 6 cache_new_entry[96]
port 283 nsew signal output
rlabel metal2 s 177946 0 178002 800 6 cache_new_entry[97]
port 284 nsew signal output
rlabel metal2 s 179694 0 179750 800 6 cache_new_entry[98]
port 285 nsew signal output
rlabel metal2 s 181442 0 181498 800 6 cache_new_entry[99]
port 286 nsew signal output
rlabel metal2 s 24122 0 24178 800 6 cache_new_entry[9]
port 287 nsew signal output
rlabel metal3 s 439200 19864 440000 19984 6 cache_rst
port 288 nsew signal output
rlabel metal2 s 164238 169200 164294 170000 6 curr_PC[0]
port 289 nsew signal output
rlabel metal2 s 174358 169200 174414 170000 6 curr_PC[10]
port 290 nsew signal output
rlabel metal2 s 175370 169200 175426 170000 6 curr_PC[11]
port 291 nsew signal output
rlabel metal2 s 176382 169200 176438 170000 6 curr_PC[12]
port 292 nsew signal output
rlabel metal2 s 177394 169200 177450 170000 6 curr_PC[13]
port 293 nsew signal output
rlabel metal2 s 178406 169200 178462 170000 6 curr_PC[14]
port 294 nsew signal output
rlabel metal2 s 179418 169200 179474 170000 6 curr_PC[15]
port 295 nsew signal output
rlabel metal2 s 180430 169200 180486 170000 6 curr_PC[16]
port 296 nsew signal output
rlabel metal2 s 181442 169200 181498 170000 6 curr_PC[17]
port 297 nsew signal output
rlabel metal2 s 182454 169200 182510 170000 6 curr_PC[18]
port 298 nsew signal output
rlabel metal2 s 183466 169200 183522 170000 6 curr_PC[19]
port 299 nsew signal output
rlabel metal2 s 165250 169200 165306 170000 6 curr_PC[1]
port 300 nsew signal output
rlabel metal2 s 184478 169200 184534 170000 6 curr_PC[20]
port 301 nsew signal output
rlabel metal2 s 185490 169200 185546 170000 6 curr_PC[21]
port 302 nsew signal output
rlabel metal2 s 186502 169200 186558 170000 6 curr_PC[22]
port 303 nsew signal output
rlabel metal2 s 187514 169200 187570 170000 6 curr_PC[23]
port 304 nsew signal output
rlabel metal2 s 188526 169200 188582 170000 6 curr_PC[24]
port 305 nsew signal output
rlabel metal2 s 189538 169200 189594 170000 6 curr_PC[25]
port 306 nsew signal output
rlabel metal2 s 190550 169200 190606 170000 6 curr_PC[26]
port 307 nsew signal output
rlabel metal2 s 191562 169200 191618 170000 6 curr_PC[27]
port 308 nsew signal output
rlabel metal2 s 166262 169200 166318 170000 6 curr_PC[2]
port 309 nsew signal output
rlabel metal2 s 167274 169200 167330 170000 6 curr_PC[3]
port 310 nsew signal output
rlabel metal2 s 168286 169200 168342 170000 6 curr_PC[4]
port 311 nsew signal output
rlabel metal2 s 169298 169200 169354 170000 6 curr_PC[5]
port 312 nsew signal output
rlabel metal2 s 170310 169200 170366 170000 6 curr_PC[6]
port 313 nsew signal output
rlabel metal2 s 171322 169200 171378 170000 6 curr_PC[7]
port 314 nsew signal output
rlabel metal2 s 172334 169200 172390 170000 6 curr_PC[8]
port 315 nsew signal output
rlabel metal2 s 173346 169200 173402 170000 6 curr_PC[9]
port 316 nsew signal output
rlabel metal2 s 424414 0 424470 800 6 custom_settings[0]
port 317 nsew signal input
rlabel metal2 s 426162 0 426218 800 6 custom_settings[1]
port 318 nsew signal input
rlabel metal2 s 427910 0 427966 800 6 custom_settings[2]
port 319 nsew signal input
rlabel metal2 s 429658 0 429714 800 6 custom_settings[3]
port 320 nsew signal input
rlabel metal2 s 431406 0 431462 800 6 custom_settings[4]
port 321 nsew signal input
rlabel metal2 s 239126 169200 239182 170000 6 dest_idx0[0]
port 322 nsew signal input
rlabel metal2 s 240138 169200 240194 170000 6 dest_idx0[1]
port 323 nsew signal input
rlabel metal2 s 241150 169200 241206 170000 6 dest_idx0[2]
port 324 nsew signal input
rlabel metal2 s 242162 169200 242218 170000 6 dest_idx0[3]
port 325 nsew signal input
rlabel metal2 s 243174 169200 243230 170000 6 dest_idx0[4]
port 326 nsew signal input
rlabel metal2 s 244186 169200 244242 170000 6 dest_idx0[5]
port 327 nsew signal input
rlabel metal3 s 439200 45976 440000 46096 6 dest_idx1[0]
port 328 nsew signal input
rlabel metal3 s 439200 46520 440000 46640 6 dest_idx1[1]
port 329 nsew signal input
rlabel metal3 s 439200 47064 440000 47184 6 dest_idx1[2]
port 330 nsew signal input
rlabel metal3 s 439200 47608 440000 47728 6 dest_idx1[3]
port 331 nsew signal input
rlabel metal3 s 439200 48152 440000 48272 6 dest_idx1[4]
port 332 nsew signal input
rlabel metal3 s 439200 48696 440000 48816 6 dest_idx1[5]
port 333 nsew signal input
rlabel metal3 s 0 44888 800 45008 6 dest_idx2[0]
port 334 nsew signal input
rlabel metal3 s 0 45432 800 45552 6 dest_idx2[1]
port 335 nsew signal input
rlabel metal3 s 0 45976 800 46096 6 dest_idx2[2]
port 336 nsew signal input
rlabel metal3 s 0 46520 800 46640 6 dest_idx2[3]
port 337 nsew signal input
rlabel metal3 s 0 47064 800 47184 6 dest_idx2[4]
port 338 nsew signal input
rlabel metal3 s 0 47608 800 47728 6 dest_idx2[5]
port 339 nsew signal input
rlabel metal2 s 237102 169200 237158 170000 6 dest_mask0[0]
port 340 nsew signal input
rlabel metal2 s 238114 169200 238170 170000 6 dest_mask0[1]
port 341 nsew signal input
rlabel metal3 s 439200 44888 440000 45008 6 dest_mask1[0]
port 342 nsew signal input
rlabel metal3 s 439200 45432 440000 45552 6 dest_mask1[1]
port 343 nsew signal input
rlabel metal3 s 0 43800 800 43920 6 dest_mask2[0]
port 344 nsew signal input
rlabel metal3 s 0 44344 800 44464 6 dest_mask2[1]
port 345 nsew signal input
rlabel metal2 s 248234 169200 248290 170000 6 dest_pred0[0]
port 346 nsew signal input
rlabel metal2 s 249246 169200 249302 170000 6 dest_pred0[1]
port 347 nsew signal input
rlabel metal2 s 250258 169200 250314 170000 6 dest_pred0[2]
port 348 nsew signal input
rlabel metal3 s 439200 50872 440000 50992 6 dest_pred1[0]
port 349 nsew signal input
rlabel metal3 s 439200 51416 440000 51536 6 dest_pred1[1]
port 350 nsew signal input
rlabel metal3 s 439200 51960 440000 52080 6 dest_pred1[2]
port 351 nsew signal input
rlabel metal3 s 0 49784 800 49904 6 dest_pred2[0]
port 352 nsew signal input
rlabel metal3 s 0 50328 800 50448 6 dest_pred2[1]
port 353 nsew signal input
rlabel metal3 s 0 50872 800 50992 6 dest_pred2[2]
port 354 nsew signal input
rlabel metal2 s 251270 169200 251326 170000 6 dest_pred_val0
port 355 nsew signal input
rlabel metal3 s 439200 52504 440000 52624 6 dest_pred_val1
port 356 nsew signal input
rlabel metal3 s 0 51416 800 51536 6 dest_pred_val2
port 357 nsew signal input
rlabel metal2 s 204718 169200 204774 170000 6 dest_val0[0]
port 358 nsew signal input
rlabel metal2 s 214838 169200 214894 170000 6 dest_val0[10]
port 359 nsew signal input
rlabel metal2 s 215850 169200 215906 170000 6 dest_val0[11]
port 360 nsew signal input
rlabel metal2 s 216862 169200 216918 170000 6 dest_val0[12]
port 361 nsew signal input
rlabel metal2 s 217874 169200 217930 170000 6 dest_val0[13]
port 362 nsew signal input
rlabel metal2 s 218886 169200 218942 170000 6 dest_val0[14]
port 363 nsew signal input
rlabel metal2 s 219898 169200 219954 170000 6 dest_val0[15]
port 364 nsew signal input
rlabel metal2 s 220910 169200 220966 170000 6 dest_val0[16]
port 365 nsew signal input
rlabel metal2 s 221922 169200 221978 170000 6 dest_val0[17]
port 366 nsew signal input
rlabel metal2 s 222934 169200 222990 170000 6 dest_val0[18]
port 367 nsew signal input
rlabel metal2 s 223946 169200 224002 170000 6 dest_val0[19]
port 368 nsew signal input
rlabel metal2 s 205730 169200 205786 170000 6 dest_val0[1]
port 369 nsew signal input
rlabel metal2 s 224958 169200 225014 170000 6 dest_val0[20]
port 370 nsew signal input
rlabel metal2 s 225970 169200 226026 170000 6 dest_val0[21]
port 371 nsew signal input
rlabel metal2 s 226982 169200 227038 170000 6 dest_val0[22]
port 372 nsew signal input
rlabel metal2 s 227994 169200 228050 170000 6 dest_val0[23]
port 373 nsew signal input
rlabel metal2 s 229006 169200 229062 170000 6 dest_val0[24]
port 374 nsew signal input
rlabel metal2 s 230018 169200 230074 170000 6 dest_val0[25]
port 375 nsew signal input
rlabel metal2 s 231030 169200 231086 170000 6 dest_val0[26]
port 376 nsew signal input
rlabel metal2 s 232042 169200 232098 170000 6 dest_val0[27]
port 377 nsew signal input
rlabel metal2 s 233054 169200 233110 170000 6 dest_val0[28]
port 378 nsew signal input
rlabel metal2 s 234066 169200 234122 170000 6 dest_val0[29]
port 379 nsew signal input
rlabel metal2 s 206742 169200 206798 170000 6 dest_val0[2]
port 380 nsew signal input
rlabel metal2 s 235078 169200 235134 170000 6 dest_val0[30]
port 381 nsew signal input
rlabel metal2 s 236090 169200 236146 170000 6 dest_val0[31]
port 382 nsew signal input
rlabel metal2 s 207754 169200 207810 170000 6 dest_val0[3]
port 383 nsew signal input
rlabel metal2 s 208766 169200 208822 170000 6 dest_val0[4]
port 384 nsew signal input
rlabel metal2 s 209778 169200 209834 170000 6 dest_val0[5]
port 385 nsew signal input
rlabel metal2 s 210790 169200 210846 170000 6 dest_val0[6]
port 386 nsew signal input
rlabel metal2 s 211802 169200 211858 170000 6 dest_val0[7]
port 387 nsew signal input
rlabel metal2 s 212814 169200 212870 170000 6 dest_val0[8]
port 388 nsew signal input
rlabel metal2 s 213826 169200 213882 170000 6 dest_val0[9]
port 389 nsew signal input
rlabel metal3 s 439200 27480 440000 27600 6 dest_val1[0]
port 390 nsew signal input
rlabel metal3 s 439200 32920 440000 33040 6 dest_val1[10]
port 391 nsew signal input
rlabel metal3 s 439200 33464 440000 33584 6 dest_val1[11]
port 392 nsew signal input
rlabel metal3 s 439200 34008 440000 34128 6 dest_val1[12]
port 393 nsew signal input
rlabel metal3 s 439200 34552 440000 34672 6 dest_val1[13]
port 394 nsew signal input
rlabel metal3 s 439200 35096 440000 35216 6 dest_val1[14]
port 395 nsew signal input
rlabel metal3 s 439200 35640 440000 35760 6 dest_val1[15]
port 396 nsew signal input
rlabel metal3 s 439200 36184 440000 36304 6 dest_val1[16]
port 397 nsew signal input
rlabel metal3 s 439200 36728 440000 36848 6 dest_val1[17]
port 398 nsew signal input
rlabel metal3 s 439200 37272 440000 37392 6 dest_val1[18]
port 399 nsew signal input
rlabel metal3 s 439200 37816 440000 37936 6 dest_val1[19]
port 400 nsew signal input
rlabel metal3 s 439200 28024 440000 28144 6 dest_val1[1]
port 401 nsew signal input
rlabel metal3 s 439200 38360 440000 38480 6 dest_val1[20]
port 402 nsew signal input
rlabel metal3 s 439200 38904 440000 39024 6 dest_val1[21]
port 403 nsew signal input
rlabel metal3 s 439200 39448 440000 39568 6 dest_val1[22]
port 404 nsew signal input
rlabel metal3 s 439200 39992 440000 40112 6 dest_val1[23]
port 405 nsew signal input
rlabel metal3 s 439200 40536 440000 40656 6 dest_val1[24]
port 406 nsew signal input
rlabel metal3 s 439200 41080 440000 41200 6 dest_val1[25]
port 407 nsew signal input
rlabel metal3 s 439200 41624 440000 41744 6 dest_val1[26]
port 408 nsew signal input
rlabel metal3 s 439200 42168 440000 42288 6 dest_val1[27]
port 409 nsew signal input
rlabel metal3 s 439200 42712 440000 42832 6 dest_val1[28]
port 410 nsew signal input
rlabel metal3 s 439200 43256 440000 43376 6 dest_val1[29]
port 411 nsew signal input
rlabel metal3 s 439200 28568 440000 28688 6 dest_val1[2]
port 412 nsew signal input
rlabel metal3 s 439200 43800 440000 43920 6 dest_val1[30]
port 413 nsew signal input
rlabel metal3 s 439200 44344 440000 44464 6 dest_val1[31]
port 414 nsew signal input
rlabel metal3 s 439200 29112 440000 29232 6 dest_val1[3]
port 415 nsew signal input
rlabel metal3 s 439200 29656 440000 29776 6 dest_val1[4]
port 416 nsew signal input
rlabel metal3 s 439200 30200 440000 30320 6 dest_val1[5]
port 417 nsew signal input
rlabel metal3 s 439200 30744 440000 30864 6 dest_val1[6]
port 418 nsew signal input
rlabel metal3 s 439200 31288 440000 31408 6 dest_val1[7]
port 419 nsew signal input
rlabel metal3 s 439200 31832 440000 31952 6 dest_val1[8]
port 420 nsew signal input
rlabel metal3 s 439200 32376 440000 32496 6 dest_val1[9]
port 421 nsew signal input
rlabel metal3 s 0 26392 800 26512 6 dest_val2[0]
port 422 nsew signal input
rlabel metal3 s 0 31832 800 31952 6 dest_val2[10]
port 423 nsew signal input
rlabel metal3 s 0 32376 800 32496 6 dest_val2[11]
port 424 nsew signal input
rlabel metal3 s 0 32920 800 33040 6 dest_val2[12]
port 425 nsew signal input
rlabel metal3 s 0 33464 800 33584 6 dest_val2[13]
port 426 nsew signal input
rlabel metal3 s 0 34008 800 34128 6 dest_val2[14]
port 427 nsew signal input
rlabel metal3 s 0 34552 800 34672 6 dest_val2[15]
port 428 nsew signal input
rlabel metal3 s 0 35096 800 35216 6 dest_val2[16]
port 429 nsew signal input
rlabel metal3 s 0 35640 800 35760 6 dest_val2[17]
port 430 nsew signal input
rlabel metal3 s 0 36184 800 36304 6 dest_val2[18]
port 431 nsew signal input
rlabel metal3 s 0 36728 800 36848 6 dest_val2[19]
port 432 nsew signal input
rlabel metal3 s 0 26936 800 27056 6 dest_val2[1]
port 433 nsew signal input
rlabel metal3 s 0 37272 800 37392 6 dest_val2[20]
port 434 nsew signal input
rlabel metal3 s 0 37816 800 37936 6 dest_val2[21]
port 435 nsew signal input
rlabel metal3 s 0 38360 800 38480 6 dest_val2[22]
port 436 nsew signal input
rlabel metal3 s 0 38904 800 39024 6 dest_val2[23]
port 437 nsew signal input
rlabel metal3 s 0 39448 800 39568 6 dest_val2[24]
port 438 nsew signal input
rlabel metal3 s 0 39992 800 40112 6 dest_val2[25]
port 439 nsew signal input
rlabel metal3 s 0 40536 800 40656 6 dest_val2[26]
port 440 nsew signal input
rlabel metal3 s 0 41080 800 41200 6 dest_val2[27]
port 441 nsew signal input
rlabel metal3 s 0 41624 800 41744 6 dest_val2[28]
port 442 nsew signal input
rlabel metal3 s 0 42168 800 42288 6 dest_val2[29]
port 443 nsew signal input
rlabel metal3 s 0 27480 800 27600 6 dest_val2[2]
port 444 nsew signal input
rlabel metal3 s 0 42712 800 42832 6 dest_val2[30]
port 445 nsew signal input
rlabel metal3 s 0 43256 800 43376 6 dest_val2[31]
port 446 nsew signal input
rlabel metal3 s 0 28024 800 28144 6 dest_val2[3]
port 447 nsew signal input
rlabel metal3 s 0 28568 800 28688 6 dest_val2[4]
port 448 nsew signal input
rlabel metal3 s 0 29112 800 29232 6 dest_val2[5]
port 449 nsew signal input
rlabel metal3 s 0 29656 800 29776 6 dest_val2[6]
port 450 nsew signal input
rlabel metal3 s 0 30200 800 30320 6 dest_val2[7]
port 451 nsew signal input
rlabel metal3 s 0 30744 800 30864 6 dest_val2[8]
port 452 nsew signal input
rlabel metal3 s 0 31288 800 31408 6 dest_val2[9]
port 453 nsew signal input
rlabel metal2 s 325146 169200 325202 170000 6 eu0_busy
port 454 nsew signal input
rlabel metal2 s 326158 169200 326214 170000 6 eu0_instruction[0]
port 455 nsew signal output
rlabel metal2 s 336278 169200 336334 170000 6 eu0_instruction[10]
port 456 nsew signal output
rlabel metal2 s 337290 169200 337346 170000 6 eu0_instruction[11]
port 457 nsew signal output
rlabel metal2 s 338302 169200 338358 170000 6 eu0_instruction[12]
port 458 nsew signal output
rlabel metal2 s 339314 169200 339370 170000 6 eu0_instruction[13]
port 459 nsew signal output
rlabel metal2 s 340326 169200 340382 170000 6 eu0_instruction[14]
port 460 nsew signal output
rlabel metal2 s 341338 169200 341394 170000 6 eu0_instruction[15]
port 461 nsew signal output
rlabel metal2 s 342350 169200 342406 170000 6 eu0_instruction[16]
port 462 nsew signal output
rlabel metal2 s 343362 169200 343418 170000 6 eu0_instruction[17]
port 463 nsew signal output
rlabel metal2 s 344374 169200 344430 170000 6 eu0_instruction[18]
port 464 nsew signal output
rlabel metal2 s 345386 169200 345442 170000 6 eu0_instruction[19]
port 465 nsew signal output
rlabel metal2 s 327170 169200 327226 170000 6 eu0_instruction[1]
port 466 nsew signal output
rlabel metal2 s 346398 169200 346454 170000 6 eu0_instruction[20]
port 467 nsew signal output
rlabel metal2 s 347410 169200 347466 170000 6 eu0_instruction[21]
port 468 nsew signal output
rlabel metal2 s 348422 169200 348478 170000 6 eu0_instruction[22]
port 469 nsew signal output
rlabel metal2 s 349434 169200 349490 170000 6 eu0_instruction[23]
port 470 nsew signal output
rlabel metal2 s 350446 169200 350502 170000 6 eu0_instruction[24]
port 471 nsew signal output
rlabel metal2 s 351458 169200 351514 170000 6 eu0_instruction[25]
port 472 nsew signal output
rlabel metal2 s 352470 169200 352526 170000 6 eu0_instruction[26]
port 473 nsew signal output
rlabel metal2 s 353482 169200 353538 170000 6 eu0_instruction[27]
port 474 nsew signal output
rlabel metal2 s 354494 169200 354550 170000 6 eu0_instruction[28]
port 475 nsew signal output
rlabel metal2 s 355506 169200 355562 170000 6 eu0_instruction[29]
port 476 nsew signal output
rlabel metal2 s 328182 169200 328238 170000 6 eu0_instruction[2]
port 477 nsew signal output
rlabel metal2 s 356518 169200 356574 170000 6 eu0_instruction[30]
port 478 nsew signal output
rlabel metal2 s 357530 169200 357586 170000 6 eu0_instruction[31]
port 479 nsew signal output
rlabel metal2 s 358542 169200 358598 170000 6 eu0_instruction[32]
port 480 nsew signal output
rlabel metal2 s 359554 169200 359610 170000 6 eu0_instruction[33]
port 481 nsew signal output
rlabel metal2 s 360566 169200 360622 170000 6 eu0_instruction[34]
port 482 nsew signal output
rlabel metal2 s 361578 169200 361634 170000 6 eu0_instruction[35]
port 483 nsew signal output
rlabel metal2 s 362590 169200 362646 170000 6 eu0_instruction[36]
port 484 nsew signal output
rlabel metal2 s 363602 169200 363658 170000 6 eu0_instruction[37]
port 485 nsew signal output
rlabel metal2 s 364614 169200 364670 170000 6 eu0_instruction[38]
port 486 nsew signal output
rlabel metal2 s 365626 169200 365682 170000 6 eu0_instruction[39]
port 487 nsew signal output
rlabel metal2 s 329194 169200 329250 170000 6 eu0_instruction[3]
port 488 nsew signal output
rlabel metal2 s 366638 169200 366694 170000 6 eu0_instruction[40]
port 489 nsew signal output
rlabel metal2 s 367650 169200 367706 170000 6 eu0_instruction[41]
port 490 nsew signal output
rlabel metal2 s 330206 169200 330262 170000 6 eu0_instruction[4]
port 491 nsew signal output
rlabel metal2 s 331218 169200 331274 170000 6 eu0_instruction[5]
port 492 nsew signal output
rlabel metal2 s 332230 169200 332286 170000 6 eu0_instruction[6]
port 493 nsew signal output
rlabel metal2 s 333242 169200 333298 170000 6 eu0_instruction[7]
port 494 nsew signal output
rlabel metal2 s 334254 169200 334310 170000 6 eu0_instruction[8]
port 495 nsew signal output
rlabel metal2 s 335266 169200 335322 170000 6 eu0_instruction[9]
port 496 nsew signal output
rlabel metal3 s 439200 92216 440000 92336 6 eu1_busy
port 497 nsew signal input
rlabel metal3 s 439200 92760 440000 92880 6 eu1_instruction[0]
port 498 nsew signal output
rlabel metal3 s 439200 98200 440000 98320 6 eu1_instruction[10]
port 499 nsew signal output
rlabel metal3 s 439200 98744 440000 98864 6 eu1_instruction[11]
port 500 nsew signal output
rlabel metal3 s 439200 99288 440000 99408 6 eu1_instruction[12]
port 501 nsew signal output
rlabel metal3 s 439200 99832 440000 99952 6 eu1_instruction[13]
port 502 nsew signal output
rlabel metal3 s 439200 100376 440000 100496 6 eu1_instruction[14]
port 503 nsew signal output
rlabel metal3 s 439200 100920 440000 101040 6 eu1_instruction[15]
port 504 nsew signal output
rlabel metal3 s 439200 101464 440000 101584 6 eu1_instruction[16]
port 505 nsew signal output
rlabel metal3 s 439200 102008 440000 102128 6 eu1_instruction[17]
port 506 nsew signal output
rlabel metal3 s 439200 102552 440000 102672 6 eu1_instruction[18]
port 507 nsew signal output
rlabel metal3 s 439200 103096 440000 103216 6 eu1_instruction[19]
port 508 nsew signal output
rlabel metal3 s 439200 93304 440000 93424 6 eu1_instruction[1]
port 509 nsew signal output
rlabel metal3 s 439200 103640 440000 103760 6 eu1_instruction[20]
port 510 nsew signal output
rlabel metal3 s 439200 104184 440000 104304 6 eu1_instruction[21]
port 511 nsew signal output
rlabel metal3 s 439200 104728 440000 104848 6 eu1_instruction[22]
port 512 nsew signal output
rlabel metal3 s 439200 105272 440000 105392 6 eu1_instruction[23]
port 513 nsew signal output
rlabel metal3 s 439200 105816 440000 105936 6 eu1_instruction[24]
port 514 nsew signal output
rlabel metal3 s 439200 106360 440000 106480 6 eu1_instruction[25]
port 515 nsew signal output
rlabel metal3 s 439200 106904 440000 107024 6 eu1_instruction[26]
port 516 nsew signal output
rlabel metal3 s 439200 107448 440000 107568 6 eu1_instruction[27]
port 517 nsew signal output
rlabel metal3 s 439200 107992 440000 108112 6 eu1_instruction[28]
port 518 nsew signal output
rlabel metal3 s 439200 108536 440000 108656 6 eu1_instruction[29]
port 519 nsew signal output
rlabel metal3 s 439200 93848 440000 93968 6 eu1_instruction[2]
port 520 nsew signal output
rlabel metal3 s 439200 109080 440000 109200 6 eu1_instruction[30]
port 521 nsew signal output
rlabel metal3 s 439200 109624 440000 109744 6 eu1_instruction[31]
port 522 nsew signal output
rlabel metal3 s 439200 110168 440000 110288 6 eu1_instruction[32]
port 523 nsew signal output
rlabel metal3 s 439200 110712 440000 110832 6 eu1_instruction[33]
port 524 nsew signal output
rlabel metal3 s 439200 111256 440000 111376 6 eu1_instruction[34]
port 525 nsew signal output
rlabel metal3 s 439200 111800 440000 111920 6 eu1_instruction[35]
port 526 nsew signal output
rlabel metal3 s 439200 112344 440000 112464 6 eu1_instruction[36]
port 527 nsew signal output
rlabel metal3 s 439200 112888 440000 113008 6 eu1_instruction[37]
port 528 nsew signal output
rlabel metal3 s 439200 113432 440000 113552 6 eu1_instruction[38]
port 529 nsew signal output
rlabel metal3 s 439200 113976 440000 114096 6 eu1_instruction[39]
port 530 nsew signal output
rlabel metal3 s 439200 94392 440000 94512 6 eu1_instruction[3]
port 531 nsew signal output
rlabel metal3 s 439200 114520 440000 114640 6 eu1_instruction[40]
port 532 nsew signal output
rlabel metal3 s 439200 115064 440000 115184 6 eu1_instruction[41]
port 533 nsew signal output
rlabel metal3 s 439200 94936 440000 95056 6 eu1_instruction[4]
port 534 nsew signal output
rlabel metal3 s 439200 95480 440000 95600 6 eu1_instruction[5]
port 535 nsew signal output
rlabel metal3 s 439200 96024 440000 96144 6 eu1_instruction[6]
port 536 nsew signal output
rlabel metal3 s 439200 96568 440000 96688 6 eu1_instruction[7]
port 537 nsew signal output
rlabel metal3 s 439200 97112 440000 97232 6 eu1_instruction[8]
port 538 nsew signal output
rlabel metal3 s 439200 97656 440000 97776 6 eu1_instruction[9]
port 539 nsew signal output
rlabel metal3 s 0 91128 800 91248 6 eu2_busy
port 540 nsew signal input
rlabel metal3 s 0 91672 800 91792 6 eu2_instruction[0]
port 541 nsew signal output
rlabel metal3 s 0 97112 800 97232 6 eu2_instruction[10]
port 542 nsew signal output
rlabel metal3 s 0 97656 800 97776 6 eu2_instruction[11]
port 543 nsew signal output
rlabel metal3 s 0 98200 800 98320 6 eu2_instruction[12]
port 544 nsew signal output
rlabel metal3 s 0 98744 800 98864 6 eu2_instruction[13]
port 545 nsew signal output
rlabel metal3 s 0 99288 800 99408 6 eu2_instruction[14]
port 546 nsew signal output
rlabel metal3 s 0 99832 800 99952 6 eu2_instruction[15]
port 547 nsew signal output
rlabel metal3 s 0 100376 800 100496 6 eu2_instruction[16]
port 548 nsew signal output
rlabel metal3 s 0 100920 800 101040 6 eu2_instruction[17]
port 549 nsew signal output
rlabel metal3 s 0 101464 800 101584 6 eu2_instruction[18]
port 550 nsew signal output
rlabel metal3 s 0 102008 800 102128 6 eu2_instruction[19]
port 551 nsew signal output
rlabel metal3 s 0 92216 800 92336 6 eu2_instruction[1]
port 552 nsew signal output
rlabel metal3 s 0 102552 800 102672 6 eu2_instruction[20]
port 553 nsew signal output
rlabel metal3 s 0 103096 800 103216 6 eu2_instruction[21]
port 554 nsew signal output
rlabel metal3 s 0 103640 800 103760 6 eu2_instruction[22]
port 555 nsew signal output
rlabel metal3 s 0 104184 800 104304 6 eu2_instruction[23]
port 556 nsew signal output
rlabel metal3 s 0 104728 800 104848 6 eu2_instruction[24]
port 557 nsew signal output
rlabel metal3 s 0 105272 800 105392 6 eu2_instruction[25]
port 558 nsew signal output
rlabel metal3 s 0 105816 800 105936 6 eu2_instruction[26]
port 559 nsew signal output
rlabel metal3 s 0 106360 800 106480 6 eu2_instruction[27]
port 560 nsew signal output
rlabel metal3 s 0 106904 800 107024 6 eu2_instruction[28]
port 561 nsew signal output
rlabel metal3 s 0 107448 800 107568 6 eu2_instruction[29]
port 562 nsew signal output
rlabel metal3 s 0 92760 800 92880 6 eu2_instruction[2]
port 563 nsew signal output
rlabel metal3 s 0 107992 800 108112 6 eu2_instruction[30]
port 564 nsew signal output
rlabel metal3 s 0 108536 800 108656 6 eu2_instruction[31]
port 565 nsew signal output
rlabel metal3 s 0 109080 800 109200 6 eu2_instruction[32]
port 566 nsew signal output
rlabel metal3 s 0 109624 800 109744 6 eu2_instruction[33]
port 567 nsew signal output
rlabel metal3 s 0 110168 800 110288 6 eu2_instruction[34]
port 568 nsew signal output
rlabel metal3 s 0 110712 800 110832 6 eu2_instruction[35]
port 569 nsew signal output
rlabel metal3 s 0 111256 800 111376 6 eu2_instruction[36]
port 570 nsew signal output
rlabel metal3 s 0 111800 800 111920 6 eu2_instruction[37]
port 571 nsew signal output
rlabel metal3 s 0 112344 800 112464 6 eu2_instruction[38]
port 572 nsew signal output
rlabel metal3 s 0 112888 800 113008 6 eu2_instruction[39]
port 573 nsew signal output
rlabel metal3 s 0 93304 800 93424 6 eu2_instruction[3]
port 574 nsew signal output
rlabel metal3 s 0 113432 800 113552 6 eu2_instruction[40]
port 575 nsew signal output
rlabel metal3 s 0 113976 800 114096 6 eu2_instruction[41]
port 576 nsew signal output
rlabel metal3 s 0 93848 800 93968 6 eu2_instruction[4]
port 577 nsew signal output
rlabel metal3 s 0 94392 800 94512 6 eu2_instruction[5]
port 578 nsew signal output
rlabel metal3 s 0 94936 800 95056 6 eu2_instruction[6]
port 579 nsew signal output
rlabel metal3 s 0 95480 800 95600 6 eu2_instruction[7]
port 580 nsew signal output
rlabel metal3 s 0 96024 800 96144 6 eu2_instruction[8]
port 581 nsew signal output
rlabel metal3 s 0 96568 800 96688 6 eu2_instruction[9]
port 582 nsew signal output
rlabel metal2 s 434442 169200 434498 170000 6 int_return0
port 583 nsew signal input
rlabel metal3 s 439200 150968 440000 151088 6 int_return1
port 584 nsew signal input
rlabel metal3 s 0 149880 800 150000 6 int_return2
port 585 nsew signal input
rlabel metal2 s 232134 0 232190 800 6 io_in[0]
port 586 nsew signal input
rlabel metal2 s 249614 0 249670 800 6 io_in[10]
port 587 nsew signal input
rlabel metal2 s 251362 0 251418 800 6 io_in[11]
port 588 nsew signal input
rlabel metal2 s 253110 0 253166 800 6 io_in[12]
port 589 nsew signal input
rlabel metal2 s 254858 0 254914 800 6 io_in[13]
port 590 nsew signal input
rlabel metal2 s 256606 0 256662 800 6 io_in[14]
port 591 nsew signal input
rlabel metal2 s 258354 0 258410 800 6 io_in[15]
port 592 nsew signal input
rlabel metal2 s 260102 0 260158 800 6 io_in[16]
port 593 nsew signal input
rlabel metal2 s 261850 0 261906 800 6 io_in[17]
port 594 nsew signal input
rlabel metal2 s 263598 0 263654 800 6 io_in[18]
port 595 nsew signal input
rlabel metal2 s 265346 0 265402 800 6 io_in[19]
port 596 nsew signal input
rlabel metal2 s 233882 0 233938 800 6 io_in[1]
port 597 nsew signal input
rlabel metal2 s 267094 0 267150 800 6 io_in[20]
port 598 nsew signal input
rlabel metal2 s 268842 0 268898 800 6 io_in[21]
port 599 nsew signal input
rlabel metal2 s 270590 0 270646 800 6 io_in[22]
port 600 nsew signal input
rlabel metal2 s 272338 0 272394 800 6 io_in[23]
port 601 nsew signal input
rlabel metal2 s 274086 0 274142 800 6 io_in[24]
port 602 nsew signal input
rlabel metal2 s 275834 0 275890 800 6 io_in[25]
port 603 nsew signal input
rlabel metal2 s 277582 0 277638 800 6 io_in[26]
port 604 nsew signal input
rlabel metal2 s 279330 0 279386 800 6 io_in[27]
port 605 nsew signal input
rlabel metal2 s 281078 0 281134 800 6 io_in[28]
port 606 nsew signal input
rlabel metal2 s 282826 0 282882 800 6 io_in[29]
port 607 nsew signal input
rlabel metal2 s 235630 0 235686 800 6 io_in[2]
port 608 nsew signal input
rlabel metal2 s 284574 0 284630 800 6 io_in[30]
port 609 nsew signal input
rlabel metal2 s 286322 0 286378 800 6 io_in[31]
port 610 nsew signal input
rlabel metal2 s 288070 0 288126 800 6 io_in[32]
port 611 nsew signal input
rlabel metal2 s 289818 0 289874 800 6 io_in[33]
port 612 nsew signal input
rlabel metal2 s 291566 0 291622 800 6 io_in[34]
port 613 nsew signal input
rlabel metal2 s 293314 0 293370 800 6 io_in[35]
port 614 nsew signal input
rlabel metal2 s 237378 0 237434 800 6 io_in[3]
port 615 nsew signal input
rlabel metal2 s 239126 0 239182 800 6 io_in[4]
port 616 nsew signal input
rlabel metal2 s 240874 0 240930 800 6 io_in[5]
port 617 nsew signal input
rlabel metal2 s 242622 0 242678 800 6 io_in[6]
port 618 nsew signal input
rlabel metal2 s 244370 0 244426 800 6 io_in[7]
port 619 nsew signal input
rlabel metal2 s 246118 0 246174 800 6 io_in[8]
port 620 nsew signal input
rlabel metal2 s 247866 0 247922 800 6 io_in[9]
port 621 nsew signal input
rlabel metal2 s 295062 0 295118 800 6 io_oeb[0]
port 622 nsew signal output
rlabel metal2 s 312542 0 312598 800 6 io_oeb[10]
port 623 nsew signal output
rlabel metal2 s 314290 0 314346 800 6 io_oeb[11]
port 624 nsew signal output
rlabel metal2 s 316038 0 316094 800 6 io_oeb[12]
port 625 nsew signal output
rlabel metal2 s 317786 0 317842 800 6 io_oeb[13]
port 626 nsew signal output
rlabel metal2 s 319534 0 319590 800 6 io_oeb[14]
port 627 nsew signal output
rlabel metal2 s 321282 0 321338 800 6 io_oeb[15]
port 628 nsew signal output
rlabel metal2 s 323030 0 323086 800 6 io_oeb[16]
port 629 nsew signal output
rlabel metal2 s 324778 0 324834 800 6 io_oeb[17]
port 630 nsew signal output
rlabel metal2 s 326526 0 326582 800 6 io_oeb[18]
port 631 nsew signal output
rlabel metal2 s 328274 0 328330 800 6 io_oeb[19]
port 632 nsew signal output
rlabel metal2 s 296810 0 296866 800 6 io_oeb[1]
port 633 nsew signal output
rlabel metal2 s 330022 0 330078 800 6 io_oeb[20]
port 634 nsew signal output
rlabel metal2 s 331770 0 331826 800 6 io_oeb[21]
port 635 nsew signal output
rlabel metal2 s 333518 0 333574 800 6 io_oeb[22]
port 636 nsew signal output
rlabel metal2 s 335266 0 335322 800 6 io_oeb[23]
port 637 nsew signal output
rlabel metal2 s 337014 0 337070 800 6 io_oeb[24]
port 638 nsew signal output
rlabel metal2 s 338762 0 338818 800 6 io_oeb[25]
port 639 nsew signal output
rlabel metal2 s 340510 0 340566 800 6 io_oeb[26]
port 640 nsew signal output
rlabel metal2 s 342258 0 342314 800 6 io_oeb[27]
port 641 nsew signal output
rlabel metal2 s 344006 0 344062 800 6 io_oeb[28]
port 642 nsew signal output
rlabel metal2 s 345754 0 345810 800 6 io_oeb[29]
port 643 nsew signal output
rlabel metal2 s 298558 0 298614 800 6 io_oeb[2]
port 644 nsew signal output
rlabel metal2 s 347502 0 347558 800 6 io_oeb[30]
port 645 nsew signal output
rlabel metal2 s 349250 0 349306 800 6 io_oeb[31]
port 646 nsew signal output
rlabel metal2 s 350998 0 351054 800 6 io_oeb[32]
port 647 nsew signal output
rlabel metal2 s 352746 0 352802 800 6 io_oeb[33]
port 648 nsew signal output
rlabel metal2 s 354494 0 354550 800 6 io_oeb[34]
port 649 nsew signal output
rlabel metal2 s 356242 0 356298 800 6 io_oeb[35]
port 650 nsew signal output
rlabel metal2 s 300306 0 300362 800 6 io_oeb[3]
port 651 nsew signal output
rlabel metal2 s 302054 0 302110 800 6 io_oeb[4]
port 652 nsew signal output
rlabel metal2 s 303802 0 303858 800 6 io_oeb[5]
port 653 nsew signal output
rlabel metal2 s 305550 0 305606 800 6 io_oeb[6]
port 654 nsew signal output
rlabel metal2 s 307298 0 307354 800 6 io_oeb[7]
port 655 nsew signal output
rlabel metal2 s 309046 0 309102 800 6 io_oeb[8]
port 656 nsew signal output
rlabel metal2 s 310794 0 310850 800 6 io_oeb[9]
port 657 nsew signal output
rlabel metal2 s 357990 0 358046 800 6 io_out[0]
port 658 nsew signal output
rlabel metal2 s 375470 0 375526 800 6 io_out[10]
port 659 nsew signal output
rlabel metal2 s 377218 0 377274 800 6 io_out[11]
port 660 nsew signal output
rlabel metal2 s 378966 0 379022 800 6 io_out[12]
port 661 nsew signal output
rlabel metal2 s 380714 0 380770 800 6 io_out[13]
port 662 nsew signal output
rlabel metal2 s 382462 0 382518 800 6 io_out[14]
port 663 nsew signal output
rlabel metal2 s 384210 0 384266 800 6 io_out[15]
port 664 nsew signal output
rlabel metal2 s 385958 0 386014 800 6 io_out[16]
port 665 nsew signal output
rlabel metal2 s 387706 0 387762 800 6 io_out[17]
port 666 nsew signal output
rlabel metal2 s 389454 0 389510 800 6 io_out[18]
port 667 nsew signal output
rlabel metal2 s 391202 0 391258 800 6 io_out[19]
port 668 nsew signal output
rlabel metal2 s 359738 0 359794 800 6 io_out[1]
port 669 nsew signal output
rlabel metal2 s 392950 0 393006 800 6 io_out[20]
port 670 nsew signal output
rlabel metal2 s 394698 0 394754 800 6 io_out[21]
port 671 nsew signal output
rlabel metal2 s 396446 0 396502 800 6 io_out[22]
port 672 nsew signal output
rlabel metal2 s 398194 0 398250 800 6 io_out[23]
port 673 nsew signal output
rlabel metal2 s 399942 0 399998 800 6 io_out[24]
port 674 nsew signal output
rlabel metal2 s 401690 0 401746 800 6 io_out[25]
port 675 nsew signal output
rlabel metal2 s 403438 0 403494 800 6 io_out[26]
port 676 nsew signal output
rlabel metal2 s 405186 0 405242 800 6 io_out[27]
port 677 nsew signal output
rlabel metal2 s 406934 0 406990 800 6 io_out[28]
port 678 nsew signal output
rlabel metal2 s 408682 0 408738 800 6 io_out[29]
port 679 nsew signal output
rlabel metal2 s 361486 0 361542 800 6 io_out[2]
port 680 nsew signal output
rlabel metal2 s 410430 0 410486 800 6 io_out[30]
port 681 nsew signal output
rlabel metal2 s 412178 0 412234 800 6 io_out[31]
port 682 nsew signal output
rlabel metal2 s 413926 0 413982 800 6 io_out[32]
port 683 nsew signal output
rlabel metal2 s 415674 0 415730 800 6 io_out[33]
port 684 nsew signal output
rlabel metal2 s 417422 0 417478 800 6 io_out[34]
port 685 nsew signal output
rlabel metal2 s 419170 0 419226 800 6 io_out[35]
port 686 nsew signal output
rlabel metal2 s 363234 0 363290 800 6 io_out[3]
port 687 nsew signal output
rlabel metal2 s 364982 0 365038 800 6 io_out[4]
port 688 nsew signal output
rlabel metal2 s 366730 0 366786 800 6 io_out[5]
port 689 nsew signal output
rlabel metal2 s 368478 0 368534 800 6 io_out[6]
port 690 nsew signal output
rlabel metal2 s 370226 0 370282 800 6 io_out[7]
port 691 nsew signal output
rlabel metal2 s 371974 0 372030 800 6 io_out[8]
port 692 nsew signal output
rlabel metal2 s 373722 0 373778 800 6 io_out[9]
port 693 nsew signal output
rlabel metal2 s 284666 169200 284722 170000 6 is_load0
port 694 nsew signal input
rlabel metal3 s 439200 70456 440000 70576 6 is_load1
port 695 nsew signal input
rlabel metal3 s 0 69368 800 69488 6 is_load2
port 696 nsew signal input
rlabel metal2 s 285678 169200 285734 170000 6 is_store0
port 697 nsew signal input
rlabel metal3 s 439200 71000 440000 71120 6 is_store1
port 698 nsew signal input
rlabel metal3 s 0 69912 800 70032 6 is_store2
port 699 nsew signal input
rlabel metal2 s 252282 169200 252338 170000 6 loadstore_address0[0]
port 700 nsew signal input
rlabel metal2 s 262402 169200 262458 170000 6 loadstore_address0[10]
port 701 nsew signal input
rlabel metal2 s 263414 169200 263470 170000 6 loadstore_address0[11]
port 702 nsew signal input
rlabel metal2 s 264426 169200 264482 170000 6 loadstore_address0[12]
port 703 nsew signal input
rlabel metal2 s 265438 169200 265494 170000 6 loadstore_address0[13]
port 704 nsew signal input
rlabel metal2 s 266450 169200 266506 170000 6 loadstore_address0[14]
port 705 nsew signal input
rlabel metal2 s 267462 169200 267518 170000 6 loadstore_address0[15]
port 706 nsew signal input
rlabel metal2 s 268474 169200 268530 170000 6 loadstore_address0[16]
port 707 nsew signal input
rlabel metal2 s 269486 169200 269542 170000 6 loadstore_address0[17]
port 708 nsew signal input
rlabel metal2 s 270498 169200 270554 170000 6 loadstore_address0[18]
port 709 nsew signal input
rlabel metal2 s 271510 169200 271566 170000 6 loadstore_address0[19]
port 710 nsew signal input
rlabel metal2 s 253294 169200 253350 170000 6 loadstore_address0[1]
port 711 nsew signal input
rlabel metal2 s 272522 169200 272578 170000 6 loadstore_address0[20]
port 712 nsew signal input
rlabel metal2 s 273534 169200 273590 170000 6 loadstore_address0[21]
port 713 nsew signal input
rlabel metal2 s 274546 169200 274602 170000 6 loadstore_address0[22]
port 714 nsew signal input
rlabel metal2 s 275558 169200 275614 170000 6 loadstore_address0[23]
port 715 nsew signal input
rlabel metal2 s 276570 169200 276626 170000 6 loadstore_address0[24]
port 716 nsew signal input
rlabel metal2 s 277582 169200 277638 170000 6 loadstore_address0[25]
port 717 nsew signal input
rlabel metal2 s 278594 169200 278650 170000 6 loadstore_address0[26]
port 718 nsew signal input
rlabel metal2 s 279606 169200 279662 170000 6 loadstore_address0[27]
port 719 nsew signal input
rlabel metal2 s 280618 169200 280674 170000 6 loadstore_address0[28]
port 720 nsew signal input
rlabel metal2 s 281630 169200 281686 170000 6 loadstore_address0[29]
port 721 nsew signal input
rlabel metal2 s 254306 169200 254362 170000 6 loadstore_address0[2]
port 722 nsew signal input
rlabel metal2 s 282642 169200 282698 170000 6 loadstore_address0[30]
port 723 nsew signal input
rlabel metal2 s 283654 169200 283710 170000 6 loadstore_address0[31]
port 724 nsew signal input
rlabel metal2 s 255318 169200 255374 170000 6 loadstore_address0[3]
port 725 nsew signal input
rlabel metal2 s 256330 169200 256386 170000 6 loadstore_address0[4]
port 726 nsew signal input
rlabel metal2 s 257342 169200 257398 170000 6 loadstore_address0[5]
port 727 nsew signal input
rlabel metal2 s 258354 169200 258410 170000 6 loadstore_address0[6]
port 728 nsew signal input
rlabel metal2 s 259366 169200 259422 170000 6 loadstore_address0[7]
port 729 nsew signal input
rlabel metal2 s 260378 169200 260434 170000 6 loadstore_address0[8]
port 730 nsew signal input
rlabel metal2 s 261390 169200 261446 170000 6 loadstore_address0[9]
port 731 nsew signal input
rlabel metal3 s 439200 53048 440000 53168 6 loadstore_address1[0]
port 732 nsew signal input
rlabel metal3 s 439200 58488 440000 58608 6 loadstore_address1[10]
port 733 nsew signal input
rlabel metal3 s 439200 59032 440000 59152 6 loadstore_address1[11]
port 734 nsew signal input
rlabel metal3 s 439200 59576 440000 59696 6 loadstore_address1[12]
port 735 nsew signal input
rlabel metal3 s 439200 60120 440000 60240 6 loadstore_address1[13]
port 736 nsew signal input
rlabel metal3 s 439200 60664 440000 60784 6 loadstore_address1[14]
port 737 nsew signal input
rlabel metal3 s 439200 61208 440000 61328 6 loadstore_address1[15]
port 738 nsew signal input
rlabel metal3 s 439200 61752 440000 61872 6 loadstore_address1[16]
port 739 nsew signal input
rlabel metal3 s 439200 62296 440000 62416 6 loadstore_address1[17]
port 740 nsew signal input
rlabel metal3 s 439200 62840 440000 62960 6 loadstore_address1[18]
port 741 nsew signal input
rlabel metal3 s 439200 63384 440000 63504 6 loadstore_address1[19]
port 742 nsew signal input
rlabel metal3 s 439200 53592 440000 53712 6 loadstore_address1[1]
port 743 nsew signal input
rlabel metal3 s 439200 63928 440000 64048 6 loadstore_address1[20]
port 744 nsew signal input
rlabel metal3 s 439200 64472 440000 64592 6 loadstore_address1[21]
port 745 nsew signal input
rlabel metal3 s 439200 65016 440000 65136 6 loadstore_address1[22]
port 746 nsew signal input
rlabel metal3 s 439200 65560 440000 65680 6 loadstore_address1[23]
port 747 nsew signal input
rlabel metal3 s 439200 66104 440000 66224 6 loadstore_address1[24]
port 748 nsew signal input
rlabel metal3 s 439200 66648 440000 66768 6 loadstore_address1[25]
port 749 nsew signal input
rlabel metal3 s 439200 67192 440000 67312 6 loadstore_address1[26]
port 750 nsew signal input
rlabel metal3 s 439200 67736 440000 67856 6 loadstore_address1[27]
port 751 nsew signal input
rlabel metal3 s 439200 68280 440000 68400 6 loadstore_address1[28]
port 752 nsew signal input
rlabel metal3 s 439200 68824 440000 68944 6 loadstore_address1[29]
port 753 nsew signal input
rlabel metal3 s 439200 54136 440000 54256 6 loadstore_address1[2]
port 754 nsew signal input
rlabel metal3 s 439200 69368 440000 69488 6 loadstore_address1[30]
port 755 nsew signal input
rlabel metal3 s 439200 69912 440000 70032 6 loadstore_address1[31]
port 756 nsew signal input
rlabel metal3 s 439200 54680 440000 54800 6 loadstore_address1[3]
port 757 nsew signal input
rlabel metal3 s 439200 55224 440000 55344 6 loadstore_address1[4]
port 758 nsew signal input
rlabel metal3 s 439200 55768 440000 55888 6 loadstore_address1[5]
port 759 nsew signal input
rlabel metal3 s 439200 56312 440000 56432 6 loadstore_address1[6]
port 760 nsew signal input
rlabel metal3 s 439200 56856 440000 56976 6 loadstore_address1[7]
port 761 nsew signal input
rlabel metal3 s 439200 57400 440000 57520 6 loadstore_address1[8]
port 762 nsew signal input
rlabel metal3 s 439200 57944 440000 58064 6 loadstore_address1[9]
port 763 nsew signal input
rlabel metal3 s 0 51960 800 52080 6 loadstore_address2[0]
port 764 nsew signal input
rlabel metal3 s 0 57400 800 57520 6 loadstore_address2[10]
port 765 nsew signal input
rlabel metal3 s 0 57944 800 58064 6 loadstore_address2[11]
port 766 nsew signal input
rlabel metal3 s 0 58488 800 58608 6 loadstore_address2[12]
port 767 nsew signal input
rlabel metal3 s 0 59032 800 59152 6 loadstore_address2[13]
port 768 nsew signal input
rlabel metal3 s 0 59576 800 59696 6 loadstore_address2[14]
port 769 nsew signal input
rlabel metal3 s 0 60120 800 60240 6 loadstore_address2[15]
port 770 nsew signal input
rlabel metal3 s 0 60664 800 60784 6 loadstore_address2[16]
port 771 nsew signal input
rlabel metal3 s 0 61208 800 61328 6 loadstore_address2[17]
port 772 nsew signal input
rlabel metal3 s 0 61752 800 61872 6 loadstore_address2[18]
port 773 nsew signal input
rlabel metal3 s 0 62296 800 62416 6 loadstore_address2[19]
port 774 nsew signal input
rlabel metal3 s 0 52504 800 52624 6 loadstore_address2[1]
port 775 nsew signal input
rlabel metal3 s 0 62840 800 62960 6 loadstore_address2[20]
port 776 nsew signal input
rlabel metal3 s 0 63384 800 63504 6 loadstore_address2[21]
port 777 nsew signal input
rlabel metal3 s 0 63928 800 64048 6 loadstore_address2[22]
port 778 nsew signal input
rlabel metal3 s 0 64472 800 64592 6 loadstore_address2[23]
port 779 nsew signal input
rlabel metal3 s 0 65016 800 65136 6 loadstore_address2[24]
port 780 nsew signal input
rlabel metal3 s 0 65560 800 65680 6 loadstore_address2[25]
port 781 nsew signal input
rlabel metal3 s 0 66104 800 66224 6 loadstore_address2[26]
port 782 nsew signal input
rlabel metal3 s 0 66648 800 66768 6 loadstore_address2[27]
port 783 nsew signal input
rlabel metal3 s 0 67192 800 67312 6 loadstore_address2[28]
port 784 nsew signal input
rlabel metal3 s 0 67736 800 67856 6 loadstore_address2[29]
port 785 nsew signal input
rlabel metal3 s 0 53048 800 53168 6 loadstore_address2[2]
port 786 nsew signal input
rlabel metal3 s 0 68280 800 68400 6 loadstore_address2[30]
port 787 nsew signal input
rlabel metal3 s 0 68824 800 68944 6 loadstore_address2[31]
port 788 nsew signal input
rlabel metal3 s 0 53592 800 53712 6 loadstore_address2[3]
port 789 nsew signal input
rlabel metal3 s 0 54136 800 54256 6 loadstore_address2[4]
port 790 nsew signal input
rlabel metal3 s 0 54680 800 54800 6 loadstore_address2[5]
port 791 nsew signal input
rlabel metal3 s 0 55224 800 55344 6 loadstore_address2[6]
port 792 nsew signal input
rlabel metal3 s 0 55768 800 55888 6 loadstore_address2[7]
port 793 nsew signal input
rlabel metal3 s 0 56312 800 56432 6 loadstore_address2[8]
port 794 nsew signal input
rlabel metal3 s 0 56856 800 56976 6 loadstore_address2[9]
port 795 nsew signal input
rlabel metal2 s 289726 169200 289782 170000 6 loadstore_dest0[0]
port 796 nsew signal input
rlabel metal2 s 290738 169200 290794 170000 6 loadstore_dest0[1]
port 797 nsew signal input
rlabel metal2 s 291750 169200 291806 170000 6 loadstore_dest0[2]
port 798 nsew signal input
rlabel metal2 s 292762 169200 292818 170000 6 loadstore_dest0[3]
port 799 nsew signal input
rlabel metal2 s 293774 169200 293830 170000 6 loadstore_dest0[4]
port 800 nsew signal input
rlabel metal2 s 294786 169200 294842 170000 6 loadstore_dest0[5]
port 801 nsew signal input
rlabel metal3 s 439200 73176 440000 73296 6 loadstore_dest1[0]
port 802 nsew signal input
rlabel metal3 s 439200 73720 440000 73840 6 loadstore_dest1[1]
port 803 nsew signal input
rlabel metal3 s 439200 74264 440000 74384 6 loadstore_dest1[2]
port 804 nsew signal input
rlabel metal3 s 439200 74808 440000 74928 6 loadstore_dest1[3]
port 805 nsew signal input
rlabel metal3 s 439200 75352 440000 75472 6 loadstore_dest1[4]
port 806 nsew signal input
rlabel metal3 s 439200 75896 440000 76016 6 loadstore_dest1[5]
port 807 nsew signal input
rlabel metal3 s 0 72088 800 72208 6 loadstore_dest2[0]
port 808 nsew signal input
rlabel metal3 s 0 72632 800 72752 6 loadstore_dest2[1]
port 809 nsew signal input
rlabel metal3 s 0 73176 800 73296 6 loadstore_dest2[2]
port 810 nsew signal input
rlabel metal3 s 0 73720 800 73840 6 loadstore_dest2[3]
port 811 nsew signal input
rlabel metal3 s 0 74264 800 74384 6 loadstore_dest2[4]
port 812 nsew signal input
rlabel metal3 s 0 74808 800 74928 6 loadstore_dest2[5]
port 813 nsew signal input
rlabel metal2 s 287702 169200 287758 170000 6 loadstore_size0[0]
port 814 nsew signal input
rlabel metal2 s 288714 169200 288770 170000 6 loadstore_size0[1]
port 815 nsew signal input
rlabel metal3 s 439200 72088 440000 72208 6 loadstore_size1[0]
port 816 nsew signal input
rlabel metal3 s 439200 72632 440000 72752 6 loadstore_size1[1]
port 817 nsew signal input
rlabel metal3 s 0 71000 800 71120 6 loadstore_size2[0]
port 818 nsew signal input
rlabel metal3 s 0 71544 800 71664 6 loadstore_size2[1]
port 819 nsew signal input
rlabel metal2 s 296810 169200 296866 170000 6 new_PC0[0]
port 820 nsew signal input
rlabel metal2 s 306930 169200 306986 170000 6 new_PC0[10]
port 821 nsew signal input
rlabel metal2 s 307942 169200 307998 170000 6 new_PC0[11]
port 822 nsew signal input
rlabel metal2 s 308954 169200 309010 170000 6 new_PC0[12]
port 823 nsew signal input
rlabel metal2 s 309966 169200 310022 170000 6 new_PC0[13]
port 824 nsew signal input
rlabel metal2 s 310978 169200 311034 170000 6 new_PC0[14]
port 825 nsew signal input
rlabel metal2 s 311990 169200 312046 170000 6 new_PC0[15]
port 826 nsew signal input
rlabel metal2 s 313002 169200 313058 170000 6 new_PC0[16]
port 827 nsew signal input
rlabel metal2 s 314014 169200 314070 170000 6 new_PC0[17]
port 828 nsew signal input
rlabel metal2 s 315026 169200 315082 170000 6 new_PC0[18]
port 829 nsew signal input
rlabel metal2 s 316038 169200 316094 170000 6 new_PC0[19]
port 830 nsew signal input
rlabel metal2 s 297822 169200 297878 170000 6 new_PC0[1]
port 831 nsew signal input
rlabel metal2 s 317050 169200 317106 170000 6 new_PC0[20]
port 832 nsew signal input
rlabel metal2 s 318062 169200 318118 170000 6 new_PC0[21]
port 833 nsew signal input
rlabel metal2 s 319074 169200 319130 170000 6 new_PC0[22]
port 834 nsew signal input
rlabel metal2 s 320086 169200 320142 170000 6 new_PC0[23]
port 835 nsew signal input
rlabel metal2 s 321098 169200 321154 170000 6 new_PC0[24]
port 836 nsew signal input
rlabel metal2 s 322110 169200 322166 170000 6 new_PC0[25]
port 837 nsew signal input
rlabel metal2 s 323122 169200 323178 170000 6 new_PC0[26]
port 838 nsew signal input
rlabel metal2 s 324134 169200 324190 170000 6 new_PC0[27]
port 839 nsew signal input
rlabel metal2 s 298834 169200 298890 170000 6 new_PC0[2]
port 840 nsew signal input
rlabel metal2 s 299846 169200 299902 170000 6 new_PC0[3]
port 841 nsew signal input
rlabel metal2 s 300858 169200 300914 170000 6 new_PC0[4]
port 842 nsew signal input
rlabel metal2 s 301870 169200 301926 170000 6 new_PC0[5]
port 843 nsew signal input
rlabel metal2 s 302882 169200 302938 170000 6 new_PC0[6]
port 844 nsew signal input
rlabel metal2 s 303894 169200 303950 170000 6 new_PC0[7]
port 845 nsew signal input
rlabel metal2 s 304906 169200 304962 170000 6 new_PC0[8]
port 846 nsew signal input
rlabel metal2 s 305918 169200 305974 170000 6 new_PC0[9]
port 847 nsew signal input
rlabel metal3 s 439200 76984 440000 77104 6 new_PC1[0]
port 848 nsew signal input
rlabel metal3 s 439200 82424 440000 82544 6 new_PC1[10]
port 849 nsew signal input
rlabel metal3 s 439200 82968 440000 83088 6 new_PC1[11]
port 850 nsew signal input
rlabel metal3 s 439200 83512 440000 83632 6 new_PC1[12]
port 851 nsew signal input
rlabel metal3 s 439200 84056 440000 84176 6 new_PC1[13]
port 852 nsew signal input
rlabel metal3 s 439200 84600 440000 84720 6 new_PC1[14]
port 853 nsew signal input
rlabel metal3 s 439200 85144 440000 85264 6 new_PC1[15]
port 854 nsew signal input
rlabel metal3 s 439200 85688 440000 85808 6 new_PC1[16]
port 855 nsew signal input
rlabel metal3 s 439200 86232 440000 86352 6 new_PC1[17]
port 856 nsew signal input
rlabel metal3 s 439200 86776 440000 86896 6 new_PC1[18]
port 857 nsew signal input
rlabel metal3 s 439200 87320 440000 87440 6 new_PC1[19]
port 858 nsew signal input
rlabel metal3 s 439200 77528 440000 77648 6 new_PC1[1]
port 859 nsew signal input
rlabel metal3 s 439200 87864 440000 87984 6 new_PC1[20]
port 860 nsew signal input
rlabel metal3 s 439200 88408 440000 88528 6 new_PC1[21]
port 861 nsew signal input
rlabel metal3 s 439200 88952 440000 89072 6 new_PC1[22]
port 862 nsew signal input
rlabel metal3 s 439200 89496 440000 89616 6 new_PC1[23]
port 863 nsew signal input
rlabel metal3 s 439200 90040 440000 90160 6 new_PC1[24]
port 864 nsew signal input
rlabel metal3 s 439200 90584 440000 90704 6 new_PC1[25]
port 865 nsew signal input
rlabel metal3 s 439200 91128 440000 91248 6 new_PC1[26]
port 866 nsew signal input
rlabel metal3 s 439200 91672 440000 91792 6 new_PC1[27]
port 867 nsew signal input
rlabel metal3 s 439200 78072 440000 78192 6 new_PC1[2]
port 868 nsew signal input
rlabel metal3 s 439200 78616 440000 78736 6 new_PC1[3]
port 869 nsew signal input
rlabel metal3 s 439200 79160 440000 79280 6 new_PC1[4]
port 870 nsew signal input
rlabel metal3 s 439200 79704 440000 79824 6 new_PC1[5]
port 871 nsew signal input
rlabel metal3 s 439200 80248 440000 80368 6 new_PC1[6]
port 872 nsew signal input
rlabel metal3 s 439200 80792 440000 80912 6 new_PC1[7]
port 873 nsew signal input
rlabel metal3 s 439200 81336 440000 81456 6 new_PC1[8]
port 874 nsew signal input
rlabel metal3 s 439200 81880 440000 82000 6 new_PC1[9]
port 875 nsew signal input
rlabel metal3 s 0 75896 800 76016 6 new_PC2[0]
port 876 nsew signal input
rlabel metal3 s 0 81336 800 81456 6 new_PC2[10]
port 877 nsew signal input
rlabel metal3 s 0 81880 800 82000 6 new_PC2[11]
port 878 nsew signal input
rlabel metal3 s 0 82424 800 82544 6 new_PC2[12]
port 879 nsew signal input
rlabel metal3 s 0 82968 800 83088 6 new_PC2[13]
port 880 nsew signal input
rlabel metal3 s 0 83512 800 83632 6 new_PC2[14]
port 881 nsew signal input
rlabel metal3 s 0 84056 800 84176 6 new_PC2[15]
port 882 nsew signal input
rlabel metal3 s 0 84600 800 84720 6 new_PC2[16]
port 883 nsew signal input
rlabel metal3 s 0 85144 800 85264 6 new_PC2[17]
port 884 nsew signal input
rlabel metal3 s 0 85688 800 85808 6 new_PC2[18]
port 885 nsew signal input
rlabel metal3 s 0 86232 800 86352 6 new_PC2[19]
port 886 nsew signal input
rlabel metal3 s 0 76440 800 76560 6 new_PC2[1]
port 887 nsew signal input
rlabel metal3 s 0 86776 800 86896 6 new_PC2[20]
port 888 nsew signal input
rlabel metal3 s 0 87320 800 87440 6 new_PC2[21]
port 889 nsew signal input
rlabel metal3 s 0 87864 800 87984 6 new_PC2[22]
port 890 nsew signal input
rlabel metal3 s 0 88408 800 88528 6 new_PC2[23]
port 891 nsew signal input
rlabel metal3 s 0 88952 800 89072 6 new_PC2[24]
port 892 nsew signal input
rlabel metal3 s 0 89496 800 89616 6 new_PC2[25]
port 893 nsew signal input
rlabel metal3 s 0 90040 800 90160 6 new_PC2[26]
port 894 nsew signal input
rlabel metal3 s 0 90584 800 90704 6 new_PC2[27]
port 895 nsew signal input
rlabel metal3 s 0 76984 800 77104 6 new_PC2[2]
port 896 nsew signal input
rlabel metal3 s 0 77528 800 77648 6 new_PC2[3]
port 897 nsew signal input
rlabel metal3 s 0 78072 800 78192 6 new_PC2[4]
port 898 nsew signal input
rlabel metal3 s 0 78616 800 78736 6 new_PC2[5]
port 899 nsew signal input
rlabel metal3 s 0 79160 800 79280 6 new_PC2[6]
port 900 nsew signal input
rlabel metal3 s 0 79704 800 79824 6 new_PC2[7]
port 901 nsew signal input
rlabel metal3 s 0 80248 800 80368 6 new_PC2[8]
port 902 nsew signal input
rlabel metal3 s 0 80792 800 80912 6 new_PC2[9]
port 903 nsew signal input
rlabel metal2 s 245198 169200 245254 170000 6 pred_idx0[0]
port 904 nsew signal input
rlabel metal2 s 246210 169200 246266 170000 6 pred_idx0[1]
port 905 nsew signal input
rlabel metal2 s 247222 169200 247278 170000 6 pred_idx0[2]
port 906 nsew signal input
rlabel metal3 s 439200 49240 440000 49360 6 pred_idx1[0]
port 907 nsew signal input
rlabel metal3 s 439200 49784 440000 49904 6 pred_idx1[1]
port 908 nsew signal input
rlabel metal3 s 439200 50328 440000 50448 6 pred_idx1[2]
port 909 nsew signal input
rlabel metal3 s 0 48152 800 48272 6 pred_idx2[0]
port 910 nsew signal input
rlabel metal3 s 0 48696 800 48816 6 pred_idx2[1]
port 911 nsew signal input
rlabel metal3 s 0 49240 800 49360 6 pred_idx2[2]
port 912 nsew signal input
rlabel metal2 s 433430 169200 433486 170000 6 pred_val0
port 913 nsew signal output
rlabel metal3 s 439200 150424 440000 150544 6 pred_val1
port 914 nsew signal output
rlabel metal3 s 0 149336 800 149456 6 pred_val2
port 915 nsew signal output
rlabel metal2 s 192574 169200 192630 170000 6 reg1_idx0[0]
port 916 nsew signal input
rlabel metal2 s 193586 169200 193642 170000 6 reg1_idx0[1]
port 917 nsew signal input
rlabel metal2 s 194598 169200 194654 170000 6 reg1_idx0[2]
port 918 nsew signal input
rlabel metal2 s 195610 169200 195666 170000 6 reg1_idx0[3]
port 919 nsew signal input
rlabel metal2 s 196622 169200 196678 170000 6 reg1_idx0[4]
port 920 nsew signal input
rlabel metal2 s 197634 169200 197690 170000 6 reg1_idx0[5]
port 921 nsew signal input
rlabel metal3 s 439200 20952 440000 21072 6 reg1_idx1[0]
port 922 nsew signal input
rlabel metal3 s 439200 21496 440000 21616 6 reg1_idx1[1]
port 923 nsew signal input
rlabel metal3 s 439200 22040 440000 22160 6 reg1_idx1[2]
port 924 nsew signal input
rlabel metal3 s 439200 22584 440000 22704 6 reg1_idx1[3]
port 925 nsew signal input
rlabel metal3 s 439200 23128 440000 23248 6 reg1_idx1[4]
port 926 nsew signal input
rlabel metal3 s 439200 23672 440000 23792 6 reg1_idx1[5]
port 927 nsew signal input
rlabel metal3 s 0 19864 800 19984 6 reg1_idx2[0]
port 928 nsew signal input
rlabel metal3 s 0 20408 800 20528 6 reg1_idx2[1]
port 929 nsew signal input
rlabel metal3 s 0 20952 800 21072 6 reg1_idx2[2]
port 930 nsew signal input
rlabel metal3 s 0 21496 800 21616 6 reg1_idx2[3]
port 931 nsew signal input
rlabel metal3 s 0 22040 800 22160 6 reg1_idx2[4]
port 932 nsew signal input
rlabel metal3 s 0 22584 800 22704 6 reg1_idx2[5]
port 933 nsew signal input
rlabel metal2 s 368662 169200 368718 170000 6 reg1_val0[0]
port 934 nsew signal output
rlabel metal2 s 378782 169200 378838 170000 6 reg1_val0[10]
port 935 nsew signal output
rlabel metal2 s 379794 169200 379850 170000 6 reg1_val0[11]
port 936 nsew signal output
rlabel metal2 s 380806 169200 380862 170000 6 reg1_val0[12]
port 937 nsew signal output
rlabel metal2 s 381818 169200 381874 170000 6 reg1_val0[13]
port 938 nsew signal output
rlabel metal2 s 382830 169200 382886 170000 6 reg1_val0[14]
port 939 nsew signal output
rlabel metal2 s 383842 169200 383898 170000 6 reg1_val0[15]
port 940 nsew signal output
rlabel metal2 s 384854 169200 384910 170000 6 reg1_val0[16]
port 941 nsew signal output
rlabel metal2 s 385866 169200 385922 170000 6 reg1_val0[17]
port 942 nsew signal output
rlabel metal2 s 386878 169200 386934 170000 6 reg1_val0[18]
port 943 nsew signal output
rlabel metal2 s 387890 169200 387946 170000 6 reg1_val0[19]
port 944 nsew signal output
rlabel metal2 s 369674 169200 369730 170000 6 reg1_val0[1]
port 945 nsew signal output
rlabel metal2 s 388902 169200 388958 170000 6 reg1_val0[20]
port 946 nsew signal output
rlabel metal2 s 389914 169200 389970 170000 6 reg1_val0[21]
port 947 nsew signal output
rlabel metal2 s 390926 169200 390982 170000 6 reg1_val0[22]
port 948 nsew signal output
rlabel metal2 s 391938 169200 391994 170000 6 reg1_val0[23]
port 949 nsew signal output
rlabel metal2 s 392950 169200 393006 170000 6 reg1_val0[24]
port 950 nsew signal output
rlabel metal2 s 393962 169200 394018 170000 6 reg1_val0[25]
port 951 nsew signal output
rlabel metal2 s 394974 169200 395030 170000 6 reg1_val0[26]
port 952 nsew signal output
rlabel metal2 s 395986 169200 396042 170000 6 reg1_val0[27]
port 953 nsew signal output
rlabel metal2 s 396998 169200 397054 170000 6 reg1_val0[28]
port 954 nsew signal output
rlabel metal2 s 398010 169200 398066 170000 6 reg1_val0[29]
port 955 nsew signal output
rlabel metal2 s 370686 169200 370742 170000 6 reg1_val0[2]
port 956 nsew signal output
rlabel metal2 s 399022 169200 399078 170000 6 reg1_val0[30]
port 957 nsew signal output
rlabel metal2 s 400034 169200 400090 170000 6 reg1_val0[31]
port 958 nsew signal output
rlabel metal2 s 371698 169200 371754 170000 6 reg1_val0[3]
port 959 nsew signal output
rlabel metal2 s 372710 169200 372766 170000 6 reg1_val0[4]
port 960 nsew signal output
rlabel metal2 s 373722 169200 373778 170000 6 reg1_val0[5]
port 961 nsew signal output
rlabel metal2 s 374734 169200 374790 170000 6 reg1_val0[6]
port 962 nsew signal output
rlabel metal2 s 375746 169200 375802 170000 6 reg1_val0[7]
port 963 nsew signal output
rlabel metal2 s 376758 169200 376814 170000 6 reg1_val0[8]
port 964 nsew signal output
rlabel metal2 s 377770 169200 377826 170000 6 reg1_val0[9]
port 965 nsew signal output
rlabel metal3 s 439200 115608 440000 115728 6 reg1_val1[0]
port 966 nsew signal output
rlabel metal3 s 439200 121048 440000 121168 6 reg1_val1[10]
port 967 nsew signal output
rlabel metal3 s 439200 121592 440000 121712 6 reg1_val1[11]
port 968 nsew signal output
rlabel metal3 s 439200 122136 440000 122256 6 reg1_val1[12]
port 969 nsew signal output
rlabel metal3 s 439200 122680 440000 122800 6 reg1_val1[13]
port 970 nsew signal output
rlabel metal3 s 439200 123224 440000 123344 6 reg1_val1[14]
port 971 nsew signal output
rlabel metal3 s 439200 123768 440000 123888 6 reg1_val1[15]
port 972 nsew signal output
rlabel metal3 s 439200 124312 440000 124432 6 reg1_val1[16]
port 973 nsew signal output
rlabel metal3 s 439200 124856 440000 124976 6 reg1_val1[17]
port 974 nsew signal output
rlabel metal3 s 439200 125400 440000 125520 6 reg1_val1[18]
port 975 nsew signal output
rlabel metal3 s 439200 125944 440000 126064 6 reg1_val1[19]
port 976 nsew signal output
rlabel metal3 s 439200 116152 440000 116272 6 reg1_val1[1]
port 977 nsew signal output
rlabel metal3 s 439200 126488 440000 126608 6 reg1_val1[20]
port 978 nsew signal output
rlabel metal3 s 439200 127032 440000 127152 6 reg1_val1[21]
port 979 nsew signal output
rlabel metal3 s 439200 127576 440000 127696 6 reg1_val1[22]
port 980 nsew signal output
rlabel metal3 s 439200 128120 440000 128240 6 reg1_val1[23]
port 981 nsew signal output
rlabel metal3 s 439200 128664 440000 128784 6 reg1_val1[24]
port 982 nsew signal output
rlabel metal3 s 439200 129208 440000 129328 6 reg1_val1[25]
port 983 nsew signal output
rlabel metal3 s 439200 129752 440000 129872 6 reg1_val1[26]
port 984 nsew signal output
rlabel metal3 s 439200 130296 440000 130416 6 reg1_val1[27]
port 985 nsew signal output
rlabel metal3 s 439200 130840 440000 130960 6 reg1_val1[28]
port 986 nsew signal output
rlabel metal3 s 439200 131384 440000 131504 6 reg1_val1[29]
port 987 nsew signal output
rlabel metal3 s 439200 116696 440000 116816 6 reg1_val1[2]
port 988 nsew signal output
rlabel metal3 s 439200 131928 440000 132048 6 reg1_val1[30]
port 989 nsew signal output
rlabel metal3 s 439200 132472 440000 132592 6 reg1_val1[31]
port 990 nsew signal output
rlabel metal3 s 439200 117240 440000 117360 6 reg1_val1[3]
port 991 nsew signal output
rlabel metal3 s 439200 117784 440000 117904 6 reg1_val1[4]
port 992 nsew signal output
rlabel metal3 s 439200 118328 440000 118448 6 reg1_val1[5]
port 993 nsew signal output
rlabel metal3 s 439200 118872 440000 118992 6 reg1_val1[6]
port 994 nsew signal output
rlabel metal3 s 439200 119416 440000 119536 6 reg1_val1[7]
port 995 nsew signal output
rlabel metal3 s 439200 119960 440000 120080 6 reg1_val1[8]
port 996 nsew signal output
rlabel metal3 s 439200 120504 440000 120624 6 reg1_val1[9]
port 997 nsew signal output
rlabel metal3 s 0 114520 800 114640 6 reg1_val2[0]
port 998 nsew signal output
rlabel metal3 s 0 119960 800 120080 6 reg1_val2[10]
port 999 nsew signal output
rlabel metal3 s 0 120504 800 120624 6 reg1_val2[11]
port 1000 nsew signal output
rlabel metal3 s 0 121048 800 121168 6 reg1_val2[12]
port 1001 nsew signal output
rlabel metal3 s 0 121592 800 121712 6 reg1_val2[13]
port 1002 nsew signal output
rlabel metal3 s 0 122136 800 122256 6 reg1_val2[14]
port 1003 nsew signal output
rlabel metal3 s 0 122680 800 122800 6 reg1_val2[15]
port 1004 nsew signal output
rlabel metal3 s 0 123224 800 123344 6 reg1_val2[16]
port 1005 nsew signal output
rlabel metal3 s 0 123768 800 123888 6 reg1_val2[17]
port 1006 nsew signal output
rlabel metal3 s 0 124312 800 124432 6 reg1_val2[18]
port 1007 nsew signal output
rlabel metal3 s 0 124856 800 124976 6 reg1_val2[19]
port 1008 nsew signal output
rlabel metal3 s 0 115064 800 115184 6 reg1_val2[1]
port 1009 nsew signal output
rlabel metal3 s 0 125400 800 125520 6 reg1_val2[20]
port 1010 nsew signal output
rlabel metal3 s 0 125944 800 126064 6 reg1_val2[21]
port 1011 nsew signal output
rlabel metal3 s 0 126488 800 126608 6 reg1_val2[22]
port 1012 nsew signal output
rlabel metal3 s 0 127032 800 127152 6 reg1_val2[23]
port 1013 nsew signal output
rlabel metal3 s 0 127576 800 127696 6 reg1_val2[24]
port 1014 nsew signal output
rlabel metal3 s 0 128120 800 128240 6 reg1_val2[25]
port 1015 nsew signal output
rlabel metal3 s 0 128664 800 128784 6 reg1_val2[26]
port 1016 nsew signal output
rlabel metal3 s 0 129208 800 129328 6 reg1_val2[27]
port 1017 nsew signal output
rlabel metal3 s 0 129752 800 129872 6 reg1_val2[28]
port 1018 nsew signal output
rlabel metal3 s 0 130296 800 130416 6 reg1_val2[29]
port 1019 nsew signal output
rlabel metal3 s 0 115608 800 115728 6 reg1_val2[2]
port 1020 nsew signal output
rlabel metal3 s 0 130840 800 130960 6 reg1_val2[30]
port 1021 nsew signal output
rlabel metal3 s 0 131384 800 131504 6 reg1_val2[31]
port 1022 nsew signal output
rlabel metal3 s 0 116152 800 116272 6 reg1_val2[3]
port 1023 nsew signal output
rlabel metal3 s 0 116696 800 116816 6 reg1_val2[4]
port 1024 nsew signal output
rlabel metal3 s 0 117240 800 117360 6 reg1_val2[5]
port 1025 nsew signal output
rlabel metal3 s 0 117784 800 117904 6 reg1_val2[6]
port 1026 nsew signal output
rlabel metal3 s 0 118328 800 118448 6 reg1_val2[7]
port 1027 nsew signal output
rlabel metal3 s 0 118872 800 118992 6 reg1_val2[8]
port 1028 nsew signal output
rlabel metal3 s 0 119416 800 119536 6 reg1_val2[9]
port 1029 nsew signal output
rlabel metal2 s 198646 169200 198702 170000 6 reg2_idx0[0]
port 1030 nsew signal input
rlabel metal2 s 199658 169200 199714 170000 6 reg2_idx0[1]
port 1031 nsew signal input
rlabel metal2 s 200670 169200 200726 170000 6 reg2_idx0[2]
port 1032 nsew signal input
rlabel metal2 s 201682 169200 201738 170000 6 reg2_idx0[3]
port 1033 nsew signal input
rlabel metal2 s 202694 169200 202750 170000 6 reg2_idx0[4]
port 1034 nsew signal input
rlabel metal2 s 203706 169200 203762 170000 6 reg2_idx0[5]
port 1035 nsew signal input
rlabel metal3 s 439200 24216 440000 24336 6 reg2_idx1[0]
port 1036 nsew signal input
rlabel metal3 s 439200 24760 440000 24880 6 reg2_idx1[1]
port 1037 nsew signal input
rlabel metal3 s 439200 25304 440000 25424 6 reg2_idx1[2]
port 1038 nsew signal input
rlabel metal3 s 439200 25848 440000 25968 6 reg2_idx1[3]
port 1039 nsew signal input
rlabel metal3 s 439200 26392 440000 26512 6 reg2_idx1[4]
port 1040 nsew signal input
rlabel metal3 s 439200 26936 440000 27056 6 reg2_idx1[5]
port 1041 nsew signal input
rlabel metal3 s 0 23128 800 23248 6 reg2_idx2[0]
port 1042 nsew signal input
rlabel metal3 s 0 23672 800 23792 6 reg2_idx2[1]
port 1043 nsew signal input
rlabel metal3 s 0 24216 800 24336 6 reg2_idx2[2]
port 1044 nsew signal input
rlabel metal3 s 0 24760 800 24880 6 reg2_idx2[3]
port 1045 nsew signal input
rlabel metal3 s 0 25304 800 25424 6 reg2_idx2[4]
port 1046 nsew signal input
rlabel metal3 s 0 25848 800 25968 6 reg2_idx2[5]
port 1047 nsew signal input
rlabel metal2 s 401046 169200 401102 170000 6 reg2_val0[0]
port 1048 nsew signal output
rlabel metal2 s 411166 169200 411222 170000 6 reg2_val0[10]
port 1049 nsew signal output
rlabel metal2 s 412178 169200 412234 170000 6 reg2_val0[11]
port 1050 nsew signal output
rlabel metal2 s 413190 169200 413246 170000 6 reg2_val0[12]
port 1051 nsew signal output
rlabel metal2 s 414202 169200 414258 170000 6 reg2_val0[13]
port 1052 nsew signal output
rlabel metal2 s 415214 169200 415270 170000 6 reg2_val0[14]
port 1053 nsew signal output
rlabel metal2 s 416226 169200 416282 170000 6 reg2_val0[15]
port 1054 nsew signal output
rlabel metal2 s 417238 169200 417294 170000 6 reg2_val0[16]
port 1055 nsew signal output
rlabel metal2 s 418250 169200 418306 170000 6 reg2_val0[17]
port 1056 nsew signal output
rlabel metal2 s 419262 169200 419318 170000 6 reg2_val0[18]
port 1057 nsew signal output
rlabel metal2 s 420274 169200 420330 170000 6 reg2_val0[19]
port 1058 nsew signal output
rlabel metal2 s 402058 169200 402114 170000 6 reg2_val0[1]
port 1059 nsew signal output
rlabel metal2 s 421286 169200 421342 170000 6 reg2_val0[20]
port 1060 nsew signal output
rlabel metal2 s 422298 169200 422354 170000 6 reg2_val0[21]
port 1061 nsew signal output
rlabel metal2 s 423310 169200 423366 170000 6 reg2_val0[22]
port 1062 nsew signal output
rlabel metal2 s 424322 169200 424378 170000 6 reg2_val0[23]
port 1063 nsew signal output
rlabel metal2 s 425334 169200 425390 170000 6 reg2_val0[24]
port 1064 nsew signal output
rlabel metal2 s 426346 169200 426402 170000 6 reg2_val0[25]
port 1065 nsew signal output
rlabel metal2 s 427358 169200 427414 170000 6 reg2_val0[26]
port 1066 nsew signal output
rlabel metal2 s 428370 169200 428426 170000 6 reg2_val0[27]
port 1067 nsew signal output
rlabel metal2 s 429382 169200 429438 170000 6 reg2_val0[28]
port 1068 nsew signal output
rlabel metal2 s 430394 169200 430450 170000 6 reg2_val0[29]
port 1069 nsew signal output
rlabel metal2 s 403070 169200 403126 170000 6 reg2_val0[2]
port 1070 nsew signal output
rlabel metal2 s 431406 169200 431462 170000 6 reg2_val0[30]
port 1071 nsew signal output
rlabel metal2 s 432418 169200 432474 170000 6 reg2_val0[31]
port 1072 nsew signal output
rlabel metal2 s 404082 169200 404138 170000 6 reg2_val0[3]
port 1073 nsew signal output
rlabel metal2 s 405094 169200 405150 170000 6 reg2_val0[4]
port 1074 nsew signal output
rlabel metal2 s 406106 169200 406162 170000 6 reg2_val0[5]
port 1075 nsew signal output
rlabel metal2 s 407118 169200 407174 170000 6 reg2_val0[6]
port 1076 nsew signal output
rlabel metal2 s 408130 169200 408186 170000 6 reg2_val0[7]
port 1077 nsew signal output
rlabel metal2 s 409142 169200 409198 170000 6 reg2_val0[8]
port 1078 nsew signal output
rlabel metal2 s 410154 169200 410210 170000 6 reg2_val0[9]
port 1079 nsew signal output
rlabel metal3 s 439200 133016 440000 133136 6 reg2_val1[0]
port 1080 nsew signal output
rlabel metal3 s 439200 138456 440000 138576 6 reg2_val1[10]
port 1081 nsew signal output
rlabel metal3 s 439200 139000 440000 139120 6 reg2_val1[11]
port 1082 nsew signal output
rlabel metal3 s 439200 139544 440000 139664 6 reg2_val1[12]
port 1083 nsew signal output
rlabel metal3 s 439200 140088 440000 140208 6 reg2_val1[13]
port 1084 nsew signal output
rlabel metal3 s 439200 140632 440000 140752 6 reg2_val1[14]
port 1085 nsew signal output
rlabel metal3 s 439200 141176 440000 141296 6 reg2_val1[15]
port 1086 nsew signal output
rlabel metal3 s 439200 141720 440000 141840 6 reg2_val1[16]
port 1087 nsew signal output
rlabel metal3 s 439200 142264 440000 142384 6 reg2_val1[17]
port 1088 nsew signal output
rlabel metal3 s 439200 142808 440000 142928 6 reg2_val1[18]
port 1089 nsew signal output
rlabel metal3 s 439200 143352 440000 143472 6 reg2_val1[19]
port 1090 nsew signal output
rlabel metal3 s 439200 133560 440000 133680 6 reg2_val1[1]
port 1091 nsew signal output
rlabel metal3 s 439200 143896 440000 144016 6 reg2_val1[20]
port 1092 nsew signal output
rlabel metal3 s 439200 144440 440000 144560 6 reg2_val1[21]
port 1093 nsew signal output
rlabel metal3 s 439200 144984 440000 145104 6 reg2_val1[22]
port 1094 nsew signal output
rlabel metal3 s 439200 145528 440000 145648 6 reg2_val1[23]
port 1095 nsew signal output
rlabel metal3 s 439200 146072 440000 146192 6 reg2_val1[24]
port 1096 nsew signal output
rlabel metal3 s 439200 146616 440000 146736 6 reg2_val1[25]
port 1097 nsew signal output
rlabel metal3 s 439200 147160 440000 147280 6 reg2_val1[26]
port 1098 nsew signal output
rlabel metal3 s 439200 147704 440000 147824 6 reg2_val1[27]
port 1099 nsew signal output
rlabel metal3 s 439200 148248 440000 148368 6 reg2_val1[28]
port 1100 nsew signal output
rlabel metal3 s 439200 148792 440000 148912 6 reg2_val1[29]
port 1101 nsew signal output
rlabel metal3 s 439200 134104 440000 134224 6 reg2_val1[2]
port 1102 nsew signal output
rlabel metal3 s 439200 149336 440000 149456 6 reg2_val1[30]
port 1103 nsew signal output
rlabel metal3 s 439200 149880 440000 150000 6 reg2_val1[31]
port 1104 nsew signal output
rlabel metal3 s 439200 134648 440000 134768 6 reg2_val1[3]
port 1105 nsew signal output
rlabel metal3 s 439200 135192 440000 135312 6 reg2_val1[4]
port 1106 nsew signal output
rlabel metal3 s 439200 135736 440000 135856 6 reg2_val1[5]
port 1107 nsew signal output
rlabel metal3 s 439200 136280 440000 136400 6 reg2_val1[6]
port 1108 nsew signal output
rlabel metal3 s 439200 136824 440000 136944 6 reg2_val1[7]
port 1109 nsew signal output
rlabel metal3 s 439200 137368 440000 137488 6 reg2_val1[8]
port 1110 nsew signal output
rlabel metal3 s 439200 137912 440000 138032 6 reg2_val1[9]
port 1111 nsew signal output
rlabel metal3 s 0 131928 800 132048 6 reg2_val2[0]
port 1112 nsew signal output
rlabel metal3 s 0 137368 800 137488 6 reg2_val2[10]
port 1113 nsew signal output
rlabel metal3 s 0 137912 800 138032 6 reg2_val2[11]
port 1114 nsew signal output
rlabel metal3 s 0 138456 800 138576 6 reg2_val2[12]
port 1115 nsew signal output
rlabel metal3 s 0 139000 800 139120 6 reg2_val2[13]
port 1116 nsew signal output
rlabel metal3 s 0 139544 800 139664 6 reg2_val2[14]
port 1117 nsew signal output
rlabel metal3 s 0 140088 800 140208 6 reg2_val2[15]
port 1118 nsew signal output
rlabel metal3 s 0 140632 800 140752 6 reg2_val2[16]
port 1119 nsew signal output
rlabel metal3 s 0 141176 800 141296 6 reg2_val2[17]
port 1120 nsew signal output
rlabel metal3 s 0 141720 800 141840 6 reg2_val2[18]
port 1121 nsew signal output
rlabel metal3 s 0 142264 800 142384 6 reg2_val2[19]
port 1122 nsew signal output
rlabel metal3 s 0 132472 800 132592 6 reg2_val2[1]
port 1123 nsew signal output
rlabel metal3 s 0 142808 800 142928 6 reg2_val2[20]
port 1124 nsew signal output
rlabel metal3 s 0 143352 800 143472 6 reg2_val2[21]
port 1125 nsew signal output
rlabel metal3 s 0 143896 800 144016 6 reg2_val2[22]
port 1126 nsew signal output
rlabel metal3 s 0 144440 800 144560 6 reg2_val2[23]
port 1127 nsew signal output
rlabel metal3 s 0 144984 800 145104 6 reg2_val2[24]
port 1128 nsew signal output
rlabel metal3 s 0 145528 800 145648 6 reg2_val2[25]
port 1129 nsew signal output
rlabel metal3 s 0 146072 800 146192 6 reg2_val2[26]
port 1130 nsew signal output
rlabel metal3 s 0 146616 800 146736 6 reg2_val2[27]
port 1131 nsew signal output
rlabel metal3 s 0 147160 800 147280 6 reg2_val2[28]
port 1132 nsew signal output
rlabel metal3 s 0 147704 800 147824 6 reg2_val2[29]
port 1133 nsew signal output
rlabel metal3 s 0 133016 800 133136 6 reg2_val2[2]
port 1134 nsew signal output
rlabel metal3 s 0 148248 800 148368 6 reg2_val2[30]
port 1135 nsew signal output
rlabel metal3 s 0 148792 800 148912 6 reg2_val2[31]
port 1136 nsew signal output
rlabel metal3 s 0 133560 800 133680 6 reg2_val2[3]
port 1137 nsew signal output
rlabel metal3 s 0 134104 800 134224 6 reg2_val2[4]
port 1138 nsew signal output
rlabel metal3 s 0 134648 800 134768 6 reg2_val2[5]
port 1139 nsew signal output
rlabel metal3 s 0 135192 800 135312 6 reg2_val2[6]
port 1140 nsew signal output
rlabel metal3 s 0 135736 800 135856 6 reg2_val2[7]
port 1141 nsew signal output
rlabel metal3 s 0 136280 800 136400 6 reg2_val2[8]
port 1142 nsew signal output
rlabel metal3 s 0 136824 800 136944 6 reg2_val2[9]
port 1143 nsew signal output
rlabel metal2 s 163226 169200 163282 170000 6 rst_eu
port 1144 nsew signal output
rlabel metal2 s 422666 0 422722 800 6 rst_n
port 1145 nsew signal input
rlabel metal2 s 286690 169200 286746 170000 6 sign_extend0
port 1146 nsew signal input
rlabel metal3 s 439200 71544 440000 71664 6 sign_extend1
port 1147 nsew signal input
rlabel metal3 s 0 70456 800 70576 6 sign_extend2
port 1148 nsew signal input
rlabel metal2 s 295798 169200 295854 170000 6 take_branch0
port 1149 nsew signal input
rlabel metal3 s 439200 76440 440000 76560 6 take_branch1
port 1150 nsew signal input
rlabel metal3 s 0 75352 800 75472 6 take_branch2
port 1151 nsew signal input
rlabel metal4 s 4208 2128 4528 167600 6 vccd1
port 1152 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 167600 6 vccd1
port 1152 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 167600 6 vccd1
port 1152 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 167600 6 vccd1
port 1152 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 167600 6 vccd1
port 1152 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 167600 6 vccd1
port 1152 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 167600 6 vccd1
port 1152 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 167600 6 vccd1
port 1152 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 167600 6 vccd1
port 1152 nsew power bidirectional
rlabel metal4 s 280688 2128 281008 167600 6 vccd1
port 1152 nsew power bidirectional
rlabel metal4 s 311408 2128 311728 167600 6 vccd1
port 1152 nsew power bidirectional
rlabel metal4 s 342128 2128 342448 167600 6 vccd1
port 1152 nsew power bidirectional
rlabel metal4 s 372848 2128 373168 167600 6 vccd1
port 1152 nsew power bidirectional
rlabel metal4 s 403568 2128 403888 167600 6 vccd1
port 1152 nsew power bidirectional
rlabel metal4 s 434288 2128 434608 167600 6 vccd1
port 1152 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 167600 6 vssd1
port 1153 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 167600 6 vssd1
port 1153 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 167600 6 vssd1
port 1153 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 167600 6 vssd1
port 1153 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 167600 6 vssd1
port 1153 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 167600 6 vssd1
port 1153 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 167600 6 vssd1
port 1153 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 167600 6 vssd1
port 1153 nsew ground bidirectional
rlabel metal4 s 265328 2128 265648 167600 6 vssd1
port 1153 nsew ground bidirectional
rlabel metal4 s 296048 2128 296368 167600 6 vssd1
port 1153 nsew ground bidirectional
rlabel metal4 s 326768 2128 327088 167600 6 vssd1
port 1153 nsew ground bidirectional
rlabel metal4 s 357488 2128 357808 167600 6 vssd1
port 1153 nsew ground bidirectional
rlabel metal4 s 388208 2128 388528 167600 6 vssd1
port 1153 nsew ground bidirectional
rlabel metal4 s 418928 2128 419248 167600 6 vssd1
port 1153 nsew ground bidirectional
rlabel metal2 s 420918 0 420974 800 6 wb_clk_i
port 1154 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 440000 170000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 162567086
string GDS_FILE /home/tholin/Desktop/ci2406-rej-pommedeterrible-tholin/openlane/VLIW/runs/24_06_04_23_19/results/signoff/vliw.magic.gds
string GDS_START 1467820
<< end >>

