// This is the unpowered netlist.
module ci2406_z80 (rst_n,
    wb_clk_i,
    custom_settings,
    io_in,
    io_oeb,
    io_out);
 input rst_n;
 input wb_clk_i;
 input [4:0] custom_settings;
 input [35:0] io_in;
 output [35:0] io_oeb;
 output [35:0] io_out;

 wire net186;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net187;
 wire net205;
 wire net206;
 wire net188;
 wire net215;
 wire net216;
 wire net207;
 wire net208;
 wire net209;
 wire net217;
 wire net189;
 wire net214;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net211;
 wire net212;
 wire net213;
 wire net210;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire clknet_0_wb_clk_i;
 wire clknet_2_0__leaf_wb_clk_i;
 wire clknet_2_1__leaf_wb_clk_i;
 wire clknet_2_2__leaf_wb_clk_i;
 wire clknet_2_3__leaf_wb_clk_i;
 wire clknet_leaf_0_wb_clk_i;
 wire clknet_leaf_10_wb_clk_i;
 wire clknet_leaf_11_wb_clk_i;
 wire clknet_leaf_12_wb_clk_i;
 wire clknet_leaf_13_wb_clk_i;
 wire clknet_leaf_14_wb_clk_i;
 wire clknet_leaf_15_wb_clk_i;
 wire clknet_leaf_16_wb_clk_i;
 wire clknet_leaf_18_wb_clk_i;
 wire clknet_leaf_19_wb_clk_i;
 wire clknet_leaf_1_wb_clk_i;
 wire clknet_leaf_20_wb_clk_i;
 wire clknet_leaf_21_wb_clk_i;
 wire clknet_leaf_22_wb_clk_i;
 wire clknet_leaf_23_wb_clk_i;
 wire clknet_leaf_24_wb_clk_i;
 wire clknet_leaf_25_wb_clk_i;
 wire clknet_leaf_26_wb_clk_i;
 wire clknet_leaf_27_wb_clk_i;
 wire clknet_leaf_28_wb_clk_i;
 wire clknet_leaf_29_wb_clk_i;
 wire clknet_leaf_2_wb_clk_i;
 wire clknet_leaf_30_wb_clk_i;
 wire clknet_leaf_31_wb_clk_i;
 wire clknet_leaf_32_wb_clk_i;
 wire clknet_leaf_33_wb_clk_i;
 wire clknet_leaf_34_wb_clk_i;
 wire clknet_leaf_35_wb_clk_i;
 wire clknet_leaf_36_wb_clk_i;
 wire clknet_leaf_37_wb_clk_i;
 wire clknet_leaf_38_wb_clk_i;
 wire clknet_leaf_39_wb_clk_i;
 wire clknet_leaf_3_wb_clk_i;
 wire clknet_leaf_40_wb_clk_i;
 wire clknet_leaf_41_wb_clk_i;
 wire clknet_leaf_42_wb_clk_i;
 wire clknet_leaf_43_wb_clk_i;
 wire clknet_leaf_44_wb_clk_i;
 wire clknet_leaf_45_wb_clk_i;
 wire clknet_leaf_46_wb_clk_i;
 wire clknet_leaf_47_wb_clk_i;
 wire clknet_leaf_48_wb_clk_i;
 wire clknet_leaf_49_wb_clk_i;
 wire clknet_leaf_4_wb_clk_i;
 wire clknet_leaf_50_wb_clk_i;
 wire clknet_leaf_5_wb_clk_i;
 wire clknet_leaf_6_wb_clk_i;
 wire clknet_leaf_7_wb_clk_i;
 wire clknet_leaf_8_wb_clk_i;
 wire clknet_leaf_9_wb_clk_i;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net79;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net8;
 wire net80;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net81;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net82;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net83;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net84;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net85;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net86;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net87;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net88;
 wire net880;
 wire net881;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire \z80.early_iorq_n ;
 wire \z80.early_mreq_n ;
 wire \z80.early_rd_n ;
 wire \z80.normal_iorq_n ;
 wire \z80.normal_mreq_n ;
 wire \z80.normal_rd_n ;
 wire \z80.tv80s.di_reg[0] ;
 wire \z80.tv80s.di_reg[1] ;
 wire \z80.tv80s.di_reg[2] ;
 wire \z80.tv80s.di_reg[3] ;
 wire \z80.tv80s.di_reg[4] ;
 wire \z80.tv80s.di_reg[5] ;
 wire \z80.tv80s.di_reg[6] ;
 wire \z80.tv80s.di_reg[7] ;
 wire \z80.tv80s.i_tv80_core.ACC[0] ;
 wire \z80.tv80s.i_tv80_core.ACC[1] ;
 wire \z80.tv80s.i_tv80_core.ACC[2] ;
 wire \z80.tv80s.i_tv80_core.ACC[3] ;
 wire \z80.tv80s.i_tv80_core.ACC[4] ;
 wire \z80.tv80s.i_tv80_core.ACC[5] ;
 wire \z80.tv80s.i_tv80_core.ACC[6] ;
 wire \z80.tv80s.i_tv80_core.ACC[7] ;
 wire \z80.tv80s.i_tv80_core.ALU_Op_r[0] ;
 wire \z80.tv80s.i_tv80_core.ALU_Op_r[1] ;
 wire \z80.tv80s.i_tv80_core.ALU_Op_r[2] ;
 wire \z80.tv80s.i_tv80_core.ALU_Op_r[3] ;
 wire \z80.tv80s.i_tv80_core.Alternate ;
 wire \z80.tv80s.i_tv80_core.Ap[0] ;
 wire \z80.tv80s.i_tv80_core.Ap[1] ;
 wire \z80.tv80s.i_tv80_core.Ap[2] ;
 wire \z80.tv80s.i_tv80_core.Ap[3] ;
 wire \z80.tv80s.i_tv80_core.Ap[4] ;
 wire \z80.tv80s.i_tv80_core.Ap[5] ;
 wire \z80.tv80s.i_tv80_core.Ap[6] ;
 wire \z80.tv80s.i_tv80_core.Ap[7] ;
 wire \z80.tv80s.i_tv80_core.Arith16_r ;
 wire \z80.tv80s.i_tv80_core.Auto_Wait_t1 ;
 wire \z80.tv80s.i_tv80_core.Auto_Wait_t2 ;
 wire \z80.tv80s.i_tv80_core.BTR_r ;
 wire \z80.tv80s.i_tv80_core.BusA[0] ;
 wire \z80.tv80s.i_tv80_core.BusA[1] ;
 wire \z80.tv80s.i_tv80_core.BusA[2] ;
 wire \z80.tv80s.i_tv80_core.BusA[3] ;
 wire \z80.tv80s.i_tv80_core.BusA[4] ;
 wire \z80.tv80s.i_tv80_core.BusA[5] ;
 wire \z80.tv80s.i_tv80_core.BusA[6] ;
 wire \z80.tv80s.i_tv80_core.BusA[7] ;
 wire \z80.tv80s.i_tv80_core.BusAck ;
 wire \z80.tv80s.i_tv80_core.BusB[0] ;
 wire \z80.tv80s.i_tv80_core.BusB[1] ;
 wire \z80.tv80s.i_tv80_core.BusB[2] ;
 wire \z80.tv80s.i_tv80_core.BusB[3] ;
 wire \z80.tv80s.i_tv80_core.BusB[4] ;
 wire \z80.tv80s.i_tv80_core.BusB[5] ;
 wire \z80.tv80s.i_tv80_core.BusB[6] ;
 wire \z80.tv80s.i_tv80_core.BusB[7] ;
 wire \z80.tv80s.i_tv80_core.BusReq_s ;
 wire \z80.tv80s.i_tv80_core.F[0] ;
 wire \z80.tv80s.i_tv80_core.F[1] ;
 wire \z80.tv80s.i_tv80_core.F[2] ;
 wire \z80.tv80s.i_tv80_core.F[3] ;
 wire \z80.tv80s.i_tv80_core.F[4] ;
 wire \z80.tv80s.i_tv80_core.F[5] ;
 wire \z80.tv80s.i_tv80_core.F[6] ;
 wire \z80.tv80s.i_tv80_core.F[7] ;
 wire \z80.tv80s.i_tv80_core.Fp[0] ;
 wire \z80.tv80s.i_tv80_core.Fp[1] ;
 wire \z80.tv80s.i_tv80_core.Fp[2] ;
 wire \z80.tv80s.i_tv80_core.Fp[3] ;
 wire \z80.tv80s.i_tv80_core.Fp[4] ;
 wire \z80.tv80s.i_tv80_core.Fp[5] ;
 wire \z80.tv80s.i_tv80_core.Fp[6] ;
 wire \z80.tv80s.i_tv80_core.Fp[7] ;
 wire \z80.tv80s.i_tv80_core.Halt_FF ;
 wire \z80.tv80s.i_tv80_core.INT_s ;
 wire \z80.tv80s.i_tv80_core.IR[0] ;
 wire \z80.tv80s.i_tv80_core.IR[1] ;
 wire \z80.tv80s.i_tv80_core.IR[2] ;
 wire \z80.tv80s.i_tv80_core.IR[3] ;
 wire \z80.tv80s.i_tv80_core.IR[4] ;
 wire \z80.tv80s.i_tv80_core.IR[5] ;
 wire \z80.tv80s.i_tv80_core.IR[6] ;
 wire \z80.tv80s.i_tv80_core.IR[7] ;
 wire \z80.tv80s.i_tv80_core.ISet[0] ;
 wire \z80.tv80s.i_tv80_core.ISet[1] ;
 wire \z80.tv80s.i_tv80_core.ISet[2] ;
 wire \z80.tv80s.i_tv80_core.ISet[3] ;
 wire \z80.tv80s.i_tv80_core.IStatus[1] ;
 wire \z80.tv80s.i_tv80_core.IStatus[2] ;
 wire \z80.tv80s.i_tv80_core.I[0] ;
 wire \z80.tv80s.i_tv80_core.I[1] ;
 wire \z80.tv80s.i_tv80_core.I[2] ;
 wire \z80.tv80s.i_tv80_core.I[3] ;
 wire \z80.tv80s.i_tv80_core.I[4] ;
 wire \z80.tv80s.i_tv80_core.I[5] ;
 wire \z80.tv80s.i_tv80_core.I[6] ;
 wire \z80.tv80s.i_tv80_core.I[7] ;
 wire \z80.tv80s.i_tv80_core.IncDecZ ;
 wire \z80.tv80s.i_tv80_core.IntCycle ;
 wire \z80.tv80s.i_tv80_core.IntE ;
 wire \z80.tv80s.i_tv80_core.IntE_FF2 ;
 wire \z80.tv80s.i_tv80_core.NMICycle ;
 wire \z80.tv80s.i_tv80_core.NMI_s ;
 wire \z80.tv80s.i_tv80_core.No_BTR ;
 wire \z80.tv80s.i_tv80_core.Oldnmi_n ;
 wire \z80.tv80s.i_tv80_core.PC[0] ;
 wire \z80.tv80s.i_tv80_core.PC[10] ;
 wire \z80.tv80s.i_tv80_core.PC[11] ;
 wire \z80.tv80s.i_tv80_core.PC[12] ;
 wire \z80.tv80s.i_tv80_core.PC[13] ;
 wire \z80.tv80s.i_tv80_core.PC[14] ;
 wire \z80.tv80s.i_tv80_core.PC[15] ;
 wire \z80.tv80s.i_tv80_core.PC[1] ;
 wire \z80.tv80s.i_tv80_core.PC[2] ;
 wire \z80.tv80s.i_tv80_core.PC[3] ;
 wire \z80.tv80s.i_tv80_core.PC[4] ;
 wire \z80.tv80s.i_tv80_core.PC[5] ;
 wire \z80.tv80s.i_tv80_core.PC[6] ;
 wire \z80.tv80s.i_tv80_core.PC[7] ;
 wire \z80.tv80s.i_tv80_core.PC[8] ;
 wire \z80.tv80s.i_tv80_core.PC[9] ;
 wire \z80.tv80s.i_tv80_core.Pre_XY_F_M[1] ;
 wire \z80.tv80s.i_tv80_core.Pre_XY_F_M[2] ;
 wire \z80.tv80s.i_tv80_core.Pre_XY_F_M[3] ;
 wire \z80.tv80s.i_tv80_core.Pre_XY_F_M[4] ;
 wire \z80.tv80s.i_tv80_core.Pre_XY_F_M[5] ;
 wire \z80.tv80s.i_tv80_core.Pre_XY_F_M[6] ;
 wire \z80.tv80s.i_tv80_core.Pre_XY_F_M[7] ;
 wire \z80.tv80s.i_tv80_core.PreserveC_r ;
 wire \z80.tv80s.i_tv80_core.R[0] ;
 wire \z80.tv80s.i_tv80_core.R[1] ;
 wire \z80.tv80s.i_tv80_core.R[2] ;
 wire \z80.tv80s.i_tv80_core.R[3] ;
 wire \z80.tv80s.i_tv80_core.R[4] ;
 wire \z80.tv80s.i_tv80_core.R[5] ;
 wire \z80.tv80s.i_tv80_core.R[6] ;
 wire \z80.tv80s.i_tv80_core.R[7] ;
 wire \z80.tv80s.i_tv80_core.Read_To_Reg_r[0] ;
 wire \z80.tv80s.i_tv80_core.Read_To_Reg_r[1] ;
 wire \z80.tv80s.i_tv80_core.Read_To_Reg_r[2] ;
 wire \z80.tv80s.i_tv80_core.Read_To_Reg_r[3] ;
 wire \z80.tv80s.i_tv80_core.Read_To_Reg_r[4] ;
 wire \z80.tv80s.i_tv80_core.RegAddrA_r[0] ;
 wire \z80.tv80s.i_tv80_core.RegAddrA_r[1] ;
 wire \z80.tv80s.i_tv80_core.RegAddrA_r[2] ;
 wire \z80.tv80s.i_tv80_core.RegAddrB_r[0] ;
 wire \z80.tv80s.i_tv80_core.RegAddrB_r[1] ;
 wire \z80.tv80s.i_tv80_core.RegAddrB_r[2] ;
 wire \z80.tv80s.i_tv80_core.RegAddrC[0] ;
 wire \z80.tv80s.i_tv80_core.RegAddrC[1] ;
 wire \z80.tv80s.i_tv80_core.RegAddrC[2] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[0] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[10] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[11] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[12] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[13] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[14] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[15] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[1] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[2] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[3] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[4] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[5] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[6] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[7] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[8] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[9] ;
 wire \z80.tv80s.i_tv80_core.SP[0] ;
 wire \z80.tv80s.i_tv80_core.SP[10] ;
 wire \z80.tv80s.i_tv80_core.SP[11] ;
 wire \z80.tv80s.i_tv80_core.SP[12] ;
 wire \z80.tv80s.i_tv80_core.SP[13] ;
 wire \z80.tv80s.i_tv80_core.SP[14] ;
 wire \z80.tv80s.i_tv80_core.SP[15] ;
 wire \z80.tv80s.i_tv80_core.SP[1] ;
 wire \z80.tv80s.i_tv80_core.SP[2] ;
 wire \z80.tv80s.i_tv80_core.SP[3] ;
 wire \z80.tv80s.i_tv80_core.SP[4] ;
 wire \z80.tv80s.i_tv80_core.SP[5] ;
 wire \z80.tv80s.i_tv80_core.SP[6] ;
 wire \z80.tv80s.i_tv80_core.SP[7] ;
 wire \z80.tv80s.i_tv80_core.SP[8] ;
 wire \z80.tv80s.i_tv80_core.SP[9] ;
 wire \z80.tv80s.i_tv80_core.Save_ALU_r ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[0] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[10] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[11] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[12] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[13] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[14] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[15] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[1] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[2] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[3] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[4] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[5] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[6] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[7] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[8] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[9] ;
 wire \z80.tv80s.i_tv80_core.XY_Ind ;
 wire \z80.tv80s.i_tv80_core.XY_State[0] ;
 wire \z80.tv80s.i_tv80_core.XY_State[1] ;
 wire \z80.tv80s.i_tv80_core.Z16_r ;
 wire \z80.tv80s.i_tv80_core.i_mcode.MCycle[0] ;
 wire \z80.tv80s.i_tv80_core.i_mcode.MCycle[1] ;
 wire \z80.tv80s.i_tv80_core.i_mcode.MCycle[2] ;
 wire \z80.tv80s.i_tv80_core.i_mcode.MCycle[3] ;
 wire \z80.tv80s.i_tv80_core.i_mcode.MCycle[4] ;
 wire \z80.tv80s.i_tv80_core.i_mcode.MCycle[5] ;
 wire \z80.tv80s.i_tv80_core.i_mcode.MCycle[6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[0][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[0][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[0][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[0][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[0][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[0][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[0][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[0][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[1][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[1][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[1][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[1][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[1][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[1][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[1][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[1][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[2][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[2][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[2][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[2][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[2][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[2][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[2][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[2][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[3][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[3][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[3][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[3][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[3][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[3][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[3][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[3][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[4][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[4][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[4][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[4][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[4][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[4][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[4][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[4][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[5][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[5][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[5][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[5][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[5][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[5][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[5][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[5][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[6][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[6][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[6][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[6][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[6][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[6][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[6][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[6][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[7][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[7][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[7][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[7][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[7][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[7][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[7][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[7][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[0][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[0][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[0][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[0][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[0][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[0][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[0][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[0][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[1][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[1][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[1][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[1][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[1][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[1][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[1][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[1][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[2][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[2][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[2][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[2][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[2][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[2][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[2][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[2][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[3][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[3][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[3][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[3][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[3][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[3][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[3][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[3][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[4][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[4][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[4][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[4][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[4][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[4][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[4][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[4][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[5][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[5][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[5][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[5][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[5][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[5][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[5][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[5][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[6][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[6][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[6][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[6][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[6][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[6][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[6][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[6][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[7][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[7][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[7][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[7][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[7][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[7][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[7][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[7][7] ;
 wire \z80.tv80s.i_tv80_core.mcycles[1] ;
 wire \z80.tv80s.i_tv80_core.mcycles[2] ;
 wire \z80.tv80s.i_tv80_core.mcycles[4] ;
 wire \z80.tv80s.i_tv80_core.mcycles[5] ;
 wire \z80.tv80s.i_tv80_core.ts[0] ;
 wire \z80.tv80s.i_tv80_core.ts[1] ;
 wire \z80.tv80s.i_tv80_core.ts[2] ;
 wire \z80.tv80s.i_tv80_core.ts[3] ;
 wire \z80.tv80s.i_tv80_core.ts[4] ;
 wire \z80.tv80s.i_tv80_core.ts[5] ;
 wire \z80.tv80s.i_tv80_core.ts[6] ;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_0475_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_0498_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_1245_));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_2526_));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_2872_));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(\z80.tv80s.i_tv80_core.BusAck ));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(\z80.tv80s.i_tv80_core.F[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(_1822_));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(_2992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3054__A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__3055__A (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__3059__A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__3062__A (.DIODE(\z80.tv80s.i_tv80_core.ISet[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3063__A (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__3066__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__3070__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__3071__A (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__3072__A (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__3074__A (.DIODE(\z80.tv80s.i_tv80_core.Halt_FF ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3078__A (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__3079__A (.DIODE(\z80.tv80s.i_tv80_core.BusA[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3080__A (.DIODE(\z80.tv80s.i_tv80_core.BusA[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3082__A (.DIODE(\z80.tv80s.i_tv80_core.BusB[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3085__A (.DIODE(\z80.tv80s.di_reg[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3086__A (.DIODE(\z80.tv80s.di_reg[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3090__A (.DIODE(\z80.tv80s.i_tv80_core.ACC[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3092__A (.DIODE(\z80.tv80s.i_tv80_core.ACC[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3093__A (.DIODE(\z80.tv80s.i_tv80_core.ACC[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3104__C_N (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__3105__A (.DIODE(_2846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3107__A_N (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__3109__B (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__3116__A (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__3116__B (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__3117__B (.DIODE(_2899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3118__A (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__3118__B (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__3119__B (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__3120__A_N (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__3120__B (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__3120__C (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__3121__A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__3122__A1 (.DIODE(_2893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3122__A2 (.DIODE(_2904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3122__B1 (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3123__B (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__3124__B (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__3125__B (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__3125__D (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__3126__B (.DIODE(_2899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3127__B (.DIODE(_2899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3128__A (.DIODE(_2846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3128__B (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__3131__A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__3132__A (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__3133__A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__3136__C_N (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__3136__D_N (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__3138__A (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__3138__B (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__3139__A (.DIODE(_2846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3139__B (.DIODE(_2847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3141__A (.DIODE(_2904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3142__A (.DIODE(_2904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3144__A (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__3144__B (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__3144__C (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__3145__B (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__3147__A (.DIODE(_2929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3148__C (.DIODE(_2929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3150__A (.DIODE(_2847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3150__C (.DIODE(_2927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3151__A (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__3151__B (.DIODE(_2847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3152__A_N (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__3152__B (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__3156__B (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__3156__D (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__3157__A (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__3167__A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__3168__A (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__3168__B (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__3169__B (.DIODE(_2899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3170__A (.DIODE(_2950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3170__B (.DIODE(_2952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3171__A1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__3172__A (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__3173__A0 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__3178__A (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__3179__A (.DIODE(_2960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3180__A (.DIODE(_2960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3181__C (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__3181__D_N (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__3184__A (.DIODE(_2847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3190__C1 (.DIODE(_2899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3194__B (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__3194__D_N (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__3195__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__3195__A2 (.DIODE(_2960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3201__A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__3202__A1 (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3202__A3 (.DIODE(_2982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3202__C1 (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3204__C (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__3205__B (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__3207__B1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__3208__A (.DIODE(_2960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3209__A (.DIODE(_2960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3210__A (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__3212__A (.DIODE(_2846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3212__B (.DIODE(_2847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3213__A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__3213__B (.DIODE(_2927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3213__D (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__3215__A (.DIODE(_2847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3215__B (.DIODE(_2927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3216__C (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__3217__A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__3217__B (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__3218__A_N (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__3218__B (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__3222__A1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__3227__A1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__3231__B (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__3232__A (.DIODE(_2899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3232__D (.DIODE(_2982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3234__A1 (.DIODE(_2846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3237__A (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__3237__D_N (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__3239__B (.DIODE(_3021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3243__B (.DIODE(_2960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3244__B (.DIODE(_2960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3245__A1 (.DIODE(_2847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3245__B2 (.DIODE(_2934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3246__A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__3246__B (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__3250__A (.DIODE(_2847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3256__A (.DIODE(_2960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3259__A (.DIODE(_2899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3260__A1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__3261__A (.DIODE(_3040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3270__C1 (.DIODE(_3052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3276__B (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__3277__B (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__3281__A (.DIODE(_2927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3281__B (.DIODE(_2934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3284__A (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__3284__B (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__3285__A (.DIODE(_2994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3286__B (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__3287__A (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__3287__B (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__3288__A2 (.DIODE(_0398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3289__B (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__3291__B1 (.DIODE(_0401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3291__B2 (.DIODE(_3040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3291__C1 (.DIODE(_2994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3292__B1 (.DIODE(_0401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3294__A (.DIODE(_2847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3296__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__3297__B (.DIODE(_2995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3298__A1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__3298__B1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__3299__B1 (.DIODE(_2982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3300__C (.DIODE(_3021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3304__B (.DIODE(_2960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3318__B (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__3319__B (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__3320__A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__3320__B (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3321__A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__3321__B (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__3321__C (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__3324__A (.DIODE(_0400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3331__A (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__3333__A (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__3337__B (.DIODE(_3052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3338__A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__3339__A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__3340__A2 (.DIODE(_0450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3342__A1 (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3343__A1 (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3345__A1 (.DIODE(_2960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3346__A1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__3351__A (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__3351__B (.DIODE(_2849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3352__B (.DIODE(_2994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3355__A_N (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__3356__B (.DIODE(\z80.tv80s.i_tv80_core.F[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3357__B (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__3357__C (.DIODE(_2847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3358__A_N (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__3358__B (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__3361__C (.DIODE(\z80.tv80s.i_tv80_core.F[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3362__B2 (.DIODE(\z80.tv80s.i_tv80_core.F[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3363__A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__3365__S (.DIODE(\z80.tv80s.i_tv80_core.F[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3366__A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__3366__B (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__3367__B1_N (.DIODE(\z80.tv80s.i_tv80_core.F[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3368__A1 (.DIODE(_0477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3369__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3371__A1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__3371__A3 (.DIODE(_0481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3371__B1 (.DIODE(_0400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3373__A (.DIODE(\z80.tv80s.i_tv80_core.IntCycle ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3375__A1 (.DIODE(_0401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3377__A (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__3378__D (.DIODE(_0398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3381__A1 (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3381__B1 (.DIODE(_0450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3385__A (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__3388__A1 (.DIODE(_2893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3388__A2 (.DIODE(_2904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3391__A1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__3391__B1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__3392__A (.DIODE(_2904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3392__D (.DIODE(_2929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3395__A2 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__3396__A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__3397__A1 (.DIODE(_2934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3400__B1 (.DIODE(_2849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3401__B (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__3402__B (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__3403__A (.DIODE(_0481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3403__B (.DIODE(_0513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3404__A (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__3406__A1 (.DIODE(_0398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3407__A1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__3408__C1 (.DIODE(_3021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3412__A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__3415__B2 (.DIODE(_0400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3418__A1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__3421__A (.DIODE(_2998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3422__A2 (.DIODE(_0400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3424__A (.DIODE(_2998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3427__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__3427__B (.DIODE(_0537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3428__A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__3429__A (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__3432__B1 (.DIODE(_2849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3434__A (.DIODE(_3021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3435__A1 (.DIODE(_3021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3436__B1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__3442__A (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__3444__A (.DIODE(_2849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3444__B (.DIODE(_0554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3445__A2 (.DIODE(_3052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3445__B1 (.DIODE(_0450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3446__B (.DIODE(_0554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3447__B (.DIODE(_0513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3448__A1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__3448__B1 (.DIODE(_2998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3451__B1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__3452__B1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__3453__B2 (.DIODE(_0400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3458__A1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__3459__C1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__3460__C (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__3466__A (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__3467__B (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__3468__A (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__3471__A (.DIODE(_0502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3472__A (.DIODE(_2893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3473__B (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA__3475__A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__3475__B (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA__3477__C (.DIODE(_0397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3481__A (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__3483__B2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__3485__A1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__3489__B (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__3490__A1 (.DIODE(_2893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3490__C1 (.DIODE(_0502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3495__A1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__3496__A1 (.DIODE(_2854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3496__B1 (.DIODE(_2849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3497__B (.DIODE(_2904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3498__A1 (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA__3498__A3 (.DIODE(_2904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3498__B1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__3499__A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__3499__B (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__3500__B (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__3501__B (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__3502__A1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__3502__A2 (.DIODE(_0604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3502__B1 (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA__3503__B (.DIODE(_0605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3504__A (.DIODE(_2849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3504__B (.DIODE(_0604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3505__B (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__3505__C (.DIODE(_0603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3506__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__3506__B (.DIODE(_0607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3509__A1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__3512__A (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__3513__A2_N (.DIODE(_2982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3515__A1 (.DIODE(_0405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3516__B1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__3517__B1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__3518__A2 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__3519__B1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__3520__A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__3521__A1 (.DIODE(_0481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3522__C (.DIODE(\z80.tv80s.i_tv80_core.IntCycle ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3523__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__3523__B (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__3525__A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__3526__A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__3526__B2 (.DIODE(_0626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3528__B2 (.DIODE(_2934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3529__A1 (.DIODE(_0405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3530__A (.DIODE(_2893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3531__A1 (.DIODE(_2849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3532__A_N (.DIODE(_0481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3532__C (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__3535__A1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__3536__A2 (.DIODE(_0481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3537__B (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__3537__C (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__3538__A2 (.DIODE(_2994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3540__B1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__3542__A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__3543__B2 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__3544__A2 (.DIODE(_0626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3549__A (.DIODE(_2846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3549__B (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__3549__C (.DIODE(_2982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3550__A (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__3550__C (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__3551__B1 (.DIODE(_0626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3552__A1 (.DIODE(_0626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3553__A1 (.DIODE(_0626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3555__A1 (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA__3555__B2 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__3559__B1 (.DIODE(_0397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3561__A (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__3561__B (.DIODE(_0513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3562__B (.DIODE(_0513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3563__A1_N (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3563__B2 (.DIODE(_0653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3564__B1 (.DIODE(_0554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3565__A1 (.DIODE(_2899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3568__A (.DIODE(_0398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3569__A (.DIODE(_0398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3570__A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__3572__A1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__3573__C1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__3574__A (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3574__C (.DIODE(_0653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3575__A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__3576__B (.DIODE(_0554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3577__C1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__3578__A2 (.DIODE(_0653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3580__B (.DIODE(_0513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3581__B (.DIODE(_3040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3582__C1 (.DIODE(_0513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3583__A1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__3583__A2 (.DIODE(_3040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3584__A1 (.DIODE(_3040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3585__C1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__3587__A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__3588__A (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__3589__B (.DIODE(_0397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3590__B (.DIODE(_0398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3591__A3 (.DIODE(_0450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3592__A1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__3592__A3 (.DIODE(_0554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3593__A2 (.DIODE(_2893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3595__A (.DIODE(_0397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3596__A1_N (.DIODE(_3021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3596__B1 (.DIODE(_0513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3597__A_N (.DIODE(_0684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3597__B (.DIODE(_0685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3598__A1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__3598__B1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__3600__A (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA__3602__A (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__3605__A2 (.DIODE(_0653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3607__A2 (.DIODE(_2927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3612__A1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__3612__A3 (.DIODE(_2927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3616__A1 (.DIODE(_2899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3619__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__3619__C (.DIODE(_0513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3622__B1 (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA__3624__B (.DIODE(_2854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3626__A2 (.DIODE(_2854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3627__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__3627__D (.DIODE(_0400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3629__A (.DIODE(_2849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3630__A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__3632__A (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__3632__B (.DIODE(\z80.tv80s.i_tv80_core.ISet[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3632__D (.DIODE(_3021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3633__B (.DIODE(_0717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3635__A (.DIODE(_0502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3636__A (.DIODE(_0502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3637__A1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__3637__A2 (.DIODE(_0607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3639__A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__3639__B (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__3640__B (.DIODE(\z80.tv80s.i_tv80_core.INT_s ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3642__B (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__3651__A1 (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA__3651__A2 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__3652__C (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__3652__D (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__3653__A1 (.DIODE(_0577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3654__A1 (.DIODE(_2849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3655__A (.DIODE(_0577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3656__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__3661__A1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__3663__B (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__3664__A1 (.DIODE(_2854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3664__A2 (.DIODE(_0604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3664__B1 (.DIODE(_2849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3666__B (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__3667__A2 (.DIODE(_2994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3667__A3 (.DIODE(_0397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3667__B1 (.DIODE(_0653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3668__A (.DIODE(_0401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3670__A (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__3672__A1 (.DIODE(_0400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3673__B (.DIODE(_0450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3674__A (.DIODE(_0400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3675__A2 (.DIODE(_0450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3675__B2 (.DIODE(_0400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3676__B1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__3676__C1 (.DIODE(_0397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3677__A1 (.DIODE(_0400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3680__A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__3682__A1 (.DIODE(_2994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3682__B1 (.DIODE(_0397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3683__A2 (.DIODE(_0653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3683__B1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__3685__A (.DIODE(_3052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3690__B1 (.DIODE(_0398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3690__B2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__3692__B1 (.DIODE(_0400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3694__A1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__3695__A2 (.DIODE(_0603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3696__B (.DIODE(_2950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3697__B (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__3697__C (.DIODE(_2950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3698__A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__3699__C (.DIODE(_2950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3701__A (.DIODE(_0772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3701__B (.DIODE(_0774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3702__B (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__3703__C (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__3705__B (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3709__C_N (.DIODE(_0781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3710__B1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__3711__A1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__3711__C1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__3715__B1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__3716__B1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__3721__B1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__3722__C1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__3725__A2 (.DIODE(_0774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3725__B1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__3726__A2 (.DIODE(_0774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3726__B1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__3727__C1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__3728__C1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__3731__B (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3732__A (.DIODE(_0794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3732__B (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__3732__C (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__3736__A (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__3736__C (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__3741__A (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__3741__B (.DIODE(\z80.tv80s.i_tv80_core.BusB[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3742__A (.DIODE(\z80.tv80s.i_tv80_core.BusA[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3743__A (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__3744__A (.DIODE(\z80.tv80s.i_tv80_core.BusA[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3745__B (.DIODE(\z80.tv80s.i_tv80_core.F[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3747__B (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__3748__A0 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__3756__A2 (.DIODE(\z80.tv80s.i_tv80_core.BusA[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3756__A3 (.DIODE(\z80.tv80s.i_tv80_core.BusB[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3757__B (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__3760__B (.DIODE(_2899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3763__A3 (.DIODE(_2899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3763__C1 (.DIODE(\z80.tv80s.i_tv80_core.BusB[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3765__A2 (.DIODE(\z80.tv80s.i_tv80_core.F[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3765__B1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__3766__A1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__3767__A1 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__3771__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusB[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3771__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusB[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3775__B2 (.DIODE(\z80.tv80s.i_tv80_core.BusA[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3777__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusB[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3780__A2 (.DIODE(\z80.tv80s.di_reg[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3782__A (.DIODE(_0856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3783__A2 (.DIODE(_0856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3784__A (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__3785__C (.DIODE(_0398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3789__A2 (.DIODE(_0400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3790__A1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__3790__A2 (.DIODE(_0398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3791__A1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__3793__B (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__3793__C (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__3794__A (.DIODE(_0794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3794__B (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3795__B (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__3796__A (.DIODE(_0794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3796__B (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3796__C (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__3799__A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__3799__B (.DIODE(_0873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3800__A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__3800__B (.DIODE(_0873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3801__B (.DIODE(_0873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3802__B (.DIODE(_0873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3804__B (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3804__C (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__3805__A (.DIODE(_0794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3805__B (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__3806__B (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__3807__A (.DIODE(_0794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3807__B (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3807__C (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__3808__A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__3810__A (.DIODE(_0794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3810__B (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3816__C (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__3817__B (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__3817__C (.DIODE(_0873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3818__C (.DIODE(_0873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3819__A2 (.DIODE(_0868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3820__A2 (.DIODE(_0879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3820__B1 (.DIODE(_0882_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3821__A2 (.DIODE(_0806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3821__B1 (.DIODE(_0885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3824__A2 (.DIODE(_0868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3824__B1 (.DIODE(_0870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3827__A1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__3827__B1 (.DIODE(_0794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3828__A1 (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3829__A2 (.DIODE(_0806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3829__B1 (.DIODE(_0879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3834__A2 (.DIODE(_0874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3834__B1 (.DIODE(_0876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3835__A2 (.DIODE(_0868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3835__B1 (.DIODE(_0870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3836__A2 (.DIODE(_0879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3836__B1 (.DIODE(_0882_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3837__A2 (.DIODE(_0806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3837__B1 (.DIODE(_0885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3840__A2 (.DIODE(_0868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3840__B1 (.DIODE(_0870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3843__A1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__3843__B1 (.DIODE(_0794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3844__A1 (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3845__A2 (.DIODE(_0806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3845__B1 (.DIODE(_0879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3849__A2 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__3849__C1 (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3851__A2 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__3851__C1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__3852__A (.DIODE(_0794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3855__S (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3862__S (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3864__A (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3866__A1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__3866__B1 (.DIODE(_0794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3869__S (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__3871__C1 (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3872__C1 (.DIODE(_0794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3874__S (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__3876__A1 (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3881__S (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__3882__S (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__3883__S (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3884__S (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__3885__A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__3887__A1 (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3887__B1 (.DIODE(_0794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3905__A2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__3905__B1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__3906__A (.DIODE(\z80.tv80s.i_tv80_core.RegAddrB_r[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3906__B (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__3907__B (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__3908__A2 (.DIODE(_0772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3909__A2 (.DIODE(_0772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3910__S1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__3911__B2 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__3912__S (.DIODE(_0808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3913__A_N (.DIODE(\z80.tv80s.i_tv80_core.BusB[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3913__B (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__3914__A_N (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__3914__B (.DIODE(\z80.tv80s.i_tv80_core.BusB[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3915__B1 (.DIODE(\z80.tv80s.i_tv80_core.BusA[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3917__A (.DIODE(\z80.tv80s.i_tv80_core.BusA[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3924__A2 (.DIODE(\z80.tv80s.i_tv80_core.BusA[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3924__A3 (.DIODE(\z80.tv80s.i_tv80_core.BusB[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3925__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusB[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3925__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusB[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3926__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusA[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3926__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusA[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3929__B1 (.DIODE(\z80.tv80s.i_tv80_core.BusB[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3932__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusA[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3932__A2 (.DIODE(\z80.tv80s.i_tv80_core.BusA[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3932__B1 (.DIODE(\z80.tv80s.i_tv80_core.BusA[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3933__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusA[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3933__A2 (.DIODE(\z80.tv80s.i_tv80_core.BusA[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3933__B1 (.DIODE(\z80.tv80s.i_tv80_core.BusA[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3934__A (.DIODE(\z80.tv80s.i_tv80_core.F[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3935__A (.DIODE(\z80.tv80s.i_tv80_core.BusA[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3935__B (.DIODE(\z80.tv80s.i_tv80_core.F[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3936__S (.DIODE(\z80.tv80s.i_tv80_core.BusA[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3939__A0 (.DIODE(_2871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3941__A (.DIODE(_1014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3942__A2 (.DIODE(_1014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3943__A2 (.DIODE(_0874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3943__B1 (.DIODE(_0876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3944__A2 (.DIODE(_0868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3944__B1 (.DIODE(_0870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3945__A2 (.DIODE(_0879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3945__B1 (.DIODE(_0882_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3946__A2 (.DIODE(_0806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3946__B1 (.DIODE(_0885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3952__A2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__3952__B1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__3953__S0 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__3954__B2 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__3955__S (.DIODE(_0808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3956__S0 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__3957__A2 (.DIODE(_0874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3957__B1 (.DIODE(_0876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3958__A2 (.DIODE(_0868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3958__B1 (.DIODE(_0870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3959__A2 (.DIODE(_0879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3959__B1 (.DIODE(_0882_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3960__A2 (.DIODE(_0806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3960__B1 (.DIODE(_0885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3968__B (.DIODE(\z80.tv80s.i_tv80_core.BusB[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3969__A (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__3970__B1 (.DIODE(\z80.tv80s.i_tv80_core.BusA[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3972__A (.DIODE(\z80.tv80s.i_tv80_core.BusA[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3980__A0 (.DIODE(\z80.tv80s.i_tv80_core.F[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3981__A (.DIODE(\z80.tv80s.i_tv80_core.BusA[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3981__B (.DIODE(\z80.tv80s.i_tv80_core.BusA[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3983__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusB[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3983__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusB[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3984__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusA[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3984__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusA[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3984__S (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__3989__B2 (.DIODE(\z80.tv80s.i_tv80_core.BusB[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3992__A2 (.DIODE(\z80.tv80s.di_reg[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3994__A (.DIODE(_1066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3995__A2 (.DIODE(_1066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3997__A2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__3998__S (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__3999__S (.DIODE(_0808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4000__B (.DIODE(\z80.tv80s.i_tv80_core.BusB[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4001__B (.DIODE(\z80.tv80s.i_tv80_core.BusB[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4002__B1 (.DIODE(\z80.tv80s.i_tv80_core.BusA[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4003__A (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__4004__A (.DIODE(\z80.tv80s.i_tv80_core.BusA[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4011__A2 (.DIODE(\z80.tv80s.i_tv80_core.BusA[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4011__A3 (.DIODE(\z80.tv80s.i_tv80_core.BusB[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4012__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusA[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4012__A2 (.DIODE(\z80.tv80s.i_tv80_core.BusA[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4012__B1 (.DIODE(\z80.tv80s.i_tv80_core.BusA[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4013__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusA[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4013__A2 (.DIODE(\z80.tv80s.i_tv80_core.BusA[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4013__A3 (.DIODE(\z80.tv80s.i_tv80_core.BusA[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4014__A (.DIODE(\z80.tv80s.i_tv80_core.BusA[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4014__B (.DIODE(\z80.tv80s.i_tv80_core.BusA[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4014__C (.DIODE(\z80.tv80s.i_tv80_core.BusA[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4015__B1 (.DIODE(\z80.tv80s.i_tv80_core.F[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4017__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4018__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusB[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4018__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusB[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4019__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusA[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4019__S (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__4022__A (.DIODE(\z80.tv80s.i_tv80_core.BusB[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4024__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusB[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4026__A0 (.DIODE(\z80.tv80s.di_reg[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4029__A (.DIODE(_1100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4030__A2 (.DIODE(_1100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4031__A2 (.DIODE(_0868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4031__B1 (.DIODE(_0870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4032__A2 (.DIODE(_0874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4032__B1 (.DIODE(_0876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4033__A2 (.DIODE(_0879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4033__B1 (.DIODE(_0882_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4034__A2 (.DIODE(_0806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4034__B1 (.DIODE(_0885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4036__B (.DIODE(_1107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4040__A2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__4040__B1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__4041__S0 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__4041__S1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__4042__B2 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__4043__S (.DIODE(_0808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4044__A4 (.DIODE(_1107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4047__A2 (.DIODE(_0868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4047__B1 (.DIODE(_0870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4048__A2 (.DIODE(_0874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4048__B1 (.DIODE(_0876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4049__A2 (.DIODE(_0879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4049__B1 (.DIODE(_0882_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4050__A2 (.DIODE(_0806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4050__B1 (.DIODE(_0885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4054__A (.DIODE(\z80.tv80s.i_tv80_core.F[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4054__B (.DIODE(\z80.tv80s.i_tv80_core.F[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4055__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4058__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusA[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4058__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusA[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4058__S (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__4059__B (.DIODE(\z80.tv80s.i_tv80_core.BusB[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4061__B (.DIODE(\z80.tv80s.i_tv80_core.BusB[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4075__B2 (.DIODE(\z80.tv80s.i_tv80_core.BusB[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4077__A0 (.DIODE(\z80.tv80s.di_reg[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4080__A (.DIODE(_1150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4081__A2 (.DIODE(_1150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4081__B1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__4083__A2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__4083__B1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__4084__S0 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__4085__B2 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__4086__S (.DIODE(_0808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4088__B (.DIODE(\z80.tv80s.i_tv80_core.BusB[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4089__B (.DIODE(\z80.tv80s.i_tv80_core.BusB[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4090__B1 (.DIODE(\z80.tv80s.i_tv80_core.BusA[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4091__A (.DIODE(\z80.tv80s.i_tv80_core.BusA[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4096__A (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__4099__A2 (.DIODE(\z80.tv80s.i_tv80_core.BusA[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4099__A3 (.DIODE(\z80.tv80s.i_tv80_core.BusB[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4101__A (.DIODE(\z80.tv80s.i_tv80_core.BusA[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4102__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusA[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4102__A2 (.DIODE(\z80.tv80s.i_tv80_core.BusA[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4102__B1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__4103__A (.DIODE(\z80.tv80s.i_tv80_core.F[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4104__A (.DIODE(\z80.tv80s.i_tv80_core.F[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4105__B (.DIODE(\z80.tv80s.i_tv80_core.BusA[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4108__A (.DIODE(\z80.tv80s.i_tv80_core.BusA[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4109__A (.DIODE(\z80.tv80s.i_tv80_core.BusA[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4110__S (.DIODE(\z80.tv80s.i_tv80_core.F[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4113__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusA[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4114__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusA[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4114__S (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__4118__B2 (.DIODE(\z80.tv80s.i_tv80_core.BusB[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4120__A0 (.DIODE(\z80.tv80s.di_reg[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4122__A (.DIODE(_1191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4123__A2 (.DIODE(_1191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4123__B1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__4124__A2 (.DIODE(_0868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4124__B1 (.DIODE(_0870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4125__A2 (.DIODE(_0874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4125__B1 (.DIODE(_0876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4126__A2 (.DIODE(_0879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4126__B1 (.DIODE(_0882_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4127__A2 (.DIODE(_0806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4127__B1 (.DIODE(_0885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4129__B (.DIODE(_1198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4131__B (.DIODE(_1198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4136__A2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__4136__B1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__4137__S0 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__4137__S1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__4138__B2 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__4139__S (.DIODE(_0808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4140__A2 (.DIODE(_0868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4140__B1 (.DIODE(_0870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4141__A2 (.DIODE(_0874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4141__B1 (.DIODE(_0876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4142__A2 (.DIODE(_0879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4142__B1 (.DIODE(_0882_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4143__A2 (.DIODE(_0806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4143__B1 (.DIODE(_0885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4150__A (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__4150__B (.DIODE(\z80.tv80s.i_tv80_core.BusB[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4151__A (.DIODE(\z80.tv80s.i_tv80_core.BusA[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4152__A (.DIODE(\z80.tv80s.i_tv80_core.BusA[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4159__A2 (.DIODE(\z80.tv80s.i_tv80_core.BusA[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4159__A3 (.DIODE(\z80.tv80s.i_tv80_core.BusB[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4160__A (.DIODE(\z80.tv80s.i_tv80_core.BusA[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4164__A (.DIODE(\z80.tv80s.i_tv80_core.BusA[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4167__S (.DIODE(\z80.tv80s.i_tv80_core.F[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4168__A (.DIODE(_0405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4169__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusA[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4169__A1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__4169__S (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__4170__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusA[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4171__A1 (.DIODE(_0405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4172__A1 (.DIODE(_0405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4172__B2 (.DIODE(\z80.tv80s.i_tv80_core.BusB[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4175__A2 (.DIODE(\z80.tv80s.di_reg[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4177__A (.DIODE(_1245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4178__B (.DIODE(_1245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4179__C1 (.DIODE(_0774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4180__A2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__4180__B1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__4181__S0 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__4181__S1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__4182__B2 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__4183__S (.DIODE(_0808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4185__A2 (.DIODE(_0874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4185__B1 (.DIODE(_0876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4186__A2 (.DIODE(_0868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4186__B1 (.DIODE(_0870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4187__A2 (.DIODE(_0879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4187__B1 (.DIODE(_0882_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4188__A2 (.DIODE(_0806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4188__B1 (.DIODE(_0885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4193__A (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__4194__B (.DIODE(\z80.tv80s.i_tv80_core.BusB[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4197__A (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__4197__B (.DIODE(\z80.tv80s.i_tv80_core.BusB[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4198__A (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__4198__B (.DIODE(\z80.tv80s.i_tv80_core.BusB[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4202__A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__4202__A3 (.DIODE(\z80.tv80s.i_tv80_core.BusB[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4204__A (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__4204__B (.DIODE(\z80.tv80s.i_tv80_core.BusA[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4205__A0 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__4207__A (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__4207__B (.DIODE(\z80.tv80s.i_tv80_core.BusA[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4208__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusA[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4214__S (.DIODE(\z80.tv80s.i_tv80_core.F[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4217__B (.DIODE(\z80.tv80s.i_tv80_core.BusA[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4218__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__4218__A2 (.DIODE(\z80.tv80s.i_tv80_core.BusA[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4219__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4219__B2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__4220__A (.DIODE(\z80.tv80s.i_tv80_core.BusB[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4220__B (.DIODE(_0474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4222__A (.DIODE(\z80.tv80s.i_tv80_core.BusB[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4222__B (.DIODE(_0474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4226__A0 (.DIODE(\z80.tv80s.di_reg[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4228__A2 (.DIODE(_1295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4228__B1 (.DIODE(_0774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4230__A2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__4230__B1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__4231__B (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__4232__B (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__4233__B (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__4233__C (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__4234__A2 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__4234__B1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__4236__A2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__4236__C1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__4237__A2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__4237__C1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__4238__A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__4238__C1 (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4239__A1 (.DIODE(_1300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4240__B2 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__4241__S (.DIODE(_0808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4242__A (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__4243__A1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__4243__B1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__4245__A1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__4246__B (.DIODE(_0477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4248__A (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4248__C (.DIODE(_2982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4254__A1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__4254__A2 (.DIODE(_0397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4256__A1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__4257__A3 (.DIODE(_0398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4258__A1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__4258__A2 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__4258__C1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__4259__B (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__4259__C (.DIODE(_2849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4262__A_N (.DIODE(_2999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4264__A (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__4265__A1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__4267__A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__4268__A (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__4270__B1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__4272__A1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__4273__A (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__4274__A1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__4274__B1 (.DIODE(_0684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4274__C1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__4275__A1 (.DIODE(_2934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4275__A3 (.DIODE(_0398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4276__A (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__4276__B (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__4278__C1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__4279__A1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__4279__A2 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__4279__B1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__4280__A1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__4280__B2 (.DIODE(_2934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4283__A (.DIODE(_1349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4284__C (.DIODE(_1349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4285__B (.DIODE(_1333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4287__S (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__4288__A (.DIODE(_2998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4289__A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__4289__B (.DIODE(_2998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4290__A (.DIODE(_2846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4290__B (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__4290__C (.DIODE(_1355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4291__A (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__4291__B (.DIODE(_2854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4291__C_N (.DIODE(_1355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4292__A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__4292__C (.DIODE(_0603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4293__A2 (.DIODE(_0607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4293__B1 (.DIODE(_1357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4294__B1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4294__B2 (.DIODE(_1356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4295__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__4297__B1 (.DIODE(_1356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4298__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4298__A2 (.DIODE(_1356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4299__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__4300__A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__4301__A0 (.DIODE(\z80.tv80s.i_tv80_core.ACC[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4301__S (.DIODE(_1357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4304__A1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__4304__A2 (.DIODE(_0603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4305__B (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__4305__C (.DIODE(_0603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4306__A1 (.DIODE(_1357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4306__B1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__4307__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4307__A2 (.DIODE(_1356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4308__A1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__4310__A0 (.DIODE(\z80.tv80s.i_tv80_core.ACC[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4310__S (.DIODE(_1357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4311__B2 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__4312__C (.DIODE(_0603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4313__A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__4314__A1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__4315__A (.DIODE(_1356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4316__A2 (.DIODE(_1357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4317__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__4318__A1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__4319__A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__4319__C (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__4321__B1 (.DIODE(_1356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4322__A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__4322__B (.DIODE(_1356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4323__A1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__4323__B2 (.DIODE(\z80.tv80s.i_tv80_core.ACC[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4324__B (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__4325__A (.DIODE(_2849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4326__A1 (.DIODE(_0450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4327__A1 (.DIODE(_2847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4329__A2 (.DIODE(_0401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4329__B2 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__4330__A1 (.DIODE(_0401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4330__B1 (.DIODE(_0684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4330__B2 (.DIODE(_2847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4331__A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__4331__B (.DIODE(_2847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4332__B (.DIODE(_0405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4334__A2 (.DIODE(_3021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4335__A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__4336__A1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__4337__A1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__4337__C1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__4339__A1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__4339__A2 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__4341__A1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__4342__B2 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__4343__A1 (.DIODE(_2934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4343__A2 (.DIODE(_0684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4345__C1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__4346__A2 (.DIODE(_0401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4346__B2 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__4347__A1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__4347__A3 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__4350__B2 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__4351__A1 (.DIODE(_2934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4352__A1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__4353__A1_N (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4353__B2 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__4354__C (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4354__D_N (.DIODE(_1412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4356__S (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__4360__A (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__4361__A (.DIODE(_1415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4361__B (.DIODE(_1417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4362__A1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__4362__B1 (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA__4363__A (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA__4365__A0 (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA__4365__S (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__4366__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__4367__A1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__4367__A2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__4369__S (.DIODE(_1424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4370__S (.DIODE(_1424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4371__S (.DIODE(_1424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4372__S (.DIODE(_1424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4373__S (.DIODE(_1424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4374__S (.DIODE(_1424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4375__S (.DIODE(_1424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4376__S (.DIODE(_1424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4378__S (.DIODE(_1425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4379__S (.DIODE(_1425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4380__S (.DIODE(_1425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4381__S (.DIODE(_1425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4382__S (.DIODE(_1425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4383__S (.DIODE(_1425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4384__S (.DIODE(_1425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4385__S (.DIODE(_1425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4387__A1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__4388__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__4390__S (.DIODE(_1428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4391__S (.DIODE(_1428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4392__S (.DIODE(_1428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4393__S (.DIODE(_1428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4394__S (.DIODE(_1428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4395__S (.DIODE(_1428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4396__S (.DIODE(_1428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4397__S (.DIODE(_1428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4398__C_N (.DIODE(_0781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4399__B1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__4402__A2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__4403__S1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__4404__A1 (.DIODE(_0772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4405__S (.DIODE(_1431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4406__B (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__4406__C (.DIODE(_0772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4407__A2 (.DIODE(_0981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4407__B1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__4408__S (.DIODE(_0981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4409__A2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__4409__C1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__4410__A2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__4410__C1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__4411__A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__4411__C1 (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4412__A1 (.DIODE(_1300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4415__A2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__4416__A1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__4417__S (.DIODE(_1431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4418__B (.DIODE(\z80.tv80s.i_tv80_core.RegAddrB_r[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4418__C (.DIODE(_0772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4419__A2 (.DIODE(_0981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4419__B1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__4421__A2 (.DIODE(\z80.tv80s.i_tv80_core.RegAddrB_r[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4421__B1 (.DIODE(_0981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4421__C1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__4422__A2 (.DIODE(\z80.tv80s.i_tv80_core.RegAddrB_r[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4422__C1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__4423__A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__4423__C1 (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4424__A1 (.DIODE(_1300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4428__A1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__4429__S (.DIODE(_1431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4434__S0 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__4435__B2 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__4436__S (.DIODE(_1431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4439__B2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__4440__S0 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__4440__S1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__4441__S (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__4442__S (.DIODE(_1431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4446__A2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__4446__B1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__4447__S0 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__4447__S1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__4448__B2 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__4449__S (.DIODE(_1431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4453__C1 (.DIODE(_0774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4454__A2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__4454__B1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__4455__S0 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__4456__B2 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__4457__S (.DIODE(_1431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4458__S0 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__4462__A2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__4463__S (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__4464__S (.DIODE(_1431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4466__S (.DIODE(_1488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4467__S (.DIODE(_1488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4468__S (.DIODE(_1488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4469__S (.DIODE(_1488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4470__S (.DIODE(_1488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4471__S (.DIODE(_1488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4472__S (.DIODE(_1488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4473__S (.DIODE(_1488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4475__S (.DIODE(_1489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4476__S (.DIODE(_1489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4477__S (.DIODE(_1489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4478__S (.DIODE(_1489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4479__S (.DIODE(_1489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4480__S (.DIODE(_1489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4481__S (.DIODE(_1489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4482__S (.DIODE(_1489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4484__S (.DIODE(_1490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4485__S (.DIODE(_1490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4486__S (.DIODE(_1490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4487__S (.DIODE(_1490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4488__S (.DIODE(_1490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4489__S (.DIODE(_1490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4490__S (.DIODE(_1490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4491__S (.DIODE(_1490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4493__S (.DIODE(_1491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4494__S (.DIODE(_1491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4495__S (.DIODE(_1491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4496__S (.DIODE(_1491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4497__S (.DIODE(_1491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4498__S (.DIODE(_1491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4499__S (.DIODE(_1491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4500__S (.DIODE(_1491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4502__S (.DIODE(_1492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4503__S (.DIODE(_1492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4504__S (.DIODE(_1492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4505__S (.DIODE(_1492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4506__S (.DIODE(_1492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4507__S (.DIODE(_1492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4508__S (.DIODE(_1492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4509__S (.DIODE(_1492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4511__S (.DIODE(_1493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4512__S (.DIODE(_1493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4513__S (.DIODE(_1493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4514__S (.DIODE(_1493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4515__S (.DIODE(_1493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4516__S (.DIODE(_1493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4517__S (.DIODE(_1493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4518__S (.DIODE(_1493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4520__S (.DIODE(_1494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4521__S (.DIODE(_1494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4522__S (.DIODE(_1494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4523__S (.DIODE(_1494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4524__S (.DIODE(_1494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4525__S (.DIODE(_1494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4526__S (.DIODE(_1494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4527__S (.DIODE(_1494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4529__S (.DIODE(_1495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4530__S (.DIODE(_1495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4531__S (.DIODE(_1495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4532__S (.DIODE(_1495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4533__S (.DIODE(_1495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4534__S (.DIODE(_1495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4535__S (.DIODE(_1495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4536__S (.DIODE(_1495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4538__S (.DIODE(_1496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4539__S (.DIODE(_1496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4540__S (.DIODE(_1496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4541__S (.DIODE(_1496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4542__S (.DIODE(_1496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4543__S (.DIODE(_1496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4544__S (.DIODE(_1496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4545__S (.DIODE(_1496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4547__S (.DIODE(_1497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4548__S (.DIODE(_1497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4549__S (.DIODE(_1497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4550__S (.DIODE(_1497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4551__S (.DIODE(_1497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4552__S (.DIODE(_1497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4553__S (.DIODE(_1497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4554__S (.DIODE(_1497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4555__A (.DIODE(\z80.tv80s.i_tv80_core.ISet[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4555__B (.DIODE(_2952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4556__A (.DIODE(\z80.tv80s.i_tv80_core.ISet[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4556__B (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__4556__C (.DIODE(_2952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4556__D (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__4557__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__4557__C (.DIODE(_2899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4558__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__4559__A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__4560__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4561__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4562__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4563__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4564__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4565__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4566__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4567__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4568__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4569__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4570__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4571__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4572__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4573__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4574__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4575__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4576__A1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__4576__B1 (.DIODE(_2999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4577__B (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__4577__C (.DIODE(_0398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4578__A1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__4578__A2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__4579__B2 (.DIODE(\z80.tv80s.i_tv80_core.ISet[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4580__B2 (.DIODE(\z80.tv80s.i_tv80_core.ISet[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4581__A1 (.DIODE(_1333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4581__A2 (.DIODE(_1349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4582__A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__4583__A1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__4583__A2 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__4583__A3 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__4584__A1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__4584__A2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__4586__C1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__4589__A2 (.DIODE(_0554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4590__A1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__4590__B2 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__4591__A1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__4592__C1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__4593__A1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__4594__B (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__4595__B (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__4596__B2 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__4597__B1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__4598__A1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__4598__A2 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__4599__A1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__4599__A2 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__4600__B (.DIODE(_1525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4601__A (.DIODE(_1333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4601__B (.DIODE(_1349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4603__A2 (.DIODE(_1525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4604__A (.DIODE(_1333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4604__B (.DIODE(_1349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4604__D (.DIODE(_1525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4605__A (.DIODE(_1333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4605__B (.DIODE(_1349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4605__D (.DIODE(_1526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4606__A (.DIODE(_1525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4607__A (.DIODE(_1526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4608__A1 (.DIODE(\z80.tv80s.di_reg[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4608__B2 (.DIODE(\z80.tv80s.i_tv80_core.ACC[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4610__A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__4611__B (.DIODE(_1526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4612__A2 (.DIODE(_1526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4613__A1 (.DIODE(\z80.tv80s.di_reg[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4613__B2 (.DIODE(\z80.tv80s.i_tv80_core.ACC[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4616__S (.DIODE(_1525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4617__A1 (.DIODE(\z80.tv80s.di_reg[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4617__B2 (.DIODE(\z80.tv80s.i_tv80_core.ACC[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4620__B2 (.DIODE(_1544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4621__A1 (.DIODE(_1107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4621__S (.DIODE(_1525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4622__A1 (.DIODE(\z80.tv80s.di_reg[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4622__B2 (.DIODE(\z80.tv80s.i_tv80_core.ACC[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4625__A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__4625__B2 (.DIODE(_1548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4626__S (.DIODE(_1525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4627__A1 (.DIODE(\z80.tv80s.di_reg[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4627__B2 (.DIODE(\z80.tv80s.i_tv80_core.ACC[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4630__B2 (.DIODE(_1552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4631__A1 (.DIODE(_1198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4631__S (.DIODE(_1525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4632__A1 (.DIODE(\z80.tv80s.di_reg[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4632__B2 (.DIODE(\z80.tv80s.i_tv80_core.ACC[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4635__B2 (.DIODE(_1556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4636__B (.DIODE(_1525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4637__A2 (.DIODE(_1526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4638__A1 (.DIODE(\z80.tv80s.di_reg[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4638__B2 (.DIODE(\z80.tv80s.i_tv80_core.ACC[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4641__B (.DIODE(_1525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4642__A2 (.DIODE(_1526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4643__A1 (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA__4643__B2 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA__4645__A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__4647__A2 (.DIODE(_1565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4648__A1 (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA__4649__A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__4650__A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__4650__B (.DIODE(_1567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4651__A1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__4651__A2 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__4651__B1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__4652__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__4652__B (.DIODE(_0603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4653__A (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA__4654__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__4654__B1 (.DIODE(_1570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4655__A1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__4655__A2 (.DIODE(_1570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4656__A (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__4656__B (.DIODE(_1567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4657__A1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__4657__A2 (.DIODE(_1570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4658__A (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__4658__B (.DIODE(_1567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4659__A2 (.DIODE(_1570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4660__A (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__4660__B (.DIODE(_1567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4661__A2 (.DIODE(_1570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4662__A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__4662__B (.DIODE(_1567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4663__A2 (.DIODE(_1570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4664__A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__4664__B (.DIODE(_1567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4665__A2 (.DIODE(_1570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4666__A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__4666__B (.DIODE(_1567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4667__A2 (.DIODE(_1570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4668__A (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__4668__B (.DIODE(_1567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4669__A2 (.DIODE(_1570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4670__C (.DIODE(_0781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4672__A1 (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4672__A2 (.DIODE(_1581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4672__B1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__4673__A (.DIODE(_0856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4673__B (.DIODE(_1581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4674__B (.DIODE(_0554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4675__A (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__4677__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusB[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4677__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusA[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4677__S (.DIODE(_1586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4678__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusB[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4678__S (.DIODE(_1585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4679__A1 (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4679__B1 (.DIODE(_1581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4680__A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__4681__A (.DIODE(_1014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4681__B (.DIODE(_1581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4682__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusB[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4682__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusA[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4682__S (.DIODE(_1586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4683__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusB[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4683__S (.DIODE(_1585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4684__A1 (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4684__B1 (.DIODE(_1581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4685__A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__4686__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusB[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4686__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusA[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4686__S (.DIODE(_1586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4687__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusB[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4687__S (.DIODE(_1585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4688__A (.DIODE(_1066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4688__B (.DIODE(_1581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4689__A1 (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4689__B1 (.DIODE(_1581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4690__A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__4691__A (.DIODE(_1100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4691__B (.DIODE(_1581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4692__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusB[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4692__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusA[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4692__S (.DIODE(_1586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4693__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusB[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4693__S (.DIODE(_1585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4694__A1 (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4694__B1 (.DIODE(_1581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4695__A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__4696__A (.DIODE(_1150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4696__B (.DIODE(_1581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4697__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusB[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4697__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusB[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4697__S (.DIODE(_1586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4698__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusA[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4698__S (.DIODE(_1585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4699__A1 (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4699__B1 (.DIODE(_1581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4700__A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__4701__A (.DIODE(_1191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4701__B (.DIODE(_1581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4702__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusB[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4702__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusB[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4702__S (.DIODE(_1586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4703__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusA[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4703__S (.DIODE(_1585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4704__A1 (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4704__B1 (.DIODE(_1581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4705__A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__4706__A (.DIODE(_1245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4706__B (.DIODE(_1581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4707__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusB[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4707__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusB[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4707__S (.DIODE(_1586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4708__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusA[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4708__S (.DIODE(_1585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4709__A1 (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4709__B1 (.DIODE(_1581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4710__A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__4711__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusB[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4711__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusB[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4711__S (.DIODE(_1586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4712__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusA[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4712__S (.DIODE(_1585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4713__A (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4714__A0 (.DIODE(_1295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4714__S (.DIODE(_1581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4715__B2 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__4716__A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__4716__B (.DIODE(_2846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4716__C (.DIODE(\z80.tv80s.i_tv80_core.ISet[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4716__D (.DIODE(_2929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4717__A (.DIODE(_0577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4718__B1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__4720__A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__4720__D (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__4721__B1 (.DIODE(_1622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4722__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4722__B2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__4723__A (.DIODE(_2846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4723__B (.DIODE(_2854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4724__A (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__4724__B (.DIODE(\z80.tv80s.i_tv80_core.ts[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4726__S (.DIODE(_1355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4727__S (.DIODE(_1626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4728__S (.DIODE(_1627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4729__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__4730__A1_N (.DIODE(\z80.tv80s.i_tv80_core.ACC[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4730__A2_N (.DIODE(_1622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4731__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4731__B2 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__4732__S (.DIODE(_1355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4733__S (.DIODE(_1626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4734__S (.DIODE(_1627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4735__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__4736__A1_N (.DIODE(\z80.tv80s.i_tv80_core.ACC[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4736__A2_N (.DIODE(_1622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4736__B1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__4737__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4737__B2 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__4738__S (.DIODE(_1355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4739__S (.DIODE(_1626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4740__S (.DIODE(_1627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4741__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__4742__A1_N (.DIODE(\z80.tv80s.i_tv80_core.ACC[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4742__A2_N (.DIODE(_1622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4743__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4743__B2 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__4744__S (.DIODE(_1355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4745__S (.DIODE(_1626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4746__S (.DIODE(_1627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4747__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__4748__A1_N (.DIODE(\z80.tv80s.i_tv80_core.ACC[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4748__A2_N (.DIODE(_1622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4748__B1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__4749__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4749__B2 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__4750__S (.DIODE(_1355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4751__S (.DIODE(_1626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4752__S (.DIODE(_1627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4753__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__4754__A1_N (.DIODE(\z80.tv80s.i_tv80_core.ACC[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4754__A2_N (.DIODE(_1622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4755__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4755__B2 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__4756__S (.DIODE(_1355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4757__S (.DIODE(_1626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4758__S (.DIODE(_1627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4759__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__4760__A1_N (.DIODE(\z80.tv80s.i_tv80_core.ACC[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4760__A2_N (.DIODE(_1622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4761__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4761__B2 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__4762__S (.DIODE(_1355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4763__S (.DIODE(_1626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4764__S (.DIODE(_1627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4765__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__4766__A1_N (.DIODE(\z80.tv80s.i_tv80_core.ACC[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4766__A2_N (.DIODE(_1622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4767__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4767__B2 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__4768__A0 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA__4768__S (.DIODE(_1355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4769__S (.DIODE(_1626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4770__A0 (.DIODE(_1295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4770__S (.DIODE(_1627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4771__A0 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA__4771__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__4772__A1 (.DIODE(_0577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4772__A2 (.DIODE(_0598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4772__B1 (.DIODE(_0605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4773__A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__4775__A1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__4775__A2 (.DIODE(_1668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4776__A1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__4776__A2 (.DIODE(_1668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4777__S0 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__4777__S1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__4778__S0 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__4778__S1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__4779__S (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA__4780__A2 (.DIODE(_1673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4780__B1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__4781__A1 (.DIODE(_2899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4782__A (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__4783__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__4783__B (.DIODE(_0653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4786__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__4788__B (.DIODE(_0717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4789__B (.DIODE(_1682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4790__A (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4790__B (.DIODE(\z80.tv80s.i_tv80_core.IntCycle ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4791__A (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4791__B (.DIODE(\z80.tv80s.i_tv80_core.IntCycle ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4793__A (.DIODE(_1686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4796__A (.DIODE(_1689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4798__A1 (.DIODE(_1673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4798__B1 (.DIODE(_1691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4798__B2 (.DIODE(\z80.tv80s.di_reg[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4800__S (.DIODE(_0502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4801__A0 (.DIODE(_1673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4801__S (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__4804__A_N (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__4804__B_N (.DIODE(_0554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4808__A (.DIODE(_1701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4809__B (.DIODE(_1701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4810__B (.DIODE(_1701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4811__A1 (.DIODE(_1696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4811__B2 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__4814__C1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__4815__A2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__4815__C1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__4816__A2 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__4818__A2 (.DIODE(_1684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4818__B1 (.DIODE(_1682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4819__S0 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__4819__S1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__4820__B (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA__4821__S0 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__4821__S1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__4822__A1 (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA__4823__A1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__4824__A (.DIODE(_1689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4824__B (.DIODE(_1716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4825__B1 (.DIODE(_1691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4825__B2 (.DIODE(\z80.tv80s.di_reg[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4826__S (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__4827__S (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__4828__C (.DIODE(_1701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4829__A2 (.DIODE(_1701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4831__A1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__4831__B2 (.DIODE(_1696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4835__B (.DIODE(_1716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4836__C1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__4838__B (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__4839__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__4841__A2 (.DIODE(_1684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4841__B1 (.DIODE(_1682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4842__S0 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__4842__S1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__4843__S0 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__4843__S1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__4844__S (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__4845__S (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__4846__A0 (.DIODE(_1736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4846__S (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__4848__B2 (.DIODE(_1736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4849__B1 (.DIODE(_1696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4851__A1 (.DIODE(\z80.tv80s.di_reg[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4851__A2 (.DIODE(_1691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4851__B2 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__4853__B (.DIODE(_1686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4857__A1 (.DIODE(_1417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4857__A2 (.DIODE(_1736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4858__A2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__4858__C1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__4859__A2 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__4861__S0 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__4861__S1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__4862__S0 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__4862__S1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__4863__S (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__4864__A1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__4864__A2 (.DIODE(_1754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4865__A (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4866__A (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4867__A (.DIODE(_1696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4868__A1 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4868__S (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__4869__A0 (.DIODE(_1754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4869__S (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__4870__B2 (.DIODE(_1754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4871__A1 (.DIODE(\z80.tv80s.di_reg[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4871__A2 (.DIODE(_1691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4872__A2 (.DIODE(_1686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4873__A0 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4874__A1 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4876__A1 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4876__B1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__4877__A2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__4879__S0 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__4879__S1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__4880__S0 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__4880__S1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__4881__S (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__4882__A1 (.DIODE(_1417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4882__A2 (.DIODE(_1771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4882__B1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__4883__A (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4883__B (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4884__A2 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4884__B1 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4885__C (.DIODE(_1696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4886__A1 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4886__S (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__4887__A0 (.DIODE(_1771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4887__S (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__4888__B2 (.DIODE(_1771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4889__A1 (.DIODE(\z80.tv80s.di_reg[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4889__A2 (.DIODE(_1691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4889__B2 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__4890__B (.DIODE(_1686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4892__A0 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4893__A1 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4893__A2 (.DIODE(_1681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4895__A1 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4895__B1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__4896__A2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__4898__S0 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__4898__S1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__4899__S0 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__4899__S1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__4900__S (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__4901__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__4901__B (.DIODE(_1789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4902__A1 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4902__A2 (.DIODE(_1684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4902__B1 (.DIODE(_1682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4903__A1 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4903__S (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__4904__A0 (.DIODE(_1789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4904__S (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__4905__A (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4906__B2 (.DIODE(_1789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4907__A1 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4907__B1 (.DIODE(_1696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4908__A1 (.DIODE(\z80.tv80s.di_reg[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4908__A2 (.DIODE(_1691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4908__B2 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__4910__B (.DIODE(_1686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4912__A1 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4914__A0 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4915__S (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__4917__S1 (.DIODE(\z80.tv80s.i_tv80_core.RegAddrC[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4918__S1 (.DIODE(\z80.tv80s.i_tv80_core.RegAddrC[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4919__S (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA__4920__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__4920__B (.DIODE(_1807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4921__A1 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4921__A2 (.DIODE(_1684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4921__B1 (.DIODE(_1682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4922__A (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4922__B (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4923__A1 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4923__B1 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4924__C (.DIODE(_1696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4925__A1 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4925__S (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__4926__A0 (.DIODE(_1807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4926__S (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__4927__B2 (.DIODE(_1807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4928__A1 (.DIODE(\z80.tv80s.di_reg[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4928__A2 (.DIODE(_1691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4928__B2 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__4930__B (.DIODE(_1686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4932__A1 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4934__A0 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4935__S (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__4937__S0 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__4937__S1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__4938__B (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__4939__S0 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__4939__S1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__4940__A1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__4941__A (.DIODE(_1827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4942__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__4943__A (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4943__B (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4943__C (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4943__D (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4944__D (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4946__A1 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4946__C1 (.DIODE(_1696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4947__A1 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4947__S (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__4948__S (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__4949__A (.DIODE(_1689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4949__B (.DIODE(_1827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4950__B1 (.DIODE(_1691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4950__B2 (.DIODE(\z80.tv80s.di_reg[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4951__A1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__4953__A0 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4954__A1 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4956__A0 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4956__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__4957__S (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__4959__S0 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__4959__S1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__4960__S0 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__4960__S1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__4961__S (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__4962__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__4962__B (.DIODE(_1847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4963__A (.DIODE(\z80.tv80s.i_tv80_core.ACC[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4963__B (.DIODE(_1691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4964__B2 (.DIODE(_1847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4965__A0 (.DIODE(\z80.tv80s.i_tv80_core.PC[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4965__S (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__4966__A0 (.DIODE(_1847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4970__A0 (.DIODE(\z80.tv80s.di_reg[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4970__S (.DIODE(_1701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4971__A1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__4971__B2 (.DIODE(_1696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4972__A1 (.DIODE(\z80.tv80s.i_tv80_core.PC[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4976__A0 (.DIODE(\z80.tv80s.di_reg[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4976__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__4977__S (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__4979__S0 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__4979__S1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__4980__S0 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__4980__S1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__4981__S (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__4982__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__4982__B (.DIODE(_1866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4983__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4983__A2 (.DIODE(_1691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4983__B1 (.DIODE(_1866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4985__A0 (.DIODE(\z80.tv80s.i_tv80_core.PC[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4985__S (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__4986__A0 (.DIODE(_1866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4989__B1 (.DIODE(_1701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4990__A1 (.DIODE(_2871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4991__A1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__4991__B2 (.DIODE(_1696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4992__A1 (.DIODE(\z80.tv80s.i_tv80_core.PC[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4996__A0 (.DIODE(\z80.tv80s.di_reg[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4996__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__4997__S (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__4999__S0 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__4999__S1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__5000__S0 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__5000__S1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5001__S (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__5002__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__5002__B (.DIODE(_1885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5003__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5003__A2 (.DIODE(_1691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5003__B1 (.DIODE(_1885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5005__A0 (.DIODE(\z80.tv80s.i_tv80_core.PC[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5005__S (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__5006__A0 (.DIODE(_1885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5008__A0 (.DIODE(\z80.tv80s.di_reg[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5008__S (.DIODE(_1701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5009__A1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__5009__B2 (.DIODE(_1696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5010__A1 (.DIODE(\z80.tv80s.i_tv80_core.PC[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5013__A1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__5014__A (.DIODE(\z80.tv80s.di_reg[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5014__B (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__5015__A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__5016__S (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__5018__S0 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__5018__S1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__5019__S0 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__5019__S1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__5020__S (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__5021__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__5021__B (.DIODE(_1903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5022__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5022__A2 (.DIODE(_1691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5022__B1 (.DIODE(_1903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5024__A0 (.DIODE(\z80.tv80s.i_tv80_core.PC[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5024__S (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__5025__A0 (.DIODE(_1903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5029__A0 (.DIODE(\z80.tv80s.di_reg[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5029__S (.DIODE(_1701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5030__A1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__5030__B2 (.DIODE(_1696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5031__A1 (.DIODE(\z80.tv80s.i_tv80_core.PC[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5035__A0 (.DIODE(\z80.tv80s.di_reg[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5035__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__5036__S (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__5038__S0 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__5038__S1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5039__S0 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__5039__S1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5040__S (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__5041__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__5041__B (.DIODE(_1922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5042__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5042__A2 (.DIODE(_1691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5042__B1 (.DIODE(_1922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5044__A0 (.DIODE(\z80.tv80s.i_tv80_core.PC[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5044__S (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__5045__A0 (.DIODE(_1922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5048__B1 (.DIODE(_1701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5049__A1 (.DIODE(\z80.tv80s.di_reg[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5049__A2 (.DIODE(_1701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5050__A1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__5050__B2 (.DIODE(_1696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5051__A1 (.DIODE(\z80.tv80s.i_tv80_core.PC[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5055__A0 (.DIODE(\z80.tv80s.di_reg[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5055__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__5056__S (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__5058__S0 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__5058__S1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__5059__B (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__5060__S0 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__5060__S1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__5061__A1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__5062__A (.DIODE(_1942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5063__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__5064__A (.DIODE(_1689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5064__B (.DIODE(_1942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5065__B1 (.DIODE(_1691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5065__B2 (.DIODE(\z80.tv80s.i_tv80_core.ACC[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5066__A0 (.DIODE(\z80.tv80s.i_tv80_core.PC[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5066__S (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__5069__A0 (.DIODE(\z80.tv80s.di_reg[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5069__S (.DIODE(_1701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5070__A1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__5070__B2 (.DIODE(_1696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5071__A1 (.DIODE(\z80.tv80s.i_tv80_core.PC[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5072__A0 (.DIODE(\z80.tv80s.i_tv80_core.I[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5075__A0 (.DIODE(\z80.tv80s.di_reg[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5075__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__5076__A0 (.DIODE(\z80.tv80s.i_tv80_core.I[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5076__S (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__5078__S0 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__5078__S1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5079__S0 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__5079__S1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__5080__S (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__5081__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__5081__B (.DIODE(_1960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5082__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5082__A2 (.DIODE(_1691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5082__B1 (.DIODE(_1960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5084__S (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__5085__A0 (.DIODE(_1960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5088__B1 (.DIODE(_1701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5089__A1 (.DIODE(\z80.tv80s.di_reg[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5089__A2 (.DIODE(_1701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5090__A1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__5090__B2 (.DIODE(_1696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5092__A0 (.DIODE(\z80.tv80s.i_tv80_core.I[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5094__A1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__5095__A (.DIODE(\z80.tv80s.di_reg[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5095__B (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__5096__A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__5097__A0 (.DIODE(\z80.tv80s.i_tv80_core.I[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5097__S (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__5099__S0 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__5099__S1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__5100__S0 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__5100__S1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__5101__S (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__5102__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__5103__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5103__A2 (.DIODE(_1691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5105__S (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__5108__A0 (.DIODE(\z80.tv80s.di_reg[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5108__S (.DIODE(_1701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5109__A1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__5109__B2 (.DIODE(_1696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5111__A0 (.DIODE(\z80.tv80s.i_tv80_core.I[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5114__A0 (.DIODE(\z80.tv80s.di_reg[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5114__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__5115__A0 (.DIODE(\z80.tv80s.i_tv80_core.I[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5115__S (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__5117__C_N (.DIODE(_0781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5119__A (.DIODE(_0856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5119__B (.DIODE(_1996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5122__A (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__5122__B (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__5124__A (.DIODE(_2846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5124__B (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__5126__A1 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__5126__A2 (.DIODE(\z80.tv80s.i_tv80_core.F[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5127__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5129__A (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__5129__B (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__5130__A (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__5130__B (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__5133__A1_N (.DIODE(\z80.tv80s.i_tv80_core.F[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5133__B2 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__5135__A1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__5139__A2 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__5139__B1 (.DIODE(\z80.tv80s.i_tv80_core.F[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5140__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__5140__A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__5143__A1 (.DIODE(_1996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5144__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__5145__C (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__5146__D (.DIODE(_0653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5147__A (.DIODE(_1996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5147__B (.DIODE(_2022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5148__A2 (.DIODE(\z80.tv80s.i_tv80_core.F[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5149__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5151__A (.DIODE(_1626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5152__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5152__B2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__5154__A1_N (.DIODE(_1014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5154__A2_N (.DIODE(_1996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5155__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__5156__A0 (.DIODE(\z80.tv80s.i_tv80_core.F[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5157__S (.DIODE(_1626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5158__A (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__5169__A0 (.DIODE(\z80.tv80s.i_tv80_core.F[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5170__A (.DIODE(\z80.tv80s.i_tv80_core.BusA[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5178__A (.DIODE(\z80.tv80s.i_tv80_core.F[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5179__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5188__B1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__5189__A1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__5189__A2 (.DIODE(\z80.tv80s.i_tv80_core.F[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5193__B (.DIODE(\z80.tv80s.i_tv80_core.BusA[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5196__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusB[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5196__B2 (.DIODE(\z80.tv80s.i_tv80_core.BusB[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5197__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusB[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5197__B2 (.DIODE(\z80.tv80s.i_tv80_core.BusB[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5198__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusB[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5198__A2 (.DIODE(_0405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5198__B2 (.DIODE(\z80.tv80s.i_tv80_core.BusB[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5200__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusB[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5204__B2 (.DIODE(\z80.tv80s.i_tv80_core.F[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5207__A (.DIODE(\z80.tv80s.di_reg[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5207__B (.DIODE(\z80.tv80s.di_reg[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5208__A (.DIODE(\z80.tv80s.di_reg[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5208__B (.DIODE(\z80.tv80s.di_reg[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5210__A (.DIODE(\z80.tv80s.di_reg[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5210__B (.DIODE(\z80.tv80s.di_reg[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5211__A (.DIODE(\z80.tv80s.di_reg[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5211__B (.DIODE(\z80.tv80s.di_reg[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5212__A (.DIODE(\z80.tv80s.di_reg[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5212__B (.DIODE(\z80.tv80s.di_reg[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5216__B1 (.DIODE(_2022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5217__A1_N (.DIODE(_2022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5219__S (.DIODE(_1996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5220__S (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__5222__A0 (.DIODE(\z80.tv80s.i_tv80_core.F[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5223__A0 (.DIODE(\z80.tv80s.i_tv80_core.ACC[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5225__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5225__B2 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__5226__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusB[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5227__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusB[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5227__A2 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__5228__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5231__S (.DIODE(_1996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5232__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__5236__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5237__A1 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__5237__B1 (.DIODE(\z80.tv80s.i_tv80_core.F[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5239__A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__5241__A1_N (.DIODE(_1150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5241__A2_N (.DIODE(_1996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5242__S (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__5243__A0 (.DIODE(\z80.tv80s.i_tv80_core.F[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5244__A0 (.DIODE(\z80.tv80s.i_tv80_core.ACC[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5245__A2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__5246__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5246__B2 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__5247__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusB[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5248__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusB[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5248__A2 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__5249__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5252__A0 (.DIODE(_1191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5252__S (.DIODE(_1996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5254__S (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__5261__A (.DIODE(\z80.tv80s.i_tv80_core.BusA[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5265__A1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__5265__A2 (.DIODE(\z80.tv80s.i_tv80_core.F[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5266__A1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__5268__A (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__5268__C (.DIODE(\z80.tv80s.i_tv80_core.BusA[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5268__D (.DIODE(\z80.tv80s.i_tv80_core.BusA[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5272__A2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__5273__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5275__A (.DIODE(\z80.tv80s.i_tv80_core.I[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5275__C (.DIODE(\z80.tv80s.i_tv80_core.I[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5276__A1 (.DIODE(\z80.tv80s.i_tv80_core.I[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5278__A (.DIODE(\z80.tv80s.di_reg[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5278__B (.DIODE(\z80.tv80s.di_reg[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5278__C (.DIODE(\z80.tv80s.di_reg[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5278__D (.DIODE(\z80.tv80s.di_reg[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5279__A (.DIODE(\z80.tv80s.di_reg[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5279__B (.DIODE(\z80.tv80s.di_reg[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5280__S (.DIODE(_2022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5281__A0 (.DIODE(_1245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5281__S (.DIODE(_1996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5283__S (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__5284__A0 (.DIODE(\z80.tv80s.i_tv80_core.F[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5285__A0 (.DIODE(\z80.tv80s.i_tv80_core.F[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5285__S (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__5287__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5288__A0 (.DIODE(\z80.tv80s.i_tv80_core.F[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5289__A1 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA__5289__S (.DIODE(_1626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5291__A0 (.DIODE(\z80.tv80s.di_reg[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5291__S (.DIODE(_2022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5292__A0 (.DIODE(_1295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5292__S (.DIODE(_1996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5293__S (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__5297__A2 (.DIODE(_2166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5297__B1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__5298__A2 (.DIODE(_2166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5299__C (.DIODE(_2166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5305__B2 (.DIODE(_2174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5306__A1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__5308__A1 (.DIODE(_2929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5308__A2 (.DIODE(_0477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5312__A1 (.DIODE(_0397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5314__A0 (.DIODE(_0537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5314__A1 (.DIODE(_2849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5314__S (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__5315__A (.DIODE(_2847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5316__A (.DIODE(_2999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5317__B (.DIODE(_0398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5318__B1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__5319__B1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__5320__A1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__5321__A1_N (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__5322__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__5324__A1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__5325__A1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__5328__B2 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__5331__B2 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA__5332__A_N (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__5332__C (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5333__A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__5334__A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__5335__A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__5337__A1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__5337__C1 (.DIODE(_3021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5338__A1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__5338__A3 (.DIODE(_0397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5339__B2 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__5340__A1 (.DIODE(\z80.tv80s.i_tv80_core.IR[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5340__A2 (.DIODE(_0398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5341__A (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__5342__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__5343__A1 (.DIODE(_2999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5344__B (.DIODE(_2950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5347__A1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__5348__A3 (.DIODE(_2960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5349__A2 (.DIODE(_2995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5353__A1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__5353__B2 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA__5354__A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__5354__A2 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__5356__A1 (.DIODE(_2982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5356__A2 (.DIODE(_0537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5357__A1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__5358__B2 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__5359__B1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__5360__C (.DIODE(_0537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5361__B1 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA__5362__A (.DIODE(_0684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5364__A (.DIODE(_2999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5365__A1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__5369__B (.DIODE(_2929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5374__C (.DIODE(_0474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5375__A1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__5377__A1 (.DIODE(_2999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5377__A2 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__5378__A1 (.DIODE(_1525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5378__B1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__5379__S (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__5380__A1 (.DIODE(_1333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5380__B1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__5381__S (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__5382__A1 (.DIODE(_1349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5382__B1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__5384__A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__5385__A1 (.DIODE(_0577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5387__C (.DIODE(_0397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5388__A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__5390__B1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__5392__A2 (.DIODE(_0577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5393__B2 (.DIODE(_0684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5394__A2 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__5394__A3 (.DIODE(_1412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5394__B1 (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5395__A0 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__5395__S (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__5396__A1 (.DIODE(_1412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5397__A1 (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5398__A (.DIODE(_2934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5401__A1 (.DIODE(_2847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5402__A1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__5404__A0 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__5406__A (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__5409__A1 (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5409__B2 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__5411__A (.DIODE(_2854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5412__A1 (.DIODE(_2854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5412__B1 (.DIODE(_1673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5413__A (.DIODE(\z80.tv80s.di_reg[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5413__B (.DIODE(_1673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5414__A1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__5415__A (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5415__B (.DIODE(\z80.tv80s.i_tv80_core.ts[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5416__A (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5416__B (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__5417__B (.DIODE(_2266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5418__A (.DIODE(_0603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5419__A1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__5420__B2 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__5421__A0 (.DIODE(\z80.tv80s.di_reg[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5422__A (.DIODE(_0604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5423__A (.DIODE(_2266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5424__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__5424__A3 (.DIODE(_2273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5424__B1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__5425__A1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__5426__A1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__5426__C1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__5427__A (.DIODE(\z80.tv80s.i_tv80_core.ts[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5427__B (.DIODE(_2871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5428__S (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__5429__A (.DIODE(_2275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5430__A1 (.DIODE(_2275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5434__A2 (.DIODE(_2273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5434__B2 (.DIODE(_2265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5435__A1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__5436__S (.DIODE(_0598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5437__A0 (.DIODE(\z80.tv80s.di_reg[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5438__S (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__5439__A (.DIODE(_2854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5439__B (.DIODE(\z80.tv80s.di_reg[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5440__A1 (.DIODE(_1736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5440__S (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__5441__A (.DIODE(_2275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5442__A1 (.DIODE(_2275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5446__A2 (.DIODE(_2273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5446__B2 (.DIODE(_2265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5447__A1 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__5448__S (.DIODE(_0598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5449__A0 (.DIODE(\z80.tv80s.di_reg[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5450__S (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__5451__A (.DIODE(_2854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5451__B (.DIODE(\z80.tv80s.di_reg[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5452__A1 (.DIODE(_1754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5452__S (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__5453__A (.DIODE(_2275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5454__A1 (.DIODE(_2275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5458__A0 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__5458__A1 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5459__S (.DIODE(_2266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5460__A1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__5461__S (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__5462__A0 (.DIODE(\z80.tv80s.di_reg[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5464__A (.DIODE(_2854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5464__B (.DIODE(\z80.tv80s.di_reg[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5465__A1 (.DIODE(_1771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5465__S (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__5466__A (.DIODE(_2275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5467__A1 (.DIODE(_2275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5471__A0 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__5471__A1 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5472__S (.DIODE(_2266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5473__A1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__5474__S (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__5475__A0 (.DIODE(\z80.tv80s.di_reg[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5477__A (.DIODE(_2854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5477__B (.DIODE(\z80.tv80s.di_reg[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5478__A1 (.DIODE(_1789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5478__S (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__5479__A (.DIODE(_2275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5480__A1 (.DIODE(_2275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5484__A0 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__5484__A1 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5485__S (.DIODE(_2266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5486__A1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__5487__S (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__5488__A0 (.DIODE(\z80.tv80s.di_reg[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5489__S (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__5490__A (.DIODE(_2854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5490__B (.DIODE(\z80.tv80s.di_reg[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5491__A1 (.DIODE(_1807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5491__S (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__5492__A (.DIODE(_2275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5493__A1 (.DIODE(_2275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5497__A2 (.DIODE(_2273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5497__B2 (.DIODE(_2265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5498__A1 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__5499__S (.DIODE(_0598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5500__A0 (.DIODE(\z80.tv80s.di_reg[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5503__A1 (.DIODE(_2854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5503__A2 (.DIODE(\z80.tv80s.di_reg[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5503__B1 (.DIODE(_2275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5504__S (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__5509__A2_N (.DIODE(_2273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5509__B2 (.DIODE(_2266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5510__A1 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__5511__S (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__5512__A0 (.DIODE(\z80.tv80s.di_reg[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5515__A1 (.DIODE(_1847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5515__S (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__5520__B (.DIODE(_2273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5525__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__5525__B (.DIODE(_2366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5526__A2 (.DIODE(_2266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5527__A1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__5527__A3 (.DIODE(_2366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5527__B1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__5528__B1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__5529__A1 (.DIODE(_1866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5529__S (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__5536__A0 (.DIODE(\z80.tv80s.di_reg[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5537__S (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__5540__A1 (.DIODE(_1885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5540__S (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__5546__A2 (.DIODE(_2273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5546__B2 (.DIODE(_2265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5547__S (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__5548__A0 (.DIODE(\z80.tv80s.di_reg[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5549__S (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__5550__A1 (.DIODE(_1903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5550__S (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__5555__A2 (.DIODE(_2273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5555__B2 (.DIODE(_2265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5556__S (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__5557__A0 (.DIODE(\z80.tv80s.di_reg[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5558__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__5559__A1 (.DIODE(_1922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5559__S (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__5566__A2_N (.DIODE(_2273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5566__B2 (.DIODE(_2266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5567__B (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__5568__A1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__5569__A1 (.DIODE(\z80.tv80s.di_reg[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5570__S (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__5571__S (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__5578__A2 (.DIODE(_2273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5578__B2 (.DIODE(_2265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5579__S (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__5580__A0 (.DIODE(\z80.tv80s.di_reg[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5581__S (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__5582__A1 (.DIODE(_1960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5582__S (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__5588__A2 (.DIODE(_2273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5588__B2 (.DIODE(_2265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5589__S (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__5590__A0 (.DIODE(\z80.tv80s.di_reg[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5591__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__5593__S (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__5596__A2 (.DIODE(_2273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5596__B2 (.DIODE(_2265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5597__S (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__5598__A0 (.DIODE(\z80.tv80s.di_reg[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5599__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__5600__A (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__5602__A2 (.DIODE(_0401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5602__B1 (.DIODE(_0684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5602__B2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__5604__A1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__5605__A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__5605__B (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__5605__C (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__5606__A1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__5606__B2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__5607__B2 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__5609__A (.DIODE(_2441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5610__A (.DIODE(_1412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5610__B (.DIODE(_2441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5611__A1 (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5611__B1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__5612__A (.DIODE(_1412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5613__A1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__5613__A2 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__5614__A2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__5614__B1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__5615__A1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__5615__C1 (.DIODE(_2999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5617__B (.DIODE(_0481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5618__A2 (.DIODE(_0405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5620__A1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__5621__A1 (.DIODE(_2849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5621__A2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__5621__B1 (.DIODE(_0401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5623__B2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__5626__A1_N (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__5626__B2 (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5627__A (.DIODE(_2459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5628__A (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5629__A_N (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5629__C (.DIODE(_2459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5630__A (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5630__B (.DIODE(_1412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5631__A1 (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5631__A2 (.DIODE(_1412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5631__B1 (.DIODE(_2441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5633__A2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__5633__C1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__5634__A2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__5634__C1 (.DIODE(_0984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5635__A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__5635__C1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__5636__A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__5636__C1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__5637__A (.DIODE(_1300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5638__A1 (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5639__A (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5640__A2 (.DIODE(_1300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5641__A1 (.DIODE(_2459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5642__A (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5642__B (.DIODE(_2459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5644__A (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5644__B (.DIODE(_2459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5645__A (.DIODE(_1412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5646__A_N (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5646__C (.DIODE(_2459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5648__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5648__B2 (.DIODE(\z80.tv80s.i_tv80_core.ACC[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5650__A1 (.DIODE(\z80.tv80s.di_reg[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5651__A1 (.DIODE(\z80.tv80s.i_tv80_core.PC[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5652__A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__5654__A1 (.DIODE(\z80.tv80s.i_tv80_core.PC[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5654__B2 (.DIODE(\z80.tv80s.di_reg[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5655__B (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5656__A2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__5656__C1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__5657__A2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__5657__C1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__5658__A1 (.DIODE(_1300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5659__S (.DIODE(_2459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5660__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5662__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5664__A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__5665__A1 (.DIODE(\z80.tv80s.di_reg[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5666__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5666__B2 (.DIODE(\z80.tv80s.i_tv80_core.PC[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5667__A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__5667__C1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__5668__A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__5668__C1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__5669__A (.DIODE(_1300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5670__A2 (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5671__S (.DIODE(_2459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5672__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5675__A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__5677__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5677__B2 (.DIODE(\z80.tv80s.i_tv80_core.PC[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5678__A2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__5678__C1 (.DIODE(_0984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5679__A2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__5679__C1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__5681__A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__5681__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__5681__C1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__5682__A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__5682__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__5682__C1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__5684__S0 (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5684__S1 (.DIODE(_2459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5685__A1 (.DIODE(\z80.tv80s.di_reg[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5685__B1 (.DIODE(_2514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5686__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5688__A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__5690__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5690__B2 (.DIODE(\z80.tv80s.i_tv80_core.PC[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5691__A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__5691__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__5691__C1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__5692__A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__5692__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__5692__C1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__5694__A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__5694__C1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__5695__A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__5695__C1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__5697__S0 (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5697__S1 (.DIODE(_2459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5698__A1 (.DIODE(\z80.tv80s.di_reg[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5699__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5701__A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__5703__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5703__B2 (.DIODE(\z80.tv80s.i_tv80_core.PC[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5704__A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__5704__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__5704__C1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__5705__A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__5705__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__5705__C1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__5707__A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__5707__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__5707__C1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__5708__A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__5708__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__5708__C1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__5710__S0 (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5710__S1 (.DIODE(_2459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5711__A1 (.DIODE(\z80.tv80s.di_reg[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5711__B1 (.DIODE(_2538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5712__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5714__A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__5716__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5717__A2 (.DIODE(\z80.tv80s.i_tv80_core.RegAddrB_r[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5717__C1 (.DIODE(_0984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5718__A2 (.DIODE(\z80.tv80s.i_tv80_core.RegAddrB_r[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5720__A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__5720__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__5720__C1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__5721__A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__5721__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__5721__C1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__5723__S0 (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5723__S1 (.DIODE(_2459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5724__A1 (.DIODE(\z80.tv80s.di_reg[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5725__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5727__A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__5728__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5729__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5730__A2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__5730__C1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__5731__A2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__5731__C1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__5732__A (.DIODE(_1300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5733__A1 (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5734__S (.DIODE(_2459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5736__B2 (.DIODE(\z80.tv80s.di_reg[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5738__A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__5739__S (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__5741__S (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__5743__S (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__5744__S (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__5745__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__5746__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__5747__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__5748__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__5749__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__5750__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__5751__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__5752__A1 (.DIODE(_1107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5752__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__5753__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__5754__A1 (.DIODE(_1198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5754__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__5755__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__5756__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__5757__A (.DIODE(_2854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5757__B (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__5757__C (.DIODE(_0477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5758__A0 (.DIODE(\z80.tv80s.i_tv80_core.ACC[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5758__S (.DIODE(_2566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5759__A0 (.DIODE(\z80.tv80s.i_tv80_core.ACC[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5759__S (.DIODE(_2566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5760__A0 (.DIODE(\z80.tv80s.i_tv80_core.ACC[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5760__S (.DIODE(_2566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5761__A0 (.DIODE(\z80.tv80s.i_tv80_core.ACC[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5761__S (.DIODE(_2566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5762__A0 (.DIODE(\z80.tv80s.i_tv80_core.ACC[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5762__S (.DIODE(_2566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5763__A0 (.DIODE(\z80.tv80s.i_tv80_core.ACC[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5763__S (.DIODE(_2566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5764__A0 (.DIODE(\z80.tv80s.i_tv80_core.ACC[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5764__S (.DIODE(_2566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5765__A0 (.DIODE(\z80.tv80s.i_tv80_core.ACC[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5765__A1 (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA__5765__S (.DIODE(_2566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5766__A0 (.DIODE(\z80.tv80s.i_tv80_core.ACC[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5767__A (.DIODE(_1333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5768__S (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__5769__S (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__5770__A (.DIODE(\z80.tv80s.i_tv80_core.Halt_FF ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5771__A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__5771__B (.DIODE(_2568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5772__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__5772__B1 (.DIODE(_0605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5773__A2 (.DIODE(_2982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5775__A1 (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5776__B2 (.DIODE(_0397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5777__A (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__5777__B (.DIODE(_0554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5778__B1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__5779__A1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__5779__A2 (.DIODE(_0685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5780__A1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__5780__A2 (.DIODE(_2893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5780__B1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__5781__A3 (.DIODE(_0398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5781__C1 (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5782__A2 (.DIODE(_2577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5782__B1 (.DIODE(_0603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5783__A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__5784__A1 (.DIODE(_0577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5784__A2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__5784__B1 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__5785__A1 (.DIODE(_0577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5785__A2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__5785__B1 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__5788__C1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__5789__A2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__5790__A1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__5790__A3 (.DIODE(_0685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5790__B1 (.DIODE(_2577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5794__A1 (.DIODE(_2584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5794__B2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__5795__A1_N (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__5795__B1 (.DIODE(_2582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5798__C1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__5799__A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__5799__B (.DIODE(\z80.tv80s.di_reg[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5799__C (.DIODE(_0685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5800__B (.DIODE(_2577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5801__A1 (.DIODE(_2577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5806__A2 (.DIODE(_2584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5806__B2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__5807__A2 (.DIODE(_2583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5807__B2 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__5808__A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__5808__B (.DIODE(\z80.tv80s.di_reg[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5808__C (.DIODE(_0685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5809__B (.DIODE(_2577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5810__A1 (.DIODE(_2577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5816__S (.DIODE(_1681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5818__A2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__5819__A1 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__5819__B2 (.DIODE(_2584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5820__A1_N (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__5820__B1 (.DIODE(_2582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5821__A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__5821__B (.DIODE(\z80.tv80s.di_reg[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5821__C (.DIODE(_0685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5822__B (.DIODE(_2577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5823__A1 (.DIODE(_2577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5828__A0 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5829__A1 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5831__A1 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5831__A2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__5832__A1 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__5832__B2 (.DIODE(_2584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5833__A1_N (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__5833__B1 (.DIODE(_2582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5834__A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__5834__B (.DIODE(\z80.tv80s.di_reg[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5834__C (.DIODE(_0685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5835__B (.DIODE(_2577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5836__A1 (.DIODE(_2577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5841__A0 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5842__A1 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5844__A1 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5845__A1 (.DIODE(_2581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5845__B2 (.DIODE(_2584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5846__A1_N (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__5846__B1 (.DIODE(_2582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5848__A1 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5850__A0 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5850__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__5851__A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__5851__B (.DIODE(\z80.tv80s.di_reg[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5851__C (.DIODE(_0685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5852__B (.DIODE(_2577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5853__A1 (.DIODE(_2577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5858__A1 (.DIODE(_2584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5858__B2 (.DIODE(_2581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5859__A2 (.DIODE(_2583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5859__B2 (.DIODE(_2570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5860__A2 (.DIODE(_1685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5861__A1 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5863__A0 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5864__A1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__5864__B1_N (.DIODE(_2581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5865__A2 (.DIODE(_0577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5866__A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__5866__B (.DIODE(\z80.tv80s.di_reg[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5866__C (.DIODE(_0685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5867__B (.DIODE(_2577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5869__A1 (.DIODE(_2577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5873__A1 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__5874__S (.DIODE(_2570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5875__A0 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5876__A1 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5878__A0 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5878__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__5879__S (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__5880__A1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__5880__A2 (.DIODE(\z80.tv80s.di_reg[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5880__A3 (.DIODE(_0685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5880__B1 (.DIODE(_2577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5881__B (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__5882__B (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__5887__S (.DIODE(_2581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5888__S (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__5889__A (.DIODE(\z80.tv80s.i_tv80_core.PC[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5889__B (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__5892__A1 (.DIODE(\z80.tv80s.i_tv80_core.PC[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5895__B1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__5896__A1 (.DIODE(\z80.tv80s.di_reg[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5896__A2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__5896__C1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__5897__A2 (.DIODE(_0577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5897__B1_N (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__5898__A (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__5900__S (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__5902__A1 (.DIODE(\z80.tv80s.i_tv80_core.PC[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5902__A2 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__5904__A1 (.DIODE(\z80.tv80s.i_tv80_core.PC[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5907__A0 (.DIODE(\z80.tv80s.di_reg[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5907__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__5908__A1 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__5908__B2 (.DIODE(_2584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5909__A2 (.DIODE(_2583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5909__B2 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__5910__A (.DIODE(\z80.tv80s.i_tv80_core.PC[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5910__B (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__5911__A1 (.DIODE(\z80.tv80s.i_tv80_core.PC[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5911__A2 (.DIODE(\z80.tv80s.i_tv80_core.PC[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5916__A1 (.DIODE(\z80.tv80s.i_tv80_core.PC[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5919__B1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__5920__A2 (.DIODE(_2584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5920__B2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__5921__A1_N (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__5921__B1 (.DIODE(_2582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5922__B (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__5923__A1 (.DIODE(\z80.tv80s.i_tv80_core.PC[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5923__A2 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__5925__A1 (.DIODE(\z80.tv80s.i_tv80_core.PC[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5928__A0 (.DIODE(\z80.tv80s.di_reg[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5928__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__5929__S (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__5930__S (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__5931__S (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__5932__B (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__5933__B (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__5935__A1 (.DIODE(\z80.tv80s.i_tv80_core.PC[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5935__A2 (.DIODE(\z80.tv80s.i_tv80_core.PC[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5935__A3 (.DIODE(\z80.tv80s.i_tv80_core.PC[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5935__A4 (.DIODE(\z80.tv80s.i_tv80_core.PC[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5935__B1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__5938__A1 (.DIODE(\z80.tv80s.i_tv80_core.PC[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5941__A0 (.DIODE(\z80.tv80s.di_reg[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5941__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__5942__S (.DIODE(_0576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5943__S (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__5944__S (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__5945__A0 (.DIODE(\z80.tv80s.i_tv80_core.I[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5945__A1 (.DIODE(\z80.tv80s.i_tv80_core.PC[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5948__A0 (.DIODE(\z80.tv80s.di_reg[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5948__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__5949__B (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__5950__A (.DIODE(\z80.tv80s.i_tv80_core.PC[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5950__B (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__5951__B (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__5955__A1 (.DIODE(_2584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5955__B2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__5956__A2 (.DIODE(_2583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5956__B2 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__5957__B (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__5958__B (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__5962__A0 (.DIODE(\z80.tv80s.i_tv80_core.I[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5965__B1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__5966__A2 (.DIODE(_2584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5966__B2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__5967__A1_N (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__5967__B1 (.DIODE(_2582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5970__A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__5971__A0 (.DIODE(\z80.tv80s.i_tv80_core.I[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5974__A0 (.DIODE(\z80.tv80s.di_reg[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5974__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__5975__S (.DIODE(_0576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5976__S (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__5977__S (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__5978__A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__5983__A1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__5986__A1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__5990__A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__5991__B1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__5993__A1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__5995__C (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__5997__B1 (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA__5998__A1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__5999__B2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__6000__A1 (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA__6001__A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__6001__B1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__6004__S (.DIODE(_2775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6005__S (.DIODE(_2775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6006__S (.DIODE(_2775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6007__S (.DIODE(_2775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6008__S (.DIODE(_2775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6009__S (.DIODE(_2775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6010__S (.DIODE(_2775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6011__S (.DIODE(_2775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6012__A0 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__6012__S (.DIODE(_0604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6013__A0 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__6013__S (.DIODE(_0604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6014__A0 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__6014__S (.DIODE(_0604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6015__A0 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__6015__S (.DIODE(_0604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6016__A0 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__6016__S (.DIODE(_0604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6017__A0 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__6017__S (.DIODE(_0604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6018__A0 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__6018__S (.DIODE(_0604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6019__A0 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__6019__A1 (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA__6019__S (.DIODE(_0604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6020__A1 (.DIODE(_2849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6021__S (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__6023__A (.DIODE(_0577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6028__A1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__6029__B2 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__6033__D_N (.DIODE(_0781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6034__B1 (.DIODE(_0603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6037__A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__6038__A1 (.DIODE(_1416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6038__A2 (.DIODE(_2785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6040__B1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__6041__A1 (.DIODE(_1416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6041__A2 (.DIODE(_1673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6041__B2 (.DIODE(_2785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6042__A1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__6043__A (.DIODE(_0856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6044__A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__6045__A1 (.DIODE(_1416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6045__B2 (.DIODE(_2785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6046__A1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__6047__A (.DIODE(_1014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6048__A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__6049__A1 (.DIODE(_1416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6049__A2 (.DIODE(_1736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6049__B2 (.DIODE(_2785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6050__A1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__6051__A (.DIODE(_1066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6052__A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__6053__A1 (.DIODE(_1416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6053__A2 (.DIODE(_1754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6053__B2 (.DIODE(_2785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6055__A (.DIODE(_1100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6056__A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__6057__A1 (.DIODE(_1416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6057__A2 (.DIODE(_1771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6057__B2 (.DIODE(_2785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6059__A (.DIODE(_1150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6060__A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__6061__A1 (.DIODE(_1416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6061__A2 (.DIODE(_1789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6061__B2 (.DIODE(_2785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6063__A (.DIODE(_1191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6064__A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__6065__A1 (.DIODE(_1416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6065__A2 (.DIODE(_1807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6065__B2 (.DIODE(_2785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6067__A (.DIODE(_1245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6068__A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__6069__A1 (.DIODE(_1415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6069__A2 (.DIODE(_1827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6070__A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__6071__A0 (.DIODE(_1295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6072__B2 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__6074__B1 (.DIODE(_1416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6074__B2 (.DIODE(_1847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6075__B1 (.DIODE(_2814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6076__A (.DIODE(_0856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6076__B (.DIODE(_2814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6077__A2 (.DIODE(_2814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6077__B1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__6078__A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__6079__A1 (.DIODE(_1416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6079__A2 (.DIODE(_1866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6079__B2 (.DIODE(_2785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6080__B1 (.DIODE(_2814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6081__A (.DIODE(_1014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6081__B (.DIODE(_2814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6082__A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__6083__A1 (.DIODE(_1416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6083__A2 (.DIODE(_1885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6083__B2 (.DIODE(_2785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6084__B1 (.DIODE(_2814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6085__A (.DIODE(_1066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6085__B (.DIODE(_2814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6086__A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__6087__A1 (.DIODE(_1416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6087__A2 (.DIODE(_1903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6087__B2 (.DIODE(_2785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6088__B1 (.DIODE(_2814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6089__A (.DIODE(_1100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6089__B (.DIODE(_2814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6090__A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__6091__B1 (.DIODE(_1416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6091__B2 (.DIODE(_1922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6092__B1 (.DIODE(_2814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6093__A (.DIODE(_1150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6093__B (.DIODE(_2814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6094__A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__6095__A1 (.DIODE(_1416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6095__B2 (.DIODE(_2785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6096__B1 (.DIODE(_2814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6097__A (.DIODE(_1191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6097__B (.DIODE(_2814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6098__A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__6100__A (.DIODE(_1415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6101__B (.DIODE(_1416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6101__C (.DIODE(_1960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6102__A2 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__6102__B1 (.DIODE(_2814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6103__A1_N (.DIODE(_1245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6103__A2_N (.DIODE(_2814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6104__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__6105__A1 (.DIODE(_1416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6105__B2 (.DIODE(_2785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6107__A0 (.DIODE(_1295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6107__S (.DIODE(_2814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6108__S (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__6130__RESET_B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__6131__RESET_B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__6133__RESET_B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__6150__RESET_B (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__6163__D (.DIODE(_0020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6242__RESET_B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__6245__RESET_B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__6246__RESET_B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__6247__RESET_B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__6248__RESET_B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__6257__RESET_B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__6258__RESET_B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__6275__SET_B (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__6276__SET_B (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__6279__SET_B (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__6292__RESET_B (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__6301__RESET_B (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__6302__RESET_B (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__6303__RESET_B (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__6304__RESET_B (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__6305__RESET_B (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__6306__RESET_B (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__6307__RESET_B (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__6308__RESET_B (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__6333__SET_B (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__6334__SET_B (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__6336__SET_B (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__6337__SET_B (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__6338__SET_B (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__6339__SET_B (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__6340__SET_B (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__6348__RESET_B (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__6349__RESET_B (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__6350__RESET_B (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__6361__RESET_B (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__6362__RESET_B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__6363__RESET_B (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__6364__RESET_B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__6365__RESET_B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__6366__RESET_B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__6367__RESET_B (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__6368__RESET_B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__6369__RESET_B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6370__RESET_B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6371__RESET_B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6372__RESET_B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6373__RESET_B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6374__RESET_B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6375__RESET_B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6376__RESET_B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6377__RESET_B (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__6427__RESET_B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6428__RESET_B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6441__RESET_B (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__6442__RESET_B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__6446__RESET_B (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__6448__CLK (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__6448__RESET_B (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__6458__RESET_B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__6459__RESET_B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__6460__RESET_B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__6461__RESET_B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__6462__RESET_B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__6463__RESET_B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__6464__RESET_B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__6465__RESET_B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__6474__RESET_B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__6475__SET_B (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__6476__SET_B (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__6477__SET_B (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__6478__SET_B (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__6479__SET_B (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__6480__SET_B (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__6481__SET_B (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__6482__SET_B (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__6483__SET_B (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__6484__SET_B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6485__SET_B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6486__SET_B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6487__SET_B (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__6488__SET_B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6489__SET_B (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__6490__SET_B (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__6523__A (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__6524__A (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__6525__A (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__6526__A (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__6527__A (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__6528__A (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__6529__A (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_14_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_15_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_18_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_19_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_20_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_21_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_22_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_23_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_24_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_25_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_26_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_27_wb_clk_i_A (.DIODE(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_28_wb_clk_i_A (.DIODE(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_29_wb_clk_i_A (.DIODE(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_30_wb_clk_i_A (.DIODE(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_31_wb_clk_i_A (.DIODE(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_32_wb_clk_i_A (.DIODE(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_33_wb_clk_i_A (.DIODE(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_34_wb_clk_i_A (.DIODE(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_35_wb_clk_i_A (.DIODE(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_36_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_37_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_38_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_39_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_40_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_41_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_42_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_43_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_44_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_45_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_46_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_47_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_48_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_49_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_50_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout100_A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout101_A (.DIODE(_0598_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout102_A (.DIODE(_0598_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout103_A (.DIODE(_0501_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout104_A (.DIODE(_0501_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout112_A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout113_A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout114_A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout115_A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout116_A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout117_A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout118_A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout121_A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout123_A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout124_A (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout125_A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout126_A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout127_A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout128_A (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout131_A (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout132_A (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout133_A (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout134_A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout135_A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout136_A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout138_A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout141_A (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout144_A (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout145_A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout148_A (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout149_A (.DIODE(\z80.tv80s.i_tv80_core.IR[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout150_A (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout151_A (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout153_A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout155_A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout156_A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout158_A (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout160_A (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout163_A (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout164_A (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout165_A (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout166_A (.DIODE(\z80.tv80s.i_tv80_core.ISet[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout167_A (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout171_A (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout172_A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout173_A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout174_A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout175_A (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout176_A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout177_A (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout178_A (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout179_A (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout180_A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout181_A (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout182_A (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout183_A (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout184_A (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout185_A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout60_A (.DIODE(_0576_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout63_A (.DIODE(_2570_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout64_A (.DIODE(_2581_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout68_A (.DIODE(_1681_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout73_A (.DIODE(_0984_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout74_A (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout82_A (.DIODE(_0981_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout83_A (.DIODE(_0981_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout84_A (.DIODE(_0981_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout88_A (.DIODE(_1418_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout89_A (.DIODE(_0772_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout90_A (.DIODE(_1417_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout93_A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout94_A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout96_A (.DIODE(_2995_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout99_A (.DIODE(_1685_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1_A (.DIODE(\z80.tv80s.i_tv80_core.BusReq_s ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold387_A (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold389_A (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold399_A (.DIODE(\z80.tv80s.i_tv80_core.BusB[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold409_A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold411_A (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold419_A (.DIODE(\z80.tv80s.i_tv80_core.BusB[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold423_A (.DIODE(\z80.tv80s.i_tv80_core.BusB[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold425_A (.DIODE(\z80.tv80s.i_tv80_core.BusB[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold427_A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold429_A (.DIODE(\z80.tv80s.i_tv80_core.BusB[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold431_A (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold452_A (.DIODE(\z80.tv80s.i_tv80_core.BusA[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold470_A (.DIODE(\z80.tv80s.i_tv80_core.BusA[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold489_A (.DIODE(\z80.tv80s.i_tv80_core.BusB[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold491_A (.DIODE(\z80.tv80s.i_tv80_core.Halt_FF ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold502_A (.DIODE(\z80.tv80s.i_tv80_core.I[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold504_A (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold506_A (.DIODE(\z80.tv80s.i_tv80_core.BusA[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold508_A (.DIODE(\z80.tv80s.i_tv80_core.BusB[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold512_A (.DIODE(\z80.tv80s.i_tv80_core.I[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold516_A (.DIODE(\z80.tv80s.i_tv80_core.ts[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold529_A (.DIODE(\z80.tv80s.i_tv80_core.BusA[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold548_A (.DIODE(\z80.tv80s.i_tv80_core.BusA[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold552_A (.DIODE(\z80.tv80s.i_tv80_core.PC[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold554_A (.DIODE(\z80.tv80s.i_tv80_core.BusB[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold558_A (.DIODE(\z80.tv80s.i_tv80_core.IntCycle ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold560_A (.DIODE(\z80.tv80s.i_tv80_core.PC[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold564_A (.DIODE(\z80.tv80s.i_tv80_core.BusA[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold566_A (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold568_A (.DIODE(\z80.tv80s.i_tv80_core.PC[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold572_A (.DIODE(\z80.tv80s.i_tv80_core.I[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold579_A (.DIODE(\z80.tv80s.i_tv80_core.PC[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold586_A (.DIODE(\z80.tv80s.i_tv80_core.PC[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold588_A (.DIODE(\z80.tv80s.i_tv80_core.PC[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold590_A (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold592_A (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold595_A (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold598_A (.DIODE(\z80.tv80s.i_tv80_core.F[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold601_A (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold603_A (.DIODE(\z80.tv80s.i_tv80_core.F[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold607_A (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold610_A (.DIODE(\z80.tv80s.i_tv80_core.F[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold613_A (.DIODE(\z80.tv80s.i_tv80_core.F[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold616_A (.DIODE(\z80.tv80s.di_reg[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold618_A (.DIODE(\z80.tv80s.di_reg[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold620_A (.DIODE(\z80.tv80s.di_reg[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold621_A (.DIODE(\z80.tv80s.di_reg[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold624_A (.DIODE(\z80.tv80s.di_reg[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold626_A (.DIODE(\z80.tv80s.di_reg[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold627_A (.DIODE(\z80.tv80s.di_reg[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold628_A (.DIODE(\z80.tv80s.di_reg[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold629_A (.DIODE(\z80.tv80s.i_tv80_core.ACC[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold630_A (.DIODE(\z80.tv80s.i_tv80_core.ACC[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold631_A (.DIODE(\z80.tv80s.i_tv80_core.ACC[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold632_A (.DIODE(\z80.tv80s.i_tv80_core.ACC[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold634_A (.DIODE(\z80.tv80s.i_tv80_core.F[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold635_A (.DIODE(\z80.tv80s.i_tv80_core.ACC[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold636_A (.DIODE(\z80.tv80s.i_tv80_core.F[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold637_A (.DIODE(\z80.tv80s.i_tv80_core.ACC[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold639_A (.DIODE(\z80.tv80s.i_tv80_core.ACC[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold641_A (.DIODE(\z80.tv80s.i_tv80_core.RegAddrC[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold642_A (.DIODE(\z80.tv80s.i_tv80_core.ACC[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold643_A (.DIODE(\z80.tv80s.i_tv80_core.F[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold645_A (.DIODE(\z80.tv80s.i_tv80_core.F[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold648_A (.DIODE(\z80.tv80s.i_tv80_core.IR[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold652_A (.DIODE(\z80.tv80s.i_tv80_core.RegAddrB_r[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap91_A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_output26_A (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_output27_A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_output34_A (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_output36_A (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_output37_A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_output38_A (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_output39_A (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_output40_A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_output49_A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_output51_A (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_output52_A (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_output54_A (.DIODE(net54));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_562 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_560 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_588 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_282 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_543 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_562 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_30 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_8 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_538 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_394 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_476 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_170 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_499 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_366 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_592 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_583 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_594 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_594 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_171 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_594 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_560 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_507 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_90 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__inv_2 _3054_ (.A(net129),
    .Y(_2842_));
 sky130_fd_sc_hd__inv_2 _3055_ (.A(net160),
    .Y(_2843_));
 sky130_fd_sc_hd__inv_2 _3056_ (.A(net155),
    .Y(_2844_));
 sky130_fd_sc_hd__inv_2 _3057_ (.A(net153),
    .Y(_2845_));
 sky130_fd_sc_hd__inv_2 _3058_ (.A(net148),
    .Y(_2846_));
 sky130_fd_sc_hd__inv_6 _3059_ (.A(net146),
    .Y(_2847_));
 sky130_fd_sc_hd__inv_4 _3060_ (.A(net131),
    .Y(_2848_));
 sky130_fd_sc_hd__inv_6 _3061_ (.A(net136),
    .Y(_2849_));
 sky130_fd_sc_hd__inv_2 _3062_ (.A(\z80.tv80s.i_tv80_core.ISet[0] ),
    .Y(_2850_));
 sky130_fd_sc_hd__inv_2 _3063_ (.A(net163),
    .Y(_2851_));
 sky130_fd_sc_hd__inv_2 _3064_ (.A(net854),
    .Y(_2852_));
 sky130_fd_sc_hd__inv_2 _3065_ (.A(\z80.tv80s.i_tv80_core.i_mcode.MCycle[3] ),
    .Y(_2853_));
 sky130_fd_sc_hd__inv_4 _3066_ (.A(net121),
    .Y(_2854_));
 sky130_fd_sc_hd__inv_2 _3067_ (.A(\z80.tv80s.i_tv80_core.ts[1] ),
    .Y(_2855_));
 sky130_fd_sc_hd__inv_4 _3068_ (.A(net829),
    .Y(_2856_));
 sky130_fd_sc_hd__inv_2 _3069_ (.A(net523),
    .Y(_2857_));
 sky130_fd_sc_hd__inv_2 _3070_ (.A(net123),
    .Y(net27));
 sky130_fd_sc_hd__inv_2 _3071_ (.A(net221),
    .Y(_2858_));
 sky130_fd_sc_hd__inv_2 _3072_ (.A(net140),
    .Y(_2859_));
 sky130_fd_sc_hd__inv_2 _3073_ (.A(net605),
    .Y(_2860_));
 sky130_fd_sc_hd__inv_2 _3074_ (.A(\z80.tv80s.i_tv80_core.Halt_FF ),
    .Y(net50));
 sky130_fd_sc_hd__inv_2 _3075_ (.A(\z80.tv80s.i_tv80_core.Save_ALU_r ),
    .Y(_2861_));
 sky130_fd_sc_hd__inv_2 _3076_ (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ),
    .Y(_2862_));
 sky130_fd_sc_hd__inv_2 _3077_ (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[0] ),
    .Y(_2863_));
 sky130_fd_sc_hd__inv_2 _3078_ (.A(net143),
    .Y(_2864_));
 sky130_fd_sc_hd__inv_2 _3079_ (.A(\z80.tv80s.i_tv80_core.BusA[1] ),
    .Y(_2865_));
 sky130_fd_sc_hd__inv_2 _3080_ (.A(\z80.tv80s.i_tv80_core.BusA[2] ),
    .Y(_2866_));
 sky130_fd_sc_hd__inv_2 _3081_ (.A(net645),
    .Y(_2867_));
 sky130_fd_sc_hd__inv_2 _3082_ (.A(\z80.tv80s.i_tv80_core.BusB[2] ),
    .Y(_2868_));
 sky130_fd_sc_hd__inv_2 _3083_ (.A(net619),
    .Y(_2869_));
 sky130_fd_sc_hd__inv_2 _3084_ (.A(\z80.tv80s.i_tv80_core.Arith16_r ),
    .Y(_2870_));
 sky130_fd_sc_hd__inv_2 _3085_ (.A(\z80.tv80s.di_reg[1] ),
    .Y(_2871_));
 sky130_fd_sc_hd__inv_2 _3086_ (.A(\z80.tv80s.di_reg[0] ),
    .Y(_2872_));
 sky130_fd_sc_hd__inv_2 _3087_ (.A(\z80.tv80s.i_tv80_core.Read_To_Reg_r[0] ),
    .Y(_2873_));
 sky130_fd_sc_hd__inv_2 _3088_ (.A(net464),
    .Y(_2874_));
 sky130_fd_sc_hd__inv_2 _3089_ (.A(net720),
    .Y(_2875_));
 sky130_fd_sc_hd__inv_2 _3090_ (.A(\z80.tv80s.i_tv80_core.ACC[0] ),
    .Y(_2876_));
 sky130_fd_sc_hd__inv_2 _3091_ (.A(net544),
    .Y(_2877_));
 sky130_fd_sc_hd__inv_2 _3092_ (.A(\z80.tv80s.i_tv80_core.ACC[3] ),
    .Y(_2878_));
 sky130_fd_sc_hd__inv_2 _3093_ (.A(\z80.tv80s.i_tv80_core.ACC[5] ),
    .Y(_2879_));
 sky130_fd_sc_hd__inv_2 _3094_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[2] ),
    .Y(_2880_));
 sky130_fd_sc_hd__inv_2 _3095_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[8] ),
    .Y(_2881_));
 sky130_fd_sc_hd__inv_2 _3096_ (.A(net563),
    .Y(_2882_));
 sky130_fd_sc_hd__inv_2 _3097_ (.A(net562),
    .Y(_2883_));
 sky130_fd_sc_hd__inv_2 _3098_ (.A(net5),
    .Y(_2884_));
 sky130_fd_sc_hd__inv_2 _3099_ (.A(net15),
    .Y(_0025_));
 sky130_fd_sc_hd__inv_2 _3100_ (.A(net16),
    .Y(_0023_));
 sky130_fd_sc_hd__inv_2 _3101__1 (.A(clknet_leaf_9_wb_clk_i),
    .Y(net218));
 sky130_fd_sc_hd__nor2_1 _3102_ (.A(\z80.tv80s.i_tv80_core.IR[7] ),
    .B(\z80.tv80s.i_tv80_core.IR[6] ),
    .Y(_2885_));
 sky130_fd_sc_hd__or2_1 _3103_ (.A(\z80.tv80s.i_tv80_core.IR[7] ),
    .B(\z80.tv80s.i_tv80_core.IR[6] ),
    .X(_2886_));
 sky130_fd_sc_hd__or3b_2 _3104_ (.A(\z80.tv80s.i_tv80_core.IR[7] ),
    .B(\z80.tv80s.i_tv80_core.IR[6] ),
    .C_N(net145),
    .X(_2887_));
 sky130_fd_sc_hd__or2_2 _3105_ (.A(_2846_),
    .B(_2887_),
    .X(_2888_));
 sky130_fd_sc_hd__inv_2 _3106_ (.A(_2888_),
    .Y(_2889_));
 sky130_fd_sc_hd__and2b_2 _3107_ (.A_N(net160),
    .B(net158),
    .X(_2890_));
 sky130_fd_sc_hd__nand2_2 _3108_ (.A(net158),
    .B(_2843_),
    .Y(_2891_));
 sky130_fd_sc_hd__and3_2 _3109_ (.A(net156),
    .B(net120),
    .C(_2890_),
    .X(_2892_));
 sky130_fd_sc_hd__and2_4 _3110_ (.A(_2889_),
    .B(_2892_),
    .X(_2893_));
 sky130_fd_sc_hd__o31a_2 _3111_ (.A1(net164),
    .A2(net567),
    .A3(net478),
    .B1(net651),
    .X(_2894_));
 sky130_fd_sc_hd__inv_2 _3112_ (.A(_2894_),
    .Y(_2895_));
 sky130_fd_sc_hd__and2_1 _3113_ (.A(\z80.tv80s.i_tv80_core.IR[7] ),
    .B(\z80.tv80s.i_tv80_core.IR[6] ),
    .X(_2896_));
 sky130_fd_sc_hd__nand2_8 _3114_ (.A(\z80.tv80s.i_tv80_core.IR[7] ),
    .B(\z80.tv80s.i_tv80_core.IR[6] ),
    .Y(_2897_));
 sky130_fd_sc_hd__nor2_1 _3115_ (.A(net148),
    .B(net144),
    .Y(_2898_));
 sky130_fd_sc_hd__or2_4 _3116_ (.A(net149),
    .B(net145),
    .X(_2899_));
 sky130_fd_sc_hd__nor2_1 _3117_ (.A(_2897_),
    .B(_2899_),
    .Y(_2900_));
 sky130_fd_sc_hd__or4bb_4 _3118_ (.A(net149),
    .B(net145),
    .C_N(\z80.tv80s.i_tv80_core.IR[7] ),
    .D_N(\z80.tv80s.i_tv80_core.IR[6] ),
    .X(_2901_));
 sky130_fd_sc_hd__and3_1 _3119_ (.A(net158),
    .B(net160),
    .C(_2844_),
    .X(_2902_));
 sky130_fd_sc_hd__nand3b_4 _3120_ (.A_N(net157),
    .B(net161),
    .C(net159),
    .Y(_2903_));
 sky130_fd_sc_hd__and3_2 _3121_ (.A(net150),
    .B(_2900_),
    .C(_2902_),
    .X(_2904_));
 sky130_fd_sc_hd__o21ai_1 _3122_ (.A1(_2893_),
    .A2(_2904_),
    .B1(\z80.tv80s.i_tv80_core.i_mcode.MCycle[5] ),
    .Y(_2905_));
 sky130_fd_sc_hd__nor2_1 _3123_ (.A(net158),
    .B(net160),
    .Y(_2906_));
 sky130_fd_sc_hd__or3_4 _3124_ (.A(net158),
    .B(net160),
    .C(net155),
    .X(_2907_));
 sky130_fd_sc_hd__or4_4 _3125_ (.A(net158),
    .B(net160),
    .C(net155),
    .D(net150),
    .X(_2908_));
 sky130_fd_sc_hd__nor3_4 _3126_ (.A(net110),
    .B(_2899_),
    .C(_2908_),
    .Y(_2909_));
 sky130_fd_sc_hd__or3_2 _3127_ (.A(net110),
    .B(_2899_),
    .C(_2908_),
    .X(_2910_));
 sky130_fd_sc_hd__or3_2 _3128_ (.A(_2846_),
    .B(net145),
    .C(_2897_),
    .X(_2911_));
 sky130_fd_sc_hd__nor2_4 _3129_ (.A(_2903_),
    .B(_2911_),
    .Y(_2912_));
 sky130_fd_sc_hd__or2_1 _3130_ (.A(_2903_),
    .B(_2911_),
    .X(_2913_));
 sky130_fd_sc_hd__nor2_1 _3131_ (.A(net150),
    .B(_2913_),
    .Y(_2914_));
 sky130_fd_sc_hd__nor2_1 _3132_ (.A(net152),
    .B(_2903_),
    .Y(_2915_));
 sky130_fd_sc_hd__or2_2 _3133_ (.A(net150),
    .B(_2903_),
    .X(_2916_));
 sky130_fd_sc_hd__nor2_1 _3134_ (.A(_2901_),
    .B(_2916_),
    .Y(_2917_));
 sky130_fd_sc_hd__or3_4 _3135_ (.A(net158),
    .B(_2843_),
    .C(net156),
    .X(_2918_));
 sky130_fd_sc_hd__or4bb_4 _3136_ (.A(net158),
    .B(net155),
    .C_N(net150),
    .D_N(net160),
    .X(_2919_));
 sky130_fd_sc_hd__inv_2 _3137_ (.A(_2919_),
    .Y(_2920_));
 sky130_fd_sc_hd__and3_1 _3138_ (.A(net149),
    .B(net145),
    .C(_2896_),
    .X(_2921_));
 sky130_fd_sc_hd__or3_2 _3139_ (.A(_2846_),
    .B(_2847_),
    .C(_2897_),
    .X(_2922_));
 sky130_fd_sc_hd__nor2_2 _3140_ (.A(_2919_),
    .B(_2922_),
    .Y(_2923_));
 sky130_fd_sc_hd__nor2_1 _3141_ (.A(_2904_),
    .B(_2923_),
    .Y(_2924_));
 sky130_fd_sc_hd__or2_1 _3142_ (.A(_2904_),
    .B(_2923_),
    .X(_2925_));
 sky130_fd_sc_hd__nor2_2 _3143_ (.A(_2903_),
    .B(_2922_),
    .Y(_2926_));
 sky130_fd_sc_hd__and3_2 _3144_ (.A(net159),
    .B(net161),
    .C(net157),
    .X(_2927_));
 sky130_fd_sc_hd__nand3_4 _3145_ (.A(net158),
    .B(net160),
    .C(net155),
    .Y(_2928_));
 sky130_fd_sc_hd__nor2_2 _3146_ (.A(_2887_),
    .B(_2928_),
    .Y(_2929_));
 sky130_fd_sc_hd__inv_2 _3147_ (.A(_2929_),
    .Y(_2930_));
 sky130_fd_sc_hd__or3_1 _3148_ (.A(_2925_),
    .B(_2926_),
    .C(_2929_),
    .X(_2931_));
 sky130_fd_sc_hd__or3_1 _3149_ (.A(_2909_),
    .B(_2912_),
    .C(_2917_),
    .X(_2932_));
 sky130_fd_sc_hd__and3_1 _3150_ (.A(_2847_),
    .B(_2885_),
    .C(_2927_),
    .X(_2933_));
 sky130_fd_sc_hd__nor2_4 _3151_ (.A(net147),
    .B(_2847_),
    .Y(_2934_));
 sky130_fd_sc_hd__nand2b_2 _3152_ (.A_N(net147),
    .B(net146),
    .Y(_2935_));
 sky130_fd_sc_hd__nor2_2 _3153_ (.A(_2897_),
    .B(_2935_),
    .Y(_2936_));
 sky130_fd_sc_hd__or2_1 _3154_ (.A(_2897_),
    .B(_2935_),
    .X(_2937_));
 sky130_fd_sc_hd__nor2_1 _3155_ (.A(_2919_),
    .B(_2937_),
    .Y(_2938_));
 sky130_fd_sc_hd__and4b_2 _3156_ (.A_N(net158),
    .B(net160),
    .C(net155),
    .D(net150),
    .X(_2939_));
 sky130_fd_sc_hd__and3_1 _3157_ (.A(net149),
    .B(_2896_),
    .C(_2939_),
    .X(_2940_));
 sky130_fd_sc_hd__a21o_1 _3158_ (.A1(_2936_),
    .A2(_2939_),
    .B1(_2940_),
    .X(_2941_));
 sky130_fd_sc_hd__or2_1 _3159_ (.A(_2938_),
    .B(_2941_),
    .X(_2942_));
 sky130_fd_sc_hd__or2_1 _3160_ (.A(_2933_),
    .B(_2942_),
    .X(_2943_));
 sky130_fd_sc_hd__nor2_1 _3161_ (.A(_2916_),
    .B(_2937_),
    .Y(_2944_));
 sky130_fd_sc_hd__nand2_4 _3162_ (.A(_2915_),
    .B(_2936_),
    .Y(_2945_));
 sky130_fd_sc_hd__nor2_1 _3163_ (.A(_2911_),
    .B(_2919_),
    .Y(_2946_));
 sky130_fd_sc_hd__or2_2 _3164_ (.A(_2944_),
    .B(_2946_),
    .X(_2947_));
 sky130_fd_sc_hd__nor2_4 _3165_ (.A(_2897_),
    .B(_2928_),
    .Y(_2948_));
 sky130_fd_sc_hd__nor2_2 _3166_ (.A(_2897_),
    .B(_2907_),
    .Y(_2949_));
 sky130_fd_sc_hd__and3_2 _3167_ (.A(net150),
    .B(_2902_),
    .C(_2936_),
    .X(_2950_));
 sky130_fd_sc_hd__or4b_4 _3168_ (.A(net159),
    .B(net160),
    .C(net156),
    .D_N(net151),
    .X(_2951_));
 sky130_fd_sc_hd__nor3_4 _3169_ (.A(net110),
    .B(_2899_),
    .C(_2951_),
    .Y(_2952_));
 sky130_fd_sc_hd__or2_1 _3170_ (.A(_2950_),
    .B(_2952_),
    .X(_2953_));
 sky130_fd_sc_hd__a211o_1 _3171_ (.A1(net145),
    .A2(_2949_),
    .B1(_2953_),
    .C1(_2948_),
    .X(_2954_));
 sky130_fd_sc_hd__nand2_1 _3172_ (.A(net161),
    .B(net151),
    .Y(_2955_));
 sky130_fd_sc_hd__mux2_1 _3173_ (.A0(net159),
    .A1(_2955_),
    .S(_2844_),
    .X(_2956_));
 sky130_fd_sc_hd__and2_1 _3174_ (.A(_2951_),
    .B(_2956_),
    .X(_2957_));
 sky130_fd_sc_hd__a21oi_1 _3175_ (.A1(_2916_),
    .A2(_2957_),
    .B1(_2888_),
    .Y(_2958_));
 sky130_fd_sc_hd__nor2_1 _3176_ (.A(net155),
    .B(_2891_),
    .Y(_2959_));
 sky130_fd_sc_hd__nand2_4 _3177_ (.A(_2844_),
    .B(_2890_),
    .Y(_2960_));
 sky130_fd_sc_hd__or2_2 _3178_ (.A(net149),
    .B(_2887_),
    .X(_2961_));
 sky130_fd_sc_hd__nor2_2 _3179_ (.A(_2960_),
    .B(_2961_),
    .Y(_2962_));
 sky130_fd_sc_hd__or2_1 _3180_ (.A(_2960_),
    .B(_2961_),
    .X(_2963_));
 sky130_fd_sc_hd__or4b_4 _3181_ (.A(net158),
    .B(net155),
    .C(net150),
    .D_N(net160),
    .X(_2964_));
 sky130_fd_sc_hd__nor2_4 _3182_ (.A(net110),
    .B(_2964_),
    .Y(_2965_));
 sky130_fd_sc_hd__or2_1 _3183_ (.A(_2886_),
    .B(_2964_),
    .X(_2966_));
 sky130_fd_sc_hd__nand2_1 _3184_ (.A(_2847_),
    .B(_2965_),
    .Y(_2967_));
 sky130_fd_sc_hd__nand2_1 _3185_ (.A(_2963_),
    .B(_2967_),
    .Y(_2968_));
 sky130_fd_sc_hd__or4_1 _3186_ (.A(_2947_),
    .B(_2954_),
    .C(_2958_),
    .D(_2968_),
    .X(_2969_));
 sky130_fd_sc_hd__or4_1 _3187_ (.A(_2931_),
    .B(_2932_),
    .C(_2943_),
    .D(_2969_),
    .X(_2970_));
 sky130_fd_sc_hd__and2b_2 _3188_ (.A_N(\z80.tv80s.i_tv80_core.IR[6] ),
    .B(\z80.tv80s.i_tv80_core.IR[7] ),
    .X(_2971_));
 sky130_fd_sc_hd__nand2b_2 _3189_ (.A_N(\z80.tv80s.i_tv80_core.IR[6] ),
    .B(\z80.tv80s.i_tv80_core.IR[7] ),
    .Y(_2972_));
 sky130_fd_sc_hd__a211o_1 _3190_ (.A1(_2908_),
    .A2(_2919_),
    .B1(_2972_),
    .C1(_2899_),
    .X(_2973_));
 sky130_fd_sc_hd__nor2_1 _3191_ (.A(net155),
    .B(net151),
    .Y(_2974_));
 sky130_fd_sc_hd__nand2_1 _3192_ (.A(_2890_),
    .B(_2974_),
    .Y(_2975_));
 sky130_fd_sc_hd__and2_1 _3193_ (.A(_2964_),
    .B(_2975_),
    .X(_2976_));
 sky130_fd_sc_hd__or4bb_2 _3194_ (.A(net158),
    .B(net150),
    .C_N(net155),
    .D_N(net160),
    .X(_2977_));
 sky130_fd_sc_hd__o21ai_1 _3195_ (.A1(net120),
    .A2(_2960_),
    .B1(_2977_),
    .Y(_2978_));
 sky130_fd_sc_hd__nand2_1 _3196_ (.A(_2936_),
    .B(_2978_),
    .Y(_2979_));
 sky130_fd_sc_hd__and2b_2 _3197_ (.A_N(\z80.tv80s.i_tv80_core.IR[7] ),
    .B(\z80.tv80s.i_tv80_core.IR[6] ),
    .X(_2980_));
 sky130_fd_sc_hd__nand2b_2 _3198_ (.A_N(\z80.tv80s.i_tv80_core.IR[7] ),
    .B(\z80.tv80s.i_tv80_core.IR[6] ),
    .Y(_2981_));
 sky130_fd_sc_hd__nor2_2 _3199_ (.A(_2844_),
    .B(_2891_),
    .Y(_2982_));
 sky130_fd_sc_hd__nand2_1 _3200_ (.A(net156),
    .B(_2890_),
    .Y(_2983_));
 sky130_fd_sc_hd__nor2_1 _3201_ (.A(net129),
    .B(net133),
    .Y(_2984_));
 sky130_fd_sc_hd__a311o_1 _3202_ (.A1(\z80.tv80s.i_tv80_core.i_mcode.MCycle[1] ),
    .A2(net108),
    .A3(_2982_),
    .B1(net135),
    .C1(\z80.tv80s.i_tv80_core.i_mcode.MCycle[6] ),
    .X(_2985_));
 sky130_fd_sc_hd__o2111a_1 _3203_ (.A1(_2901_),
    .A2(_2976_),
    .B1(_2979_),
    .C1(_2985_),
    .D1(_2973_),
    .X(_2986_));
 sky130_fd_sc_hd__or3_2 _3204_ (.A(net158),
    .B(_2844_),
    .C(net150),
    .X(_2987_));
 sky130_fd_sc_hd__and3_1 _3205_ (.A(net155),
    .B(net150),
    .C(_2906_),
    .X(_2988_));
 sky130_fd_sc_hd__a21oi_1 _3206_ (.A1(net151),
    .A2(_2959_),
    .B1(_2988_),
    .Y(_2989_));
 sky130_fd_sc_hd__a211o_1 _3207_ (.A1(_2987_),
    .A2(_2989_),
    .B1(net145),
    .C1(_2897_),
    .X(_2990_));
 sky130_fd_sc_hd__nor2_2 _3208_ (.A(_2960_),
    .B(net108),
    .Y(_2991_));
 sky130_fd_sc_hd__or2_2 _3209_ (.A(_2960_),
    .B(_2981_),
    .X(_2992_));
 sky130_fd_sc_hd__nor2_1 _3210_ (.A(net152),
    .B(_2992_),
    .Y(_2993_));
 sky130_fd_sc_hd__or4_4 _3211_ (.A(net158),
    .B(_2843_),
    .C(_2844_),
    .D(_2981_),
    .X(_2994_));
 sky130_fd_sc_hd__nor2_2 _3212_ (.A(_2846_),
    .B(_2847_),
    .Y(_2995_));
 sky130_fd_sc_hd__and4_1 _3213_ (.A(net120),
    .B(_2927_),
    .C(_2980_),
    .D(net96),
    .X(_2996_));
 sky130_fd_sc_hd__nor2_1 _3214_ (.A(net144),
    .B(_2981_),
    .Y(_2997_));
 sky130_fd_sc_hd__and3_2 _3215_ (.A(_2847_),
    .B(_2927_),
    .C(_2980_),
    .X(_2998_));
 sky130_fd_sc_hd__and3_4 _3216_ (.A(net155),
    .B(_2906_),
    .C(net109),
    .X(_2999_));
 sky130_fd_sc_hd__nand2_1 _3217_ (.A(net109),
    .B(net97),
    .Y(_3000_));
 sky130_fd_sc_hd__and2b_2 _3218_ (.A_N(net145),
    .B(net149),
    .X(_3001_));
 sky130_fd_sc_hd__nand2_2 _3219_ (.A(_2971_),
    .B(_3001_),
    .Y(_3002_));
 sky130_fd_sc_hd__a21o_1 _3220_ (.A1(_2916_),
    .A2(_2987_),
    .B1(_3002_),
    .X(_3003_));
 sky130_fd_sc_hd__and4_1 _3221_ (.A(_2986_),
    .B(_2990_),
    .C(_3000_),
    .D(_3003_),
    .X(_3004_));
 sky130_fd_sc_hd__o21a_1 _3222_ (.A1(net160),
    .A2(_2987_),
    .B1(_2976_),
    .X(_3005_));
 sky130_fd_sc_hd__o2bb2a_1 _3223_ (.A1_N(_2936_),
    .A2_N(_2988_),
    .B1(_3005_),
    .B2(_2922_),
    .X(_3006_));
 sky130_fd_sc_hd__nand3b_4 _3224_ (.A_N(\z80.tv80s.i_tv80_core.IR[6] ),
    .B(\z80.tv80s.i_tv80_core.IR[7] ),
    .C(net144),
    .Y(_3007_));
 sky130_fd_sc_hd__or2_1 _3225_ (.A(net148),
    .B(_3007_),
    .X(_3008_));
 sky130_fd_sc_hd__o31a_1 _3226_ (.A1(net151),
    .A2(_2928_),
    .A3(_3002_),
    .B1(_3008_),
    .X(_3009_));
 sky130_fd_sc_hd__a31oi_1 _3227_ (.A1(net160),
    .A2(net155),
    .A3(_2845_),
    .B1(_2988_),
    .Y(_3010_));
 sky130_fd_sc_hd__and3_1 _3228_ (.A(_2908_),
    .B(_2964_),
    .C(_2975_),
    .X(_3011_));
 sky130_fd_sc_hd__and3_1 _3229_ (.A(net155),
    .B(net151),
    .C(_2891_),
    .X(_3012_));
 sky130_fd_sc_hd__inv_2 _3230_ (.A(_3012_),
    .Y(_3013_));
 sky130_fd_sc_hd__or3b_1 _3231_ (.A(_3007_),
    .B(net149),
    .C_N(_2939_),
    .X(_3014_));
 sky130_fd_sc_hd__or4_1 _3232_ (.A(_2899_),
    .B(_2972_),
    .C(_2974_),
    .D(_2982_),
    .X(_3015_));
 sky130_fd_sc_hd__o221a_1 _3233_ (.A1(_3009_),
    .A2(_3010_),
    .B1(_3011_),
    .B2(_3002_),
    .C1(_3015_),
    .X(_3016_));
 sky130_fd_sc_hd__o311a_1 _3234_ (.A1(_2846_),
    .A2(_3007_),
    .A3(_3013_),
    .B1(_3014_),
    .C1(_3016_),
    .X(_3017_));
 sky130_fd_sc_hd__and3_1 _3235_ (.A(_3004_),
    .B(_3006_),
    .C(_3017_),
    .X(_3018_));
 sky130_fd_sc_hd__nor2_1 _3236_ (.A(_2901_),
    .B(_2919_),
    .Y(_3019_));
 sky130_fd_sc_hd__or4b_4 _3237_ (.A(net145),
    .B(\z80.tv80s.i_tv80_core.IR[7] ),
    .C(\z80.tv80s.i_tv80_core.IR[6] ),
    .D_N(net149),
    .X(_3020_));
 sky130_fd_sc_hd__nor2_4 _3238_ (.A(_2908_),
    .B(_3020_),
    .Y(_3021_));
 sky130_fd_sc_hd__or2_1 _3239_ (.A(_3019_),
    .B(_3021_),
    .X(_3022_));
 sky130_fd_sc_hd__and2_1 _3240_ (.A(_2908_),
    .B(_2916_),
    .X(_3023_));
 sky130_fd_sc_hd__a211o_1 _3241_ (.A1(_2916_),
    .A2(_2956_),
    .B1(net144),
    .C1(net110),
    .X(_3024_));
 sky130_fd_sc_hd__o21a_1 _3242_ (.A1(_2961_),
    .A2(_3023_),
    .B1(_3024_),
    .X(_3025_));
 sky130_fd_sc_hd__nor2_1 _3243_ (.A(net110),
    .B(_2960_),
    .Y(_3026_));
 sky130_fd_sc_hd__or2_1 _3244_ (.A(net110),
    .B(_2960_),
    .X(_3027_));
 sky130_fd_sc_hd__o22a_1 _3245_ (.A1(_2847_),
    .A2(_2966_),
    .B1(_3027_),
    .B2(_2934_),
    .X(_3028_));
 sky130_fd_sc_hd__nand2_2 _3246_ (.A(net120),
    .B(net149),
    .Y(_3029_));
 sky130_fd_sc_hd__or2_2 _3247_ (.A(_2887_),
    .B(_2907_),
    .X(_3030_));
 sky130_fd_sc_hd__or2_2 _3248_ (.A(_2951_),
    .B(_3020_),
    .X(_3031_));
 sky130_fd_sc_hd__nand2_4 _3249_ (.A(_2900_),
    .B(_2939_),
    .Y(_3032_));
 sky130_fd_sc_hd__nand2_1 _3250_ (.A(_2847_),
    .B(_2949_),
    .Y(_3033_));
 sky130_fd_sc_hd__o22a_1 _3251_ (.A1(_2957_),
    .A2(_2961_),
    .B1(_3029_),
    .B2(_3030_),
    .X(_3034_));
 sky130_fd_sc_hd__and4b_1 _3252_ (.A_N(_3022_),
    .B(_3031_),
    .C(_3032_),
    .D(_3033_),
    .X(_3035_));
 sky130_fd_sc_hd__and3_1 _3253_ (.A(_3028_),
    .B(_3034_),
    .C(_3035_),
    .X(_3036_));
 sky130_fd_sc_hd__nand2_1 _3254_ (.A(_3025_),
    .B(_3036_),
    .Y(_3037_));
 sky130_fd_sc_hd__or2_4 _3255_ (.A(_2903_),
    .B(_3007_),
    .X(_3038_));
 sky130_fd_sc_hd__or2_4 _3256_ (.A(_2960_),
    .B(_3007_),
    .X(_3039_));
 sky130_fd_sc_hd__and2_2 _3257_ (.A(_3038_),
    .B(_3039_),
    .X(_3040_));
 sky130_fd_sc_hd__nand2_2 _3258_ (.A(_3038_),
    .B(_3039_),
    .Y(_3041_));
 sky130_fd_sc_hd__or3b_1 _3259_ (.A(_2899_),
    .B(_2972_),
    .C_N(_2974_),
    .X(_3042_));
 sky130_fd_sc_hd__o32a_1 _3260_ (.A1(net161),
    .A2(_2987_),
    .A3(_3008_),
    .B1(_3013_),
    .B2(_3002_),
    .X(_3043_));
 sky130_fd_sc_hd__and3_1 _3261_ (.A(_3040_),
    .B(_3042_),
    .C(_3043_),
    .X(_3044_));
 sky130_fd_sc_hd__o21ai_1 _3262_ (.A1(_2978_),
    .A2(_2988_),
    .B1(_2921_),
    .Y(_3045_));
 sky130_fd_sc_hd__or4_1 _3263_ (.A(_2844_),
    .B(_2890_),
    .C(_3007_),
    .D(_3029_),
    .X(_3046_));
 sky130_fd_sc_hd__o31a_1 _3264_ (.A1(_2845_),
    .A2(_2928_),
    .A3(_3008_),
    .B1(_3046_),
    .X(_3047_));
 sky130_fd_sc_hd__nor2_1 _3265_ (.A(_2907_),
    .B(_3007_),
    .Y(_3048_));
 sky130_fd_sc_hd__or2_2 _3266_ (.A(_2907_),
    .B(_3007_),
    .X(_3049_));
 sky130_fd_sc_hd__nor2_2 _3267_ (.A(_2918_),
    .B(_3007_),
    .Y(_3050_));
 sky130_fd_sc_hd__or2_2 _3268_ (.A(_2918_),
    .B(_3007_),
    .X(_3051_));
 sky130_fd_sc_hd__nor2_2 _3269_ (.A(_3048_),
    .B(_3050_),
    .Y(_3052_));
 sky130_fd_sc_hd__o311a_1 _3270_ (.A1(net155),
    .A2(_2845_),
    .A3(_3002_),
    .B1(_3047_),
    .C1(_3052_),
    .X(_3053_));
 sky130_fd_sc_hd__a21o_1 _3271_ (.A1(_2911_),
    .A2(_2937_),
    .B1(_3005_),
    .X(_0382_));
 sky130_fd_sc_hd__and4_1 _3272_ (.A(_3044_),
    .B(_3045_),
    .C(_3053_),
    .D(_0382_),
    .X(_0383_));
 sky130_fd_sc_hd__and3_1 _3273_ (.A(_3025_),
    .B(_3036_),
    .C(_0383_),
    .X(_0384_));
 sky130_fd_sc_hd__and3b_1 _3274_ (.A_N(_2970_),
    .B(_3018_),
    .C(_0384_),
    .X(_0385_));
 sky130_fd_sc_hd__o21a_1 _3275_ (.A1(_2851_),
    .A2(_0385_),
    .B1(_2905_),
    .X(_0386_));
 sky130_fd_sc_hd__nor2_1 _3276_ (.A(net164),
    .B(net163),
    .Y(_0387_));
 sky130_fd_sc_hd__or2_2 _3277_ (.A(net164),
    .B(net163),
    .X(_0388_));
 sky130_fd_sc_hd__nor2_1 _3278_ (.A(_3041_),
    .B(_3048_),
    .Y(_0389_));
 sky130_fd_sc_hd__nor2_2 _3279_ (.A(_2903_),
    .B(net108),
    .Y(_0390_));
 sky130_fd_sc_hd__or2_2 _3280_ (.A(_2903_),
    .B(net108),
    .X(_0391_));
 sky130_fd_sc_hd__and3_1 _3281_ (.A(_2927_),
    .B(_2934_),
    .C(_2980_),
    .X(_0392_));
 sky130_fd_sc_hd__or3_2 _3282_ (.A(_2928_),
    .B(_2935_),
    .C(net108),
    .X(_0393_));
 sky130_fd_sc_hd__and3_1 _3283_ (.A(_3051_),
    .B(_0391_),
    .C(_0393_),
    .X(_0394_));
 sky130_fd_sc_hd__or3_2 _3284_ (.A(net159),
    .B(net157),
    .C(net108),
    .X(_0395_));
 sky130_fd_sc_hd__nand4_1 _3285_ (.A(_2994_),
    .B(_0389_),
    .C(_0394_),
    .D(_0395_),
    .Y(_0396_));
 sky130_fd_sc_hd__nor2_4 _3286_ (.A(net131),
    .B(net130),
    .Y(_0397_));
 sky130_fd_sc_hd__or2_4 _3287_ (.A(net132),
    .B(net130),
    .X(_0398_));
 sky130_fd_sc_hd__o21a_1 _3288_ (.A1(_0393_),
    .A2(_0398_),
    .B1(_0396_),
    .X(_0399_));
 sky130_fd_sc_hd__nor2_4 _3289_ (.A(net131),
    .B(net134),
    .Y(_0400_));
 sky130_fd_sc_hd__or2_4 _3290_ (.A(net131),
    .B(net133),
    .X(_0401_));
 sky130_fd_sc_hd__o221a_1 _3291_ (.A1(net135),
    .A2(_0395_),
    .B1(_0401_),
    .B2(_3040_),
    .C1(_2994_),
    .X(_0402_));
 sky130_fd_sc_hd__o221a_1 _3292_ (.A1(net135),
    .A2(_3051_),
    .B1(_0401_),
    .B2(_3049_),
    .C1(_0391_),
    .X(_0403_));
 sky130_fd_sc_hd__a31o_1 _3293_ (.A1(_0399_),
    .A2(_0402_),
    .A3(_0403_),
    .B1(_0388_),
    .X(_0404_));
 sky130_fd_sc_hd__nor2_4 _3294_ (.A(_2847_),
    .B(_3029_),
    .Y(_0405_));
 sky130_fd_sc_hd__nand3b_4 _3295_ (.A_N(net153),
    .B(net148),
    .C(net144),
    .Y(_0406_));
 sky130_fd_sc_hd__nand2_1 _3296_ (.A(net97),
    .B(_0406_),
    .Y(_0407_));
 sky130_fd_sc_hd__nand2_1 _3297_ (.A(_2892_),
    .B(_2995_),
    .Y(_0408_));
 sky130_fd_sc_hd__a41o_1 _3298_ (.A1(net137),
    .A2(_2980_),
    .A3(_0407_),
    .A4(_0408_),
    .B1(net119),
    .X(_0409_));
 sky130_fd_sc_hd__a2bb2o_1 _3299_ (.A1_N(_2886_),
    .A2_N(_2918_),
    .B1(_2982_),
    .B2(_2896_),
    .X(_0410_));
 sky130_fd_sc_hd__or4_1 _3300_ (.A(_2931_),
    .B(_2940_),
    .C(_3021_),
    .D(_0410_),
    .X(_0411_));
 sky130_fd_sc_hd__nor2_2 _3301_ (.A(net110),
    .B(_2903_),
    .Y(_0412_));
 sky130_fd_sc_hd__or2_1 _3302_ (.A(net110),
    .B(_2903_),
    .X(_0413_));
 sky130_fd_sc_hd__a2111o_1 _3303_ (.A1(_2936_),
    .A2(_2939_),
    .B1(_0412_),
    .C1(_2938_),
    .D1(_2933_),
    .X(_0414_));
 sky130_fd_sc_hd__nor2_2 _3304_ (.A(_2897_),
    .B(_2960_),
    .Y(_0415_));
 sky130_fd_sc_hd__or2_2 _3305_ (.A(_2917_),
    .B(_0415_),
    .X(_0416_));
 sky130_fd_sc_hd__and2_1 _3306_ (.A(_3030_),
    .B(_3031_),
    .X(_0417_));
 sky130_fd_sc_hd__nand2_2 _3307_ (.A(_3030_),
    .B(_3031_),
    .Y(_0418_));
 sky130_fd_sc_hd__or2_1 _3308_ (.A(_0416_),
    .B(_0418_),
    .X(_0419_));
 sky130_fd_sc_hd__or2_1 _3309_ (.A(_2946_),
    .B(_2953_),
    .X(_0420_));
 sky130_fd_sc_hd__nor4_1 _3310_ (.A(_0411_),
    .B(_0414_),
    .C(_0419_),
    .D(_0420_),
    .Y(_0421_));
 sky130_fd_sc_hd__nor2_4 _3311_ (.A(_2897_),
    .B(_2977_),
    .Y(_0422_));
 sky130_fd_sc_hd__nor2_1 _3312_ (.A(_2948_),
    .B(_0422_),
    .Y(_0423_));
 sky130_fd_sc_hd__o22a_1 _3313_ (.A1(_2897_),
    .A2(_2907_),
    .B1(_2919_),
    .B2(_2901_),
    .X(_0424_));
 sky130_fd_sc_hd__or2_1 _3314_ (.A(_2949_),
    .B(_3019_),
    .X(_0425_));
 sky130_fd_sc_hd__nor2_1 _3315_ (.A(_2897_),
    .B(_2964_),
    .Y(_0426_));
 sky130_fd_sc_hd__or2_2 _3316_ (.A(_2897_),
    .B(_2964_),
    .X(_0427_));
 sky130_fd_sc_hd__and3_1 _3317_ (.A(_0423_),
    .B(_0424_),
    .C(_0427_),
    .X(_0428_));
 sky130_fd_sc_hd__nor2_1 _3318_ (.A(net110),
    .B(net97),
    .Y(_0429_));
 sky130_fd_sc_hd__or2_2 _3319_ (.A(net110),
    .B(net97),
    .X(_0430_));
 sky130_fd_sc_hd__nand2_1 _3320_ (.A(net120),
    .B(\z80.tv80s.i_tv80_core.i_mcode.MCycle[1] ),
    .Y(_0431_));
 sky130_fd_sc_hd__and3_1 _3321_ (.A(net120),
    .B(net132),
    .C(net96),
    .X(_0432_));
 sky130_fd_sc_hd__and3b_2 _3322_ (.A_N(net158),
    .B(net156),
    .C(_2885_),
    .X(_0433_));
 sky130_fd_sc_hd__or3_4 _3323_ (.A(net158),
    .B(_2844_),
    .C(net110),
    .X(_0434_));
 sky130_fd_sc_hd__nor2_1 _3324_ (.A(_0400_),
    .B(_0406_),
    .Y(_0435_));
 sky130_fd_sc_hd__o221a_1 _3325_ (.A1(_0430_),
    .A2(_0432_),
    .B1(_0434_),
    .B2(_0435_),
    .C1(_2910_),
    .X(_0436_));
 sky130_fd_sc_hd__or3b_4 _3326_ (.A(_2844_),
    .B(_2897_),
    .C_N(_2906_),
    .X(_0437_));
 sky130_fd_sc_hd__inv_2 _3327_ (.A(_0437_),
    .Y(_0438_));
 sky130_fd_sc_hd__nand2_1 _3328_ (.A(_3032_),
    .B(_0437_),
    .Y(_0439_));
 sky130_fd_sc_hd__and4b_1 _3329_ (.A_N(_0439_),
    .B(net108),
    .C(_2945_),
    .D(_0436_),
    .X(_0440_));
 sky130_fd_sc_hd__a31o_1 _3330_ (.A1(net155),
    .A2(net135),
    .A3(_2890_),
    .B1(_2972_),
    .X(_0441_));
 sky130_fd_sc_hd__nand2_1 _3331_ (.A(net145),
    .B(_3026_),
    .Y(_0442_));
 sky130_fd_sc_hd__nand2_1 _3332_ (.A(_2913_),
    .B(_0442_),
    .Y(_0443_));
 sky130_fd_sc_hd__or3_2 _3333_ (.A(net145),
    .B(net135),
    .C(_3027_),
    .X(_0444_));
 sky130_fd_sc_hd__and3b_1 _3334_ (.A_N(_0443_),
    .B(_0444_),
    .C(_0441_),
    .X(_0445_));
 sky130_fd_sc_hd__a41o_1 _3335_ (.A1(_0421_),
    .A2(_0428_),
    .A3(_0440_),
    .A4(_0445_),
    .B1(_0409_),
    .X(_0446_));
 sky130_fd_sc_hd__nand3_4 _3336_ (.A(_0386_),
    .B(_0404_),
    .C(_0446_),
    .Y(_0447_));
 sky130_fd_sc_hd__nor2_1 _3337_ (.A(net133),
    .B(_3052_),
    .Y(_0448_));
 sky130_fd_sc_hd__o21a_1 _3338_ (.A1(net130),
    .A2(\z80.tv80s.i_tv80_core.i_mcode.MCycle[3] ),
    .B1(_2848_),
    .X(_0449_));
 sky130_fd_sc_hd__o21ai_4 _3339_ (.A1(net130),
    .A2(\z80.tv80s.i_tv80_core.i_mcode.MCycle[3] ),
    .B1(_2848_),
    .Y(_0450_));
 sky130_fd_sc_hd__a21oi_1 _3340_ (.A1(_0390_),
    .A2(_0450_),
    .B1(_0448_),
    .Y(_0451_));
 sky130_fd_sc_hd__a31o_1 _3341_ (.A1(_0399_),
    .A2(_0402_),
    .A3(_0451_),
    .B1(_0388_),
    .X(_0452_));
 sky130_fd_sc_hd__o21a_1 _3342_ (.A1(\z80.tv80s.i_tv80_core.i_mcode.MCycle[1] ),
    .A2(_2913_),
    .B1(_0421_),
    .X(_0453_));
 sky130_fd_sc_hd__a21o_1 _3343_ (.A1(\z80.tv80s.i_tv80_core.i_mcode.MCycle[2] ),
    .A2(_0431_),
    .B1(_2888_),
    .X(_0454_));
 sky130_fd_sc_hd__o211a_1 _3344_ (.A1(_2961_),
    .A2(_0449_),
    .B1(_0454_),
    .C1(_3020_),
    .X(_0455_));
 sky130_fd_sc_hd__o211a_1 _3345_ (.A1(_2960_),
    .A2(_0455_),
    .B1(_0453_),
    .C1(_0428_),
    .X(_0456_));
 sky130_fd_sc_hd__o2111a_1 _3346_ (.A1(net149),
    .A2(_0444_),
    .B1(_0456_),
    .C1(_0440_),
    .D1(_0441_),
    .X(_0457_));
 sky130_fd_sc_hd__o211a_2 _3347_ (.A1(_0409_),
    .A2(_0457_),
    .B1(_0452_),
    .C1(_0386_),
    .X(_0458_));
 sky130_fd_sc_hd__or2_1 _3348_ (.A(_2894_),
    .B(_0458_),
    .X(_0459_));
 sky130_fd_sc_hd__a21o_1 _3349_ (.A1(_3039_),
    .A2(_0395_),
    .B1(net135),
    .X(_0460_));
 sky130_fd_sc_hd__nor2_4 _3350_ (.A(_2848_),
    .B(net133),
    .Y(_0461_));
 sky130_fd_sc_hd__nand2_2 _3351_ (.A(net132),
    .B(_2849_),
    .Y(_0462_));
 sky130_fd_sc_hd__or2_1 _3352_ (.A(net135),
    .B(_2994_),
    .X(_0463_));
 sky130_fd_sc_hd__a21o_1 _3353_ (.A1(_3038_),
    .A2(_0463_),
    .B1(_0461_),
    .X(_0464_));
 sky130_fd_sc_hd__nor2_1 _3354_ (.A(_3049_),
    .B(_0461_),
    .Y(_0465_));
 sky130_fd_sc_hd__and4bb_1 _3355_ (.A_N(net166),
    .B_N(_0465_),
    .C(_0394_),
    .D(_0460_),
    .X(_0466_));
 sky130_fd_sc_hd__xnor2_1 _3356_ (.A(net153),
    .B(\z80.tv80s.i_tv80_core.F[0] ),
    .Y(_0467_));
 sky130_fd_sc_hd__and3_1 _3357_ (.A(net153),
    .B(net149),
    .C(_2847_),
    .X(_0468_));
 sky130_fd_sc_hd__nand2b_2 _3358_ (.A_N(net147),
    .B(net154),
    .Y(_0469_));
 sky130_fd_sc_hd__and3b_2 _3359_ (.A_N(net148),
    .B(net144),
    .C(net153),
    .X(_0470_));
 sky130_fd_sc_hd__nor2_2 _3360_ (.A(net151),
    .B(_2935_),
    .Y(_0471_));
 sky130_fd_sc_hd__nor4b_1 _3361_ (.A(net153),
    .B(net148),
    .C(\z80.tv80s.i_tv80_core.F[2] ),
    .D_N(net144),
    .Y(_0472_));
 sky130_fd_sc_hd__a221oi_2 _3362_ (.A1(_3001_),
    .A2(_0467_),
    .B1(_0470_),
    .B2(\z80.tv80s.i_tv80_core.F[2] ),
    .C1(_0472_),
    .Y(_0473_));
 sky130_fd_sc_hd__and3_1 _3363_ (.A(net154),
    .B(net148),
    .C(net144),
    .X(_0474_));
 sky130_fd_sc_hd__nand3_2 _3364_ (.A(net153),
    .B(net148),
    .C(net144),
    .Y(_0475_));
 sky130_fd_sc_hd__mux2_1 _3365_ (.A0(_0406_),
    .A1(_0475_),
    .S(\z80.tv80s.i_tv80_core.F[7] ),
    .X(_0476_));
 sky130_fd_sc_hd__or2_2 _3366_ (.A(net154),
    .B(net147),
    .X(_0477_));
 sky130_fd_sc_hd__o21ba_1 _3367_ (.A1(net153),
    .A2(net148),
    .B1_N(\z80.tv80s.i_tv80_core.F[6] ),
    .X(_0478_));
 sky130_fd_sc_hd__mux2_1 _3368_ (.A0(_0469_),
    .A1(_0477_),
    .S(_2852_),
    .X(_0479_));
 sky130_fd_sc_hd__a211o_1 _3369_ (.A1(\z80.tv80s.i_tv80_core.F[6] ),
    .A2(_0469_),
    .B1(_0478_),
    .C1(net144),
    .X(_0480_));
 sky130_fd_sc_hd__and3_2 _3370_ (.A(_0473_),
    .B(_0476_),
    .C(_0480_),
    .X(_0481_));
 sky130_fd_sc_hd__a31o_1 _3371_ (.A1(net134),
    .A2(_2949_),
    .A3(_0481_),
    .B1(_0400_),
    .X(_0482_));
 sky130_fd_sc_hd__inv_2 _3372_ (.A(_0482_),
    .Y(_0483_));
 sky130_fd_sc_hd__or2_4 _3373_ (.A(\z80.tv80s.i_tv80_core.IntCycle ),
    .B(net621),
    .X(_0484_));
 sky130_fd_sc_hd__inv_2 _3374_ (.A(_0484_),
    .Y(_0485_));
 sky130_fd_sc_hd__a21o_1 _3375_ (.A1(_0401_),
    .A2(_0484_),
    .B1(_2910_),
    .X(_0486_));
 sky130_fd_sc_hd__and4_1 _3376_ (.A(net165),
    .B(_2972_),
    .C(net108),
    .D(_0434_),
    .X(_0487_));
 sky130_fd_sc_hd__nor2_1 _3377_ (.A(net134),
    .B(_2945_),
    .Y(_0488_));
 sky130_fd_sc_hd__or4_1 _3378_ (.A(net133),
    .B(\z80.tv80s.i_tv80_core.i_mcode.MCycle[3] ),
    .C(_2945_),
    .D(_0398_),
    .X(_0489_));
 sky130_fd_sc_hd__and4_1 _3379_ (.A(_0430_),
    .B(_0442_),
    .C(_0487_),
    .D(_0489_),
    .X(_0490_));
 sky130_fd_sc_hd__o2111a_1 _3380_ (.A1(_3032_),
    .A2(_0449_),
    .B1(_0486_),
    .C1(_0490_),
    .D1(_0444_),
    .X(_0491_));
 sky130_fd_sc_hd__a41o_2 _3381_ (.A1(\z80.tv80s.i_tv80_core.i_mcode.MCycle[2] ),
    .A2(_0473_),
    .A3(_0476_),
    .A4(_0480_),
    .B1(_0450_),
    .X(_0492_));
 sky130_fd_sc_hd__nand2_1 _3382_ (.A(_0438_),
    .B(_0492_),
    .Y(_0493_));
 sky130_fd_sc_hd__o211a_1 _3383_ (.A1(_0428_),
    .A2(_0483_),
    .B1(_0491_),
    .C1(_0493_),
    .X(_0494_));
 sky130_fd_sc_hd__a32o_1 _3384_ (.A1(_0396_),
    .A2(_0464_),
    .A3(_0466_),
    .B1(_0494_),
    .B2(_0453_),
    .X(_0495_));
 sky130_fd_sc_hd__or3b_4 _3385_ (.A(net163),
    .B(_2894_),
    .C_N(_0495_),
    .X(_0496_));
 sky130_fd_sc_hd__nand2_1 _3386_ (.A(_0459_),
    .B(_0496_),
    .Y(_0497_));
 sky130_fd_sc_hd__a21oi_2 _3387_ (.A1(_2895_),
    .A2(_0447_),
    .B1(_0497_),
    .Y(_0498_));
 sky130_fd_sc_hd__o21a_1 _3388_ (.A1(_2893_),
    .A2(_2904_),
    .B1(net136),
    .X(_0499_));
 sky130_fd_sc_hd__nor2_1 _3389_ (.A(\z80.tv80s.i_tv80_core.XY_State[1] ),
    .B(net467),
    .Y(_0500_));
 sky130_fd_sc_hd__or2_2 _3390_ (.A(\z80.tv80s.i_tv80_core.XY_State[1] ),
    .B(net467),
    .X(_0501_));
 sky130_fd_sc_hd__o211a_4 _3391_ (.A1(net61),
    .A2(_0499_),
    .B1(net103),
    .C1(_2859_),
    .X(_0502_));
 sky130_fd_sc_hd__or4_1 _3392_ (.A(_2904_),
    .B(_2912_),
    .C(_2926_),
    .D(_2929_),
    .X(_0503_));
 sky130_fd_sc_hd__or3_1 _3393_ (.A(_2962_),
    .B(_0416_),
    .C(_0503_),
    .X(_0504_));
 sky130_fd_sc_hd__or2_1 _3394_ (.A(_0420_),
    .B(_0426_),
    .X(_0505_));
 sky130_fd_sc_hd__o21a_1 _3395_ (.A1(_2897_),
    .A2(net97),
    .B1(_2972_),
    .X(_0506_));
 sky130_fd_sc_hd__or2_1 _3396_ (.A(net109),
    .B(_0429_),
    .X(_0507_));
 sky130_fd_sc_hd__o2111a_1 _3397_ (.A1(_2934_),
    .A2(_3027_),
    .B1(_0430_),
    .C1(_2966_),
    .D1(_2981_),
    .X(_0508_));
 sky130_fd_sc_hd__nand2_1 _3398_ (.A(_0506_),
    .B(_0508_),
    .Y(_0509_));
 sky130_fd_sc_hd__or4_2 _3399_ (.A(_2943_),
    .B(_0504_),
    .C(_0505_),
    .D(_0509_),
    .X(_0510_));
 sky130_fd_sc_hd__o21a_1 _3400_ (.A1(_0418_),
    .A2(_0510_),
    .B1(_2849_),
    .X(_0511_));
 sky130_fd_sc_hd__and2_4 _3401_ (.A(_2848_),
    .B(net130),
    .X(_0512_));
 sky130_fd_sc_hd__nand2_4 _3402_ (.A(_2848_),
    .B(net130),
    .Y(_0513_));
 sky130_fd_sc_hd__nor2_1 _3403_ (.A(_0481_),
    .B(_0513_),
    .Y(_0514_));
 sky130_fd_sc_hd__nor2_1 _3404_ (.A(net134),
    .B(_0514_),
    .Y(_0515_));
 sky130_fd_sc_hd__and2_1 _3405_ (.A(_0438_),
    .B(_0515_),
    .X(_0516_));
 sky130_fd_sc_hd__a21oi_2 _3406_ (.A1(_0398_),
    .A2(_0484_),
    .B1(net133),
    .Y(_0517_));
 sky130_fd_sc_hd__a21o_1 _3407_ (.A1(net134),
    .A2(_0484_),
    .B1(_0517_),
    .X(_0518_));
 sky130_fd_sc_hd__a221o_1 _3408_ (.A1(_0418_),
    .A2(_0512_),
    .B1(_0518_),
    .B2(_2909_),
    .C1(_3021_),
    .X(_0519_));
 sky130_fd_sc_hd__nor2_1 _3409_ (.A(net133),
    .B(_0512_),
    .Y(_0520_));
 sky130_fd_sc_hd__nand2_1 _3410_ (.A(_2945_),
    .B(_3032_),
    .Y(_0521_));
 sky130_fd_sc_hd__nand2_1 _3411_ (.A(_0423_),
    .B(_0424_),
    .Y(_0522_));
 sky130_fd_sc_hd__nor2_1 _3412_ (.A(net137),
    .B(_0432_),
    .Y(_0523_));
 sky130_fd_sc_hd__nor2_1 _3413_ (.A(net110),
    .B(_2919_),
    .Y(_0524_));
 sky130_fd_sc_hd__or2_2 _3414_ (.A(net110),
    .B(_2919_),
    .X(_0525_));
 sky130_fd_sc_hd__a22o_1 _3415_ (.A1(_0433_),
    .A2(_0523_),
    .B1(_0524_),
    .B2(_0400_),
    .X(_0526_));
 sky130_fd_sc_hd__a211o_1 _3416_ (.A1(_0520_),
    .A2(_0521_),
    .B1(_0522_),
    .C1(_0526_),
    .X(_0527_));
 sky130_fd_sc_hd__o41a_1 _3417_ (.A1(_0511_),
    .A2(_0516_),
    .A3(_0519_),
    .A4(_0527_),
    .B1(net165),
    .X(_0528_));
 sky130_fd_sc_hd__o21ai_1 _3418_ (.A1(net157),
    .A2(_3007_),
    .B1(_0393_),
    .Y(_0529_));
 sky130_fd_sc_hd__or2_2 _3419_ (.A(_2991_),
    .B(_0529_),
    .X(_0530_));
 sky130_fd_sc_hd__inv_2 _3420_ (.A(_0530_),
    .Y(_0531_));
 sky130_fd_sc_hd__nor2_1 _3421_ (.A(_2998_),
    .B(_0530_),
    .Y(_0532_));
 sky130_fd_sc_hd__a221o_1 _3422_ (.A1(_2991_),
    .A2(_0400_),
    .B1(_0520_),
    .B2(_0392_),
    .C1(_0532_),
    .X(_0533_));
 sky130_fd_sc_hd__o31a_1 _3423_ (.A1(net133),
    .A2(_3039_),
    .A3(_0512_),
    .B1(_3038_),
    .X(_0534_));
 sky130_fd_sc_hd__or4b_1 _3424_ (.A(_2998_),
    .B(_0448_),
    .C(_0533_),
    .D_N(_0534_),
    .X(_0535_));
 sky130_fd_sc_hd__a21oi_1 _3425_ (.A1(net133),
    .A2(_0532_),
    .B1(net105),
    .Y(_0536_));
 sky130_fd_sc_hd__nand2_2 _3426_ (.A(net131),
    .B(_2984_),
    .Y(_0537_));
 sky130_fd_sc_hd__nor2_1 _3427_ (.A(net97),
    .B(_0537_),
    .Y(_0538_));
 sky130_fd_sc_hd__nor2_1 _3428_ (.A(net137),
    .B(_0538_),
    .Y(_0539_));
 sky130_fd_sc_hd__nand2_1 _3429_ (.A(net163),
    .B(_0539_),
    .Y(_0540_));
 sky130_fd_sc_hd__a21oi_1 _3430_ (.A1(_0535_),
    .A2(_0536_),
    .B1(_0528_),
    .Y(_0541_));
 sky130_fd_sc_hd__and3_1 _3431_ (.A(_2842_),
    .B(_0540_),
    .C(_0541_),
    .X(_0542_));
 sky130_fd_sc_hd__o21a_1 _3432_ (.A1(_0510_),
    .A2(_0522_),
    .B1(_2849_),
    .X(_0543_));
 sky130_fd_sc_hd__nand2_1 _3433_ (.A(_3032_),
    .B(_0417_),
    .Y(_0544_));
 sky130_fd_sc_hd__nor2_1 _3434_ (.A(_3021_),
    .B(_0544_),
    .Y(_0545_));
 sky130_fd_sc_hd__o21a_1 _3435_ (.A1(_3021_),
    .A2(_0544_),
    .B1(_0520_),
    .X(_0546_));
 sky130_fd_sc_hd__a21oi_1 _3436_ (.A1(_2853_),
    .A2(\z80.tv80s.i_tv80_core.i_mcode.MCycle[4] ),
    .B1(net130),
    .Y(_0547_));
 sky130_fd_sc_hd__o21ai_1 _3437_ (.A1(net131),
    .A2(_0547_),
    .B1(_0488_),
    .Y(_0548_));
 sky130_fd_sc_hd__or2_1 _3438_ (.A(_2923_),
    .B(_0412_),
    .X(_0549_));
 sky130_fd_sc_hd__a211o_1 _3439_ (.A1(_2909_),
    .A2(_0517_),
    .B1(_0526_),
    .C1(_0549_),
    .X(_0550_));
 sky130_fd_sc_hd__or4b_1 _3440_ (.A(_0516_),
    .B(_0546_),
    .C(_0550_),
    .D_N(_0548_),
    .X(_0551_));
 sky130_fd_sc_hd__o21ai_1 _3441_ (.A1(_0543_),
    .A2(_0551_),
    .B1(net165),
    .Y(_0552_));
 sky130_fd_sc_hd__nor2_1 _3442_ (.A(net130),
    .B(_2853_),
    .Y(_0553_));
 sky130_fd_sc_hd__nand2_4 _3443_ (.A(_2848_),
    .B(_0553_),
    .Y(_0554_));
 sky130_fd_sc_hd__nand2_1 _3444_ (.A(_2849_),
    .B(_0554_),
    .Y(_0555_));
 sky130_fd_sc_hd__a21oi_1 _3445_ (.A1(_3039_),
    .A2(_3052_),
    .B1(_0450_),
    .Y(_0556_));
 sky130_fd_sc_hd__nor2_1 _3446_ (.A(_3038_),
    .B(_0554_),
    .Y(_0557_));
 sky130_fd_sc_hd__nor2_2 _3447_ (.A(_0393_),
    .B(_0513_),
    .Y(_0558_));
 sky130_fd_sc_hd__a2111o_1 _3448_ (.A1(net132),
    .A2(_2991_),
    .B1(_2998_),
    .C1(_0557_),
    .D1(net133),
    .X(_0559_));
 sky130_fd_sc_hd__or3_1 _3449_ (.A(_0556_),
    .B(_0558_),
    .C(_0559_),
    .X(_0560_));
 sky130_fd_sc_hd__or2_1 _3450_ (.A(net105),
    .B(_0560_),
    .X(_0561_));
 sky130_fd_sc_hd__a31o_1 _3451_ (.A1(_0540_),
    .A2(_0552_),
    .A3(_0561_),
    .B1(net129),
    .X(_0562_));
 sky130_fd_sc_hd__o21ai_1 _3452_ (.A1(_0510_),
    .A2(_0522_),
    .B1(net134),
    .Y(_0563_));
 sky130_fd_sc_hd__o22a_1 _3453_ (.A1(_2910_),
    .A2(_0517_),
    .B1(_0525_),
    .B2(_0400_),
    .X(_0564_));
 sky130_fd_sc_hd__o221ai_1 _3454_ (.A1(_0434_),
    .A2(_0523_),
    .B1(_0545_),
    .B2(_0520_),
    .C1(_0564_),
    .Y(_0565_));
 sky130_fd_sc_hd__o21ai_1 _3455_ (.A1(_0437_),
    .A2(_0515_),
    .B1(_0563_),
    .Y(_0566_));
 sky130_fd_sc_hd__or4_1 _3456_ (.A(_2944_),
    .B(_0549_),
    .C(_0565_),
    .D(_0566_),
    .X(_0567_));
 sky130_fd_sc_hd__or2_1 _3457_ (.A(_2851_),
    .B(_0539_),
    .X(_0568_));
 sky130_fd_sc_hd__a21bo_1 _3458_ (.A1(net106),
    .A2(_0560_),
    .B1_N(_0568_),
    .X(_0569_));
 sky130_fd_sc_hd__a311oi_2 _3459_ (.A1(net165),
    .A2(_0548_),
    .A3(_0567_),
    .B1(_0569_),
    .C1(net129),
    .Y(_0570_));
 sky130_fd_sc_hd__and3b_1 _3460_ (.A_N(_0542_),
    .B(_0570_),
    .C(net122),
    .X(_0571_));
 sky130_fd_sc_hd__a21o_1 _3461_ (.A1(net265),
    .A2(_0542_),
    .B1(_0571_),
    .X(_0572_));
 sky130_fd_sc_hd__mux2_1 _3462_ (.A0(net297),
    .A1(net363),
    .S(_0542_),
    .X(_0573_));
 sky130_fd_sc_hd__mux2_1 _3463_ (.A0(_0572_),
    .A1(_0573_),
    .S(_0562_),
    .X(_0574_));
 sky130_fd_sc_hd__or4_1 _3464_ (.A(_2860_),
    .B(_0542_),
    .C(_0562_),
    .D(_0570_),
    .X(_0575_));
 sky130_fd_sc_hd__and2b_4 _3465_ (.A_N(_0574_),
    .B(_0575_),
    .X(_0576_));
 sky130_fd_sc_hd__inv_6 _3466_ (.A(net60),
    .Y(_0577_));
 sky130_fd_sc_hd__nor2_1 _3467_ (.A(_2856_),
    .B(net17),
    .Y(_0578_));
 sky130_fd_sc_hd__nor2_1 _3468_ (.A(net60),
    .B(_0578_),
    .Y(_0579_));
 sky130_fd_sc_hd__nand2_4 _3469_ (.A(_2858_),
    .B(_0579_),
    .Y(_0580_));
 sky130_fd_sc_hd__inv_2 _3470_ (.A(_0580_),
    .Y(_0581_));
 sky130_fd_sc_hd__nand2_4 _3471_ (.A(_0502_),
    .B(_0581_),
    .Y(_0582_));
 sky130_fd_sc_hd__nor2_2 _3472_ (.A(_2893_),
    .B(_0582_),
    .Y(_0583_));
 sky130_fd_sc_hd__and2_1 _3473_ (.A(_2842_),
    .B(net609),
    .X(_0584_));
 sky130_fd_sc_hd__a22o_1 _3474_ (.A1(net499),
    .A2(_0582_),
    .B1(_0583_),
    .B2(_0584_),
    .X(_0008_));
 sky130_fd_sc_hd__nor2_1 _3475_ (.A(net129),
    .B(net609),
    .Y(_0585_));
 sky130_fd_sc_hd__and2_1 _3476_ (.A(_0583_),
    .B(_0585_),
    .X(_0586_));
 sky130_fd_sc_hd__and4_1 _3477_ (.A(_2853_),
    .B(_2857_),
    .C(_0397_),
    .D(_0586_),
    .X(_0587_));
 sky130_fd_sc_hd__a21o_1 _3478_ (.A1(net257),
    .A2(_0582_),
    .B1(_0587_),
    .X(_0009_));
 sky130_fd_sc_hd__a22o_1 _3479_ (.A1(net399),
    .A2(_0582_),
    .B1(_0586_),
    .B2(\z80.tv80s.i_tv80_core.i_mcode.MCycle[4] ),
    .X(_0010_));
 sky130_fd_sc_hd__nor2_1 _3480_ (.A(\z80.tv80s.i_tv80_core.i_mcode.MCycle[3] ),
    .B(net523),
    .Y(_0588_));
 sky130_fd_sc_hd__and3_1 _3481_ (.A(net130),
    .B(_0586_),
    .C(net524),
    .X(_0589_));
 sky130_fd_sc_hd__a21o_1 _3482_ (.A1(net267),
    .A2(_0582_),
    .B1(_0589_),
    .X(_0011_));
 sky130_fd_sc_hd__a22o_1 _3483_ (.A1(net521),
    .A2(_0582_),
    .B1(_0583_),
    .B2(net129),
    .X(_0012_));
 sky130_fd_sc_hd__or4_1 _3484_ (.A(net257),
    .B(net399),
    .C(net267),
    .D(net521),
    .X(_0590_));
 sky130_fd_sc_hd__a221o_1 _3485_ (.A1(net129),
    .A2(_0583_),
    .B1(_0590_),
    .B2(_0582_),
    .C1(_0587_),
    .X(_0591_));
 sky130_fd_sc_hd__a211o_1 _3486_ (.A1(net523),
    .A2(_0586_),
    .B1(_0589_),
    .C1(net652),
    .X(_0029_));
 sky130_fd_sc_hd__and2b_1 _3487_ (.A_N(_0585_),
    .B(_0583_),
    .X(_0592_));
 sky130_fd_sc_hd__nand2_1 _3488_ (.A(_0585_),
    .B(net524),
    .Y(_0593_));
 sky130_fd_sc_hd__nor3_1 _3489_ (.A(_2848_),
    .B(net130),
    .C(_0593_),
    .Y(_0594_));
 sky130_fd_sc_hd__o211a_1 _3490_ (.A1(_2893_),
    .A2(_0594_),
    .B1(_0581_),
    .C1(_0502_),
    .X(_0595_));
 sky130_fd_sc_hd__o41a_1 _3491_ (.A1(net499),
    .A2(net267),
    .A3(net521),
    .A4(net259),
    .B1(_0582_),
    .X(_0596_));
 sky130_fd_sc_hd__or4_1 _3492_ (.A(_0589_),
    .B(_0592_),
    .C(_0595_),
    .D(_0596_),
    .X(_0030_));
 sky130_fd_sc_hd__or4_1 _3493_ (.A(net499),
    .B(net399),
    .C(net521),
    .D(net255),
    .X(_0597_));
 sky130_fd_sc_hd__a22o_1 _3494_ (.A1(_0583_),
    .A2(net525),
    .B1(_0597_),
    .B2(_0582_),
    .X(_0031_));
 sky130_fd_sc_hd__o31a_4 _3495_ (.A1(net122),
    .A2(net573),
    .A3(\z80.tv80s.i_tv80_core.ts[2] ),
    .B1(net136),
    .X(_0598_));
 sky130_fd_sc_hd__a31o_1 _3496_ (.A1(_2854_),
    .A2(_2855_),
    .A3(_2856_),
    .B1(_2849_),
    .X(_0599_));
 sky130_fd_sc_hd__and2_1 _3497_ (.A(net164),
    .B(_2904_),
    .X(_0600_));
 sky130_fd_sc_hd__a31o_1 _3498_ (.A1(net609),
    .A2(net164),
    .A3(_2904_),
    .B1(net101),
    .X(_0601_));
 sky130_fd_sc_hd__nor2_1 _3499_ (.A(net124),
    .B(net101),
    .Y(_0602_));
 sky130_fd_sc_hd__and2_4 _3500_ (.A(net860),
    .B(net17),
    .X(_0603_));
 sky130_fd_sc_hd__nand2_8 _3501_ (.A(net829),
    .B(net17),
    .Y(_0604_));
 sky130_fd_sc_hd__a21oi_4 _3502_ (.A1(net101),
    .A2(_0604_),
    .B1(net746),
    .Y(_0605_));
 sky130_fd_sc_hd__nand2_1 _3503_ (.A(_0601_),
    .B(_0605_),
    .Y(_0606_));
 sky130_fd_sc_hd__nor2_2 _3504_ (.A(_2849_),
    .B(_0604_),
    .Y(_0607_));
 sky130_fd_sc_hd__and3_1 _3505_ (.A(net136),
    .B(net113),
    .C(_0603_),
    .X(_0608_));
 sky130_fd_sc_hd__nand2_1 _3506_ (.A(net113),
    .B(_0607_),
    .Y(_0609_));
 sky130_fd_sc_hd__and2_1 _3507_ (.A(net164),
    .B(_2941_),
    .X(_0610_));
 sky130_fd_sc_hd__nor2_1 _3508_ (.A(_0600_),
    .B(_0610_),
    .Y(_0611_));
 sky130_fd_sc_hd__o41a_1 _3509_ (.A1(net163),
    .A2(net567),
    .A3(net478),
    .A4(_0611_),
    .B1(_0608_),
    .X(_0612_));
 sky130_fd_sc_hd__a221o_1 _3510_ (.A1(net164),
    .A2(_0606_),
    .B1(_0610_),
    .B2(net795),
    .C1(_0612_),
    .X(_0000_));
 sky130_fd_sc_hd__nand2_1 _3511_ (.A(net148),
    .B(_0467_),
    .Y(_0613_));
 sky130_fd_sc_hd__nand3_2 _3512_ (.A(net132),
    .B(_0479_),
    .C(_0613_),
    .Y(_0614_));
 sky130_fd_sc_hd__o2bb2a_1 _3513_ (.A1_N(\z80.tv80s.i_tv80_core.IR[7] ),
    .A2_N(_2982_),
    .B1(_3027_),
    .B2(net144),
    .X(_0615_));
 sky130_fd_sc_hd__or3_1 _3514_ (.A(_2892_),
    .B(_2981_),
    .C(_0406_),
    .X(_0616_));
 sky130_fd_sc_hd__o221a_1 _3515_ (.A1(_0405_),
    .A2(_0430_),
    .B1(_0614_),
    .B2(_3030_),
    .C1(_0616_),
    .X(_0617_));
 sky130_fd_sc_hd__a21o_1 _3516_ (.A1(_0615_),
    .A2(_0617_),
    .B1(net118),
    .X(_0618_));
 sky130_fd_sc_hd__a21oi_1 _3517_ (.A1(net165),
    .A2(_0406_),
    .B1(net163),
    .Y(_0619_));
 sky130_fd_sc_hd__o32a_1 _3518_ (.A1(net108),
    .A2(net97),
    .A3(_0619_),
    .B1(_0395_),
    .B2(net105),
    .X(_0620_));
 sky130_fd_sc_hd__a21oi_1 _3519_ (.A1(_0618_),
    .A2(_0620_),
    .B1(net124),
    .Y(_0621_));
 sky130_fd_sc_hd__a21o_1 _3520_ (.A1(net124),
    .A2(net279),
    .B1(_0621_),
    .X(_0014_));
 sky130_fd_sc_hd__a21oi_1 _3521_ (.A1(_0481_),
    .A2(_0512_),
    .B1(_0437_),
    .Y(_0622_));
 sky130_fd_sc_hd__and3b_2 _3522_ (.A_N(\z80.tv80s.i_tv80_core.NMICycle ),
    .B(_2909_),
    .C(\z80.tv80s.i_tv80_core.IntCycle ),
    .X(_0623_));
 sky130_fd_sc_hd__nor2_2 _3523_ (.A(net118),
    .B(net124),
    .Y(_0624_));
 sky130_fd_sc_hd__o41a_1 _3524_ (.A1(_2962_),
    .A2(_0521_),
    .A3(_0622_),
    .A4(_0623_),
    .B1(_0624_),
    .X(_0625_));
 sky130_fd_sc_hd__nor2_2 _3525_ (.A(net124),
    .B(net105),
    .Y(_0626_));
 sky130_fd_sc_hd__a221o_1 _3526_ (.A1(net124),
    .A2(net548),
    .B1(_0390_),
    .B2(_0626_),
    .C1(_0625_),
    .X(_0015_));
 sky130_fd_sc_hd__and3_1 _3527_ (.A(net164),
    .B(_2941_),
    .C(_0608_),
    .X(_0627_));
 sky130_fd_sc_hd__a22o_1 _3528_ (.A1(net567),
    .A2(_0609_),
    .B1(_0627_),
    .B2(_2934_),
    .X(_0001_));
 sky130_fd_sc_hd__a211o_1 _3529_ (.A1(_0405_),
    .A2(_0433_),
    .B1(_0415_),
    .C1(_2948_),
    .X(_0628_));
 sky130_fd_sc_hd__or3b_1 _3530_ (.A(_2893_),
    .B(_0628_),
    .C_N(_3031_),
    .X(_0629_));
 sky130_fd_sc_hd__a2111o_1 _3531_ (.A1(_2849_),
    .A2(_2949_),
    .B1(_0426_),
    .C1(_0524_),
    .D1(_0629_),
    .X(_0630_));
 sky130_fd_sc_hd__and3b_1 _3532_ (.A_N(_0481_),
    .B(_2949_),
    .C(net134),
    .X(_0631_));
 sky130_fd_sc_hd__a211o_1 _3533_ (.A1(\z80.tv80s.i_tv80_core.NMICycle ),
    .A2(_2909_),
    .B1(_2965_),
    .C1(_0422_),
    .X(_0632_));
 sky130_fd_sc_hd__or4_1 _3534_ (.A(_2914_),
    .B(_3022_),
    .C(_0631_),
    .D(_0632_),
    .X(_0633_));
 sky130_fd_sc_hd__a2111o_1 _3535_ (.A1(net150),
    .A2(_2912_),
    .B1(_2917_),
    .C1(_0630_),
    .D1(_0633_),
    .X(_0634_));
 sky130_fd_sc_hd__a31o_1 _3536_ (.A1(_0438_),
    .A2(_0481_),
    .A3(_0512_),
    .B1(_0634_),
    .X(_0635_));
 sky130_fd_sc_hd__or3_1 _3537_ (.A(_2851_),
    .B(net109),
    .C(net97),
    .X(_0636_));
 sky130_fd_sc_hd__a21oi_1 _3538_ (.A1(_2992_),
    .A2(_2994_),
    .B1(net105),
    .Y(_0637_));
 sky130_fd_sc_hd__a21oi_1 _3539_ (.A1(net165),
    .A2(_0635_),
    .B1(_0637_),
    .Y(_0638_));
 sky130_fd_sc_hd__a21oi_1 _3540_ (.A1(_0636_),
    .A2(_0638_),
    .B1(net124),
    .Y(_0639_));
 sky130_fd_sc_hd__and3b_1 _3541_ (.A_N(_3030_),
    .B(_0614_),
    .C(_0624_),
    .X(_0640_));
 sky130_fd_sc_hd__a211o_1 _3542_ (.A1(net124),
    .A2(net412),
    .B1(_0639_),
    .C1(_0640_),
    .X(_0016_));
 sky130_fd_sc_hd__a32o_1 _3543_ (.A1(_2889_),
    .A2(_2959_),
    .A3(_0624_),
    .B1(net819),
    .B2(net124),
    .X(_0641_));
 sky130_fd_sc_hd__a21o_1 _3544_ (.A1(_0529_),
    .A2(_0626_),
    .B1(_0641_),
    .X(_0013_));
 sky130_fd_sc_hd__a21o_1 _3545_ (.A1(net259),
    .A2(_0582_),
    .B1(_0595_),
    .X(_0007_));
 sky130_fd_sc_hd__a32o_1 _3546_ (.A1(\z80.tv80s.i_tv80_core.i_mcode.MCycle[3] ),
    .A2(_2857_),
    .A3(_0586_),
    .B1(_0582_),
    .B2(net255),
    .X(_0006_));
 sky130_fd_sc_hd__and3_1 _3547_ (.A(net156),
    .B(net151),
    .C(_2890_),
    .X(_0642_));
 sky130_fd_sc_hd__a31o_1 _3548_ (.A1(net148),
    .A2(_2997_),
    .A3(_0642_),
    .B1(_2996_),
    .X(_0643_));
 sky130_fd_sc_hd__and3_1 _3549_ (.A(_2846_),
    .B(net109),
    .C(_2982_),
    .X(_0644_));
 sky130_fd_sc_hd__and3_1 _3550_ (.A(net147),
    .B(_2892_),
    .C(net109),
    .X(_0645_));
 sky130_fd_sc_hd__o31ai_1 _3551_ (.A1(_0643_),
    .A2(_0644_),
    .A3(_0645_),
    .B1(_0626_),
    .Y(_0646_));
 sky130_fd_sc_hd__a22o_1 _3552_ (.A1(_0626_),
    .A2(_0643_),
    .B1(_0646_),
    .B2(net585),
    .X(_0004_));
 sky130_fd_sc_hd__a22o_1 _3553_ (.A1(_0626_),
    .A2(_0645_),
    .B1(_0646_),
    .B2(net269),
    .X(_0005_));
 sky130_fd_sc_hd__and2_1 _3554_ (.A(net478),
    .B(_0609_),
    .X(_0003_));
 sky130_fd_sc_hd__a32o_1 _3555_ (.A1(net609),
    .A2(_0600_),
    .A3(_0602_),
    .B1(_0609_),
    .B2(net163),
    .X(_0647_));
 sky130_fd_sc_hd__a21o_1 _3556_ (.A1(_0600_),
    .A2(_0608_),
    .B1(_0647_),
    .X(_0002_));
 sky130_fd_sc_hd__or3_1 _3557_ (.A(net131),
    .B(_2945_),
    .C(_0547_),
    .X(_0648_));
 sky130_fd_sc_hd__nand2_1 _3558_ (.A(_2909_),
    .B(_0484_),
    .Y(_0649_));
 sky130_fd_sc_hd__a21o_1 _3559_ (.A1(_0423_),
    .A2(_0649_),
    .B1(_0397_),
    .X(_0650_));
 sky130_fd_sc_hd__a21o_1 _3560_ (.A1(_0648_),
    .A2(_0650_),
    .B1(net133),
    .X(_0651_));
 sky130_fd_sc_hd__nor2_1 _3561_ (.A(net134),
    .B(_0513_),
    .Y(_0652_));
 sky130_fd_sc_hd__or2_4 _3562_ (.A(net133),
    .B(_0513_),
    .X(_0653_));
 sky130_fd_sc_hd__o2bb2a_1 _3563_ (.A1_N(\z80.tv80s.i_tv80_core.i_mcode.MCycle[2] ),
    .A2_N(_0429_),
    .B1(_0434_),
    .B2(_0653_),
    .X(_0654_));
 sky130_fd_sc_hd__o22a_1 _3564_ (.A1(_3020_),
    .A2(_0462_),
    .B1(_0554_),
    .B2(_2888_),
    .X(_0655_));
 sky130_fd_sc_hd__o32a_1 _3565_ (.A1(_2899_),
    .A2(_3027_),
    .A3(_0431_),
    .B1(_0654_),
    .B2(_0406_),
    .X(_0656_));
 sky130_fd_sc_hd__o2bb2a_1 _3566_ (.A1_N(_2914_),
    .A2_N(_0512_),
    .B1(_0655_),
    .B2(_2975_),
    .X(_0657_));
 sky130_fd_sc_hd__and3_1 _3567_ (.A(net108),
    .B(_0656_),
    .C(_0657_),
    .X(_0658_));
 sky130_fd_sc_hd__nor2_1 _3568_ (.A(_0398_),
    .B(_0588_),
    .Y(_0659_));
 sky130_fd_sc_hd__or2_1 _3569_ (.A(_0398_),
    .B(_0588_),
    .X(_0660_));
 sky130_fd_sc_hd__nand2_1 _3570_ (.A(net120),
    .B(_2962_),
    .Y(_0661_));
 sky130_fd_sc_hd__a31o_1 _3571_ (.A1(_3032_),
    .A2(_0437_),
    .A3(_0661_),
    .B1(_0660_),
    .X(_0662_));
 sky130_fd_sc_hd__a21oi_1 _3572_ (.A1(net97),
    .A2(_0432_),
    .B1(net108),
    .Y(_0663_));
 sky130_fd_sc_hd__a311o_1 _3573_ (.A1(_0651_),
    .A2(_0658_),
    .A3(_0662_),
    .B1(_0663_),
    .C1(net118),
    .X(_0664_));
 sky130_fd_sc_hd__or3_1 _3574_ (.A(\z80.tv80s.i_tv80_core.i_mcode.MCycle[6] ),
    .B(_0636_),
    .C(_0653_),
    .X(_0665_));
 sky130_fd_sc_hd__nand2_1 _3575_ (.A(net120),
    .B(_0390_),
    .Y(_0666_));
 sky130_fd_sc_hd__or2_1 _3576_ (.A(_0393_),
    .B(_0554_),
    .X(_0667_));
 sky130_fd_sc_hd__o311a_1 _3577_ (.A1(_2918_),
    .A2(net108),
    .A3(_0462_),
    .B1(_0667_),
    .C1(net106),
    .X(_0668_));
 sky130_fd_sc_hd__o221a_1 _3578_ (.A1(_0389_),
    .A2(_0653_),
    .B1(_0660_),
    .B2(_0666_),
    .C1(_0668_),
    .X(_0669_));
 sky130_fd_sc_hd__a31o_4 _3579_ (.A1(_0388_),
    .A2(_0664_),
    .A3(_0665_),
    .B1(_0669_),
    .X(net26));
 sky130_fd_sc_hd__or2_2 _3580_ (.A(net105),
    .B(_0513_),
    .X(_0670_));
 sky130_fd_sc_hd__nor2_1 _3581_ (.A(net135),
    .B(_3040_),
    .Y(_0671_));
 sky130_fd_sc_hd__a2111o_2 _3582_ (.A1(_3049_),
    .A2(_3051_),
    .B1(net105),
    .C1(_0513_),
    .D1(net135),
    .X(_0672_));
 sky130_fd_sc_hd__o31a_1 _3583_ (.A1(net137),
    .A2(_3040_),
    .A3(_0670_),
    .B1(_0672_),
    .X(_0673_));
 sky130_fd_sc_hd__a211o_1 _3584_ (.A1(_3040_),
    .A2(_3051_),
    .B1(_0670_),
    .C1(net135),
    .X(_0674_));
 sky130_fd_sc_hd__o221a_1 _3585_ (.A1(net856),
    .A2(_0672_),
    .B1(_0674_),
    .B2(_2852_),
    .C1(net147),
    .X(_0675_));
 sky130_fd_sc_hd__nor2_1 _3586_ (.A(_0673_),
    .B(_0675_),
    .Y(_0028_));
 sky130_fd_sc_hd__nor2_1 _3587_ (.A(net120),
    .B(_0393_),
    .Y(_0676_));
 sky130_fd_sc_hd__nand2_1 _3588_ (.A(net132),
    .B(_0676_),
    .Y(_0677_));
 sky130_fd_sc_hd__nor2_1 _3589_ (.A(_2992_),
    .B(_0397_),
    .Y(_0678_));
 sky130_fd_sc_hd__nand2_1 _3590_ (.A(_2991_),
    .B(_0398_),
    .Y(_0679_));
 sky130_fd_sc_hd__o311a_1 _3591_ (.A1(net135),
    .A2(_3051_),
    .A3(_0450_),
    .B1(_0677_),
    .C1(_0679_),
    .X(_0680_));
 sky130_fd_sc_hd__o31a_1 _3592_ (.A1(net134),
    .A2(_0389_),
    .A3(_0554_),
    .B1(_0680_),
    .X(_0681_));
 sky130_fd_sc_hd__o22a_1 _3593_ (.A1(_2842_),
    .A2(_2893_),
    .B1(_0681_),
    .B2(net164),
    .X(_0682_));
 sky130_fd_sc_hd__nor2_1 _3594_ (.A(net573),
    .B(_0578_),
    .Y(_0683_));
 sky130_fd_sc_hd__nor2_2 _3595_ (.A(_0397_),
    .B(_0525_),
    .Y(_0684_));
 sky130_fd_sc_hd__o2bb2a_4 _3596_ (.A1_N(_3021_),
    .A2_N(_0652_),
    .B1(_0513_),
    .B2(_0417_),
    .X(_0685_));
 sky130_fd_sc_hd__nand2b_1 _3597_ (.A_N(_0684_),
    .B(_0685_),
    .Y(_0686_));
 sky130_fd_sc_hd__o21ai_1 _3598_ (.A1(net163),
    .A2(_0682_),
    .B1(net26),
    .Y(_0687_));
 sky130_fd_sc_hd__a211o_1 _3599_ (.A1(net164),
    .A2(_0686_),
    .B1(_0687_),
    .C1(_0683_),
    .X(_0688_));
 sky130_fd_sc_hd__or2_1 _3600_ (.A(net778),
    .B(_0683_),
    .X(_0689_));
 sky130_fd_sc_hd__mux2_1 _3601_ (.A0(_0688_),
    .A1(_0689_),
    .S(net136),
    .X(_0019_));
 sky130_fd_sc_hd__or2_1 _3602_ (.A(net26),
    .B(_0683_),
    .X(_0690_));
 sky130_fd_sc_hd__nand2_1 _3603_ (.A(_0688_),
    .B(_0690_),
    .Y(_0691_));
 sky130_fd_sc_hd__a21o_1 _3604_ (.A1(_3039_),
    .A2(_0395_),
    .B1(_0462_),
    .X(_0692_));
 sky130_fd_sc_hd__o21a_1 _3605_ (.A1(_3038_),
    .A2(_0653_),
    .B1(_0692_),
    .X(_0693_));
 sky130_fd_sc_hd__o211a_1 _3606_ (.A1(_2928_),
    .A2(_2961_),
    .B1(_3028_),
    .C1(_2924_),
    .X(_0694_));
 sky130_fd_sc_hd__a2111o_1 _3607_ (.A1(_2889_),
    .A2(_2927_),
    .B1(_2940_),
    .C1(_0507_),
    .D1(_2926_),
    .X(_0695_));
 sky130_fd_sc_hd__nor2_1 _3608_ (.A(_0414_),
    .B(_0695_),
    .Y(_0696_));
 sky130_fd_sc_hd__or3_2 _3609_ (.A(_2953_),
    .B(_0422_),
    .C(_0426_),
    .X(_0697_));
 sky130_fd_sc_hd__nor2_1 _3610_ (.A(_2968_),
    .B(_0697_),
    .Y(_0698_));
 sky130_fd_sc_hd__nand3_1 _3611_ (.A(_0694_),
    .B(_0696_),
    .C(_0698_),
    .Y(_0699_));
 sky130_fd_sc_hd__a31o_1 _3612_ (.A1(net150),
    .A2(_2921_),
    .A3(_2927_),
    .B1(_0544_),
    .X(_0700_));
 sky130_fd_sc_hd__a21o_1 _3613_ (.A1(_2948_),
    .A2(_0475_),
    .B1(_0438_),
    .X(_0701_));
 sky130_fd_sc_hd__nor2_1 _3614_ (.A(_2901_),
    .B(_2907_),
    .Y(_0702_));
 sky130_fd_sc_hd__or4_1 _3615_ (.A(_3022_),
    .B(_0700_),
    .C(_0701_),
    .D(_0702_),
    .X(_0703_));
 sky130_fd_sc_hd__a211o_1 _3616_ (.A1(_2899_),
    .A2(_2949_),
    .B1(_0416_),
    .C1(_0703_),
    .X(_0704_));
 sky130_fd_sc_hd__and3_1 _3617_ (.A(_2910_),
    .B(_0506_),
    .C(_0525_),
    .X(_0705_));
 sky130_fd_sc_hd__nand2_1 _3618_ (.A(_0434_),
    .B(_0705_),
    .Y(_0706_));
 sky130_fd_sc_hd__or4_1 _3619_ (.A(net118),
    .B(_2947_),
    .C(_0513_),
    .D(_0706_),
    .X(_0707_));
 sky130_fd_sc_hd__o32a_2 _3620_ (.A1(_0699_),
    .A2(_0704_),
    .A3(_0707_),
    .B1(_0693_),
    .B2(net105),
    .X(_0708_));
 sky130_fd_sc_hd__a21o_1 _3621_ (.A1(_0688_),
    .A2(_0690_),
    .B1(_0708_),
    .X(_0709_));
 sky130_fd_sc_hd__o21ai_1 _3622_ (.A1(net573),
    .A2(_0578_),
    .B1(net778),
    .Y(_0710_));
 sky130_fd_sc_hd__mux2_1 _3623_ (.A0(_0709_),
    .A1(_0710_),
    .S(net136),
    .X(_0017_));
 sky130_fd_sc_hd__nand2_1 _3624_ (.A(net136),
    .B(_2854_),
    .Y(_0711_));
 sky130_fd_sc_hd__a21oi_1 _3625_ (.A1(_0691_),
    .A2(_0708_),
    .B1(net136),
    .Y(_0712_));
 sky130_fd_sc_hd__a31o_1 _3626_ (.A1(net136),
    .A2(_2854_),
    .A3(_0689_),
    .B1(_0712_),
    .X(_0018_));
 sky130_fd_sc_hd__or4_4 _3627_ (.A(net118),
    .B(_2908_),
    .C(_3020_),
    .D(_0400_),
    .X(_0713_));
 sky130_fd_sc_hd__or4_1 _3628_ (.A(\z80.tv80s.i_tv80_core.mcycles[2] ),
    .B(\z80.tv80s.i_tv80_core.mcycles[4] ),
    .C(\z80.tv80s.i_tv80_core.mcycles[5] ),
    .D(\z80.tv80s.i_tv80_core.mcycles[1] ),
    .X(_0714_));
 sky130_fd_sc_hd__nor2_1 _3629_ (.A(_2849_),
    .B(_0714_),
    .Y(_0715_));
 sky130_fd_sc_hd__a221o_1 _3630_ (.A1(net130),
    .A2(net412),
    .B1(\z80.tv80s.i_tv80_core.mcycles[1] ),
    .B2(\z80.tv80s.i_tv80_core.i_mcode.MCycle[3] ),
    .C1(_0715_),
    .X(_0716_));
 sky130_fd_sc_hd__a221o_2 _3631_ (.A1(net131),
    .A2(net279),
    .B1(net548),
    .B2(\z80.tv80s.i_tv80_core.i_mcode.MCycle[4] ),
    .C1(_0716_),
    .X(_0717_));
 sky130_fd_sc_hd__and4_1 _3632_ (.A(net132),
    .B(\z80.tv80s.i_tv80_core.ISet[0] ),
    .C(net429),
    .D(_3021_),
    .X(_0718_));
 sky130_fd_sc_hd__or3_2 _3633_ (.A(net715),
    .B(_0717_),
    .C(_0718_),
    .X(_0719_));
 sky130_fd_sc_hd__nand2_1 _3634_ (.A(_2842_),
    .B(_0719_),
    .Y(_0720_));
 sky130_fd_sc_hd__nor2_2 _3635_ (.A(_0502_),
    .B(_0580_),
    .Y(_0721_));
 sky130_fd_sc_hd__or3_2 _3636_ (.A(_0502_),
    .B(_0580_),
    .C(_0720_),
    .X(_0722_));
 sky130_fd_sc_hd__o211a_1 _3637_ (.A1(net38),
    .A2(_0607_),
    .B1(_0722_),
    .C1(_2860_),
    .X(_0032_));
 sky130_fd_sc_hd__nor3_1 _3638_ (.A(_0600_),
    .B(_0610_),
    .C(_0722_),
    .Y(_0723_));
 sky130_fd_sc_hd__or4_2 _3639_ (.A(net120),
    .B(net118),
    .C(_2903_),
    .D(_2922_),
    .X(_0724_));
 sky130_fd_sc_hd__and3_1 _3640_ (.A(net763),
    .B(\z80.tv80s.i_tv80_core.INT_s ),
    .C(_0724_),
    .X(_0725_));
 sky130_fd_sc_hd__o21a_1 _3641_ (.A1(net518),
    .A2(_0725_),
    .B1(_0723_),
    .X(_0726_));
 sky130_fd_sc_hd__and4_1 _3642_ (.A(net165),
    .B(net122),
    .C(_2915_),
    .D(_2921_),
    .X(_0727_));
 sky130_fd_sc_hd__or2_2 _3643_ (.A(_0463_),
    .B(_0670_),
    .X(_0728_));
 sky130_fd_sc_hd__or3_1 _3644_ (.A(_2856_),
    .B(\z80.tv80s.i_tv80_core.IntE_FF2 ),
    .C(_0728_),
    .X(_0729_));
 sky130_fd_sc_hd__o21ai_1 _3645_ (.A1(net621),
    .A2(_0724_),
    .B1(_0728_),
    .Y(_0730_));
 sky130_fd_sc_hd__a21o_1 _3646_ (.A1(\z80.tv80s.i_tv80_core.ts[2] ),
    .A2(_0730_),
    .B1(net763),
    .X(_0731_));
 sky130_fd_sc_hd__and4bb_1 _3647_ (.A_N(_0726_),
    .B_N(_0727_),
    .C(_0729_),
    .D(net764),
    .X(_0026_));
 sky130_fd_sc_hd__and3b_1 _3648_ (.A_N(net518),
    .B(_0723_),
    .C(_0725_),
    .X(_0732_));
 sky130_fd_sc_hd__o21ba_1 _3649_ (.A1(_2856_),
    .A2(_0724_),
    .B1_N(net842),
    .X(_0733_));
 sky130_fd_sc_hd__nor3_1 _3650_ (.A(_0727_),
    .B(_0732_),
    .C(_0733_),
    .Y(_0027_));
 sky130_fd_sc_hd__a21oi_2 _3651_ (.A1(net746),
    .A2(net221),
    .B1(_0578_),
    .Y(_0734_));
 sky130_fd_sc_hd__and4_1 _3652_ (.A(net165),
    .B(_2892_),
    .C(net109),
    .D(net96),
    .X(_0735_));
 sky130_fd_sc_hd__a32o_1 _3653_ (.A1(_0577_),
    .A2(_0734_),
    .A3(_0735_),
    .B1(_0485_),
    .B2(net711),
    .X(_0024_));
 sky130_fd_sc_hd__o22a_1 _3654_ (.A1(_2849_),
    .A2(_0485_),
    .B1(_0708_),
    .B2(net405),
    .X(_0736_));
 sky130_fd_sc_hd__nor2_1 _3655_ (.A(_0577_),
    .B(net406),
    .Y(_0021_));
 sky130_fd_sc_hd__mux2_4 _3656_ (.A0(\z80.normal_rd_n ),
    .A1(\z80.early_rd_n ),
    .S(net1),
    .X(net49));
 sky130_fd_sc_hd__nor2_1 _3657_ (.A(net2),
    .B(net3),
    .Y(_0737_));
 sky130_fd_sc_hd__and2b_1 _3658_ (.A_N(net3),
    .B(net2),
    .X(_0738_));
 sky130_fd_sc_hd__o22a_4 _3659_ (.A1(\z80.early_iorq_n ),
    .A2(_0737_),
    .B1(_0738_),
    .B2(\z80.normal_iorq_n ),
    .X(net52));
 sky130_fd_sc_hd__mux2_1 _3660_ (.A0(\z80.normal_mreq_n ),
    .A1(\z80.early_mreq_n ),
    .S(net4),
    .X(_0739_));
 sky130_fd_sc_hd__o21bai_1 _3661_ (.A1(net54),
    .A2(_2884_),
    .B1_N(\z80.normal_mreq_n ),
    .Y(_0740_));
 sky130_fd_sc_hd__a22o_2 _3662_ (.A1(_2884_),
    .A2(_0739_),
    .B1(_0740_),
    .B2(\z80.early_mreq_n ),
    .X(net51));
 sky130_fd_sc_hd__nand2_1 _3663_ (.A(net136),
    .B(net122),
    .Y(_0741_));
 sky130_fd_sc_hd__a21o_1 _3664_ (.A1(_2854_),
    .A2(_0604_),
    .B1(_2849_),
    .X(_0033_));
 sky130_fd_sc_hd__or2_2 _3665_ (.A(net136),
    .B(_0690_),
    .X(_0020_));
 sky130_fd_sc_hd__and2_1 _3666_ (.A(net340),
    .B(net60),
    .X(_0022_));
 sky130_fd_sc_hd__o32a_1 _3667_ (.A1(net133),
    .A2(_2994_),
    .A3(_0397_),
    .B1(_0653_),
    .B2(_3049_),
    .X(_0742_));
 sky130_fd_sc_hd__nor2_1 _3668_ (.A(_0401_),
    .B(_0547_),
    .Y(_0743_));
 sky130_fd_sc_hd__o21ai_2 _3669_ (.A1(_2945_),
    .A2(_0743_),
    .B1(net165),
    .Y(_0744_));
 sky130_fd_sc_hd__nand2_1 _3670_ (.A(net149),
    .B(_0412_),
    .Y(_0745_));
 sky130_fd_sc_hd__nor2_1 _3671_ (.A(_0437_),
    .B(_0492_),
    .Y(_0746_));
 sky130_fd_sc_hd__o22a_1 _3672_ (.A1(_0400_),
    .A2(_0423_),
    .B1(_0437_),
    .B2(_0492_),
    .X(_0747_));
 sky130_fd_sc_hd__nor2_1 _3673_ (.A(_3032_),
    .B(_0450_),
    .Y(_0748_));
 sky130_fd_sc_hd__nor2_1 _3674_ (.A(_0400_),
    .B(_0649_),
    .Y(_0749_));
 sky130_fd_sc_hd__o221a_2 _3675_ (.A1(_3032_),
    .A2(_0450_),
    .B1(_0649_),
    .B2(_0400_),
    .C1(_2945_),
    .X(_0750_));
 sky130_fd_sc_hd__a211o_1 _3676_ (.A1(_0424_),
    .A2(_0427_),
    .B1(net134),
    .C1(_0397_),
    .X(_0751_));
 sky130_fd_sc_hd__o221a_2 _3677_ (.A1(_0400_),
    .A2(_0423_),
    .B1(_0437_),
    .B2(_0492_),
    .C1(_0751_),
    .X(_0752_));
 sky130_fd_sc_hd__a31o_1 _3678_ (.A1(_0745_),
    .A2(_0750_),
    .A3(_0752_),
    .B1(_0744_),
    .X(_0753_));
 sky130_fd_sc_hd__o21ai_4 _3679_ (.A1(net105),
    .A2(_0742_),
    .B1(_0753_),
    .Y(_0754_));
 sky130_fd_sc_hd__nand2_1 _3680_ (.A(net146),
    .B(_0412_),
    .Y(_0755_));
 sky130_fd_sc_hd__a31o_1 _3681_ (.A1(_0750_),
    .A2(_0752_),
    .A3(_0755_),
    .B1(_0744_),
    .X(_0756_));
 sky130_fd_sc_hd__a211o_1 _3682_ (.A1(_2994_),
    .A2(_3038_),
    .B1(_0397_),
    .C1(net133),
    .X(_0757_));
 sky130_fd_sc_hd__o21ai_1 _3683_ (.A1(_3039_),
    .A2(_0653_),
    .B1(net106),
    .Y(_0758_));
 sky130_fd_sc_hd__inv_2 _3684_ (.A(_0758_),
    .Y(_0759_));
 sky130_fd_sc_hd__or2_2 _3685_ (.A(_3052_),
    .B(_0462_),
    .X(_0760_));
 sky130_fd_sc_hd__a32oi_4 _3686_ (.A1(_0757_),
    .A2(_0759_),
    .A3(_0760_),
    .B1(_0756_),
    .B2(net105),
    .Y(_0761_));
 sky130_fd_sc_hd__a32o_1 _3687_ (.A1(_0757_),
    .A2(_0759_),
    .A3(_0760_),
    .B1(_0756_),
    .B2(net105),
    .X(_0762_));
 sky130_fd_sc_hd__nand2_2 _3688_ (.A(_0754_),
    .B(_0761_),
    .Y(_0763_));
 sky130_fd_sc_hd__a31oi_4 _3689_ (.A1(_0413_),
    .A2(_0750_),
    .A3(_0752_),
    .B1(_0744_),
    .Y(_0764_));
 sky130_fd_sc_hd__o2bb2a_1 _3690_ (.A1_N(_3049_),
    .A2_N(_0463_),
    .B1(_0398_),
    .B2(net134),
    .X(_0765_));
 sky130_fd_sc_hd__or2_1 _3691_ (.A(net135),
    .B(_3038_),
    .X(_0766_));
 sky130_fd_sc_hd__a21oi_1 _3692_ (.A1(_3051_),
    .A2(_0766_),
    .B1(_0400_),
    .Y(_0767_));
 sky130_fd_sc_hd__or3_2 _3693_ (.A(_0758_),
    .B(_0765_),
    .C(_0767_),
    .X(_0768_));
 sky130_fd_sc_hd__o21a_1 _3694_ (.A1(net106),
    .A2(_0764_),
    .B1(_0768_),
    .X(_0769_));
 sky130_fd_sc_hd__o2111ai_4 _3695_ (.A1(net136),
    .A2(_0603_),
    .B1(_0711_),
    .C1(_0763_),
    .D1(_0769_),
    .Y(_0770_));
 sky130_fd_sc_hd__and2_1 _3696_ (.A(net164),
    .B(_2950_),
    .X(_0771_));
 sky130_fd_sc_hd__and3_4 _3697_ (.A(net164),
    .B(net122),
    .C(_2950_),
    .X(_0772_));
 sky130_fd_sc_hd__nand2_2 _3698_ (.A(net122),
    .B(_0771_),
    .Y(_0773_));
 sky130_fd_sc_hd__and3_2 _3699_ (.A(net164),
    .B(net874),
    .C(_2950_),
    .X(_0774_));
 sky130_fd_sc_hd__nand2_4 _3700_ (.A(net363),
    .B(_0771_),
    .Y(_0775_));
 sky130_fd_sc_hd__nor2_2 _3701_ (.A(_0772_),
    .B(_0774_),
    .Y(_0776_));
 sky130_fd_sc_hd__nand2_1 _3702_ (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[0] ),
    .B(net143),
    .Y(_0777_));
 sky130_fd_sc_hd__nand3_4 _3703_ (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[2] ),
    .B(\z80.tv80s.i_tv80_core.ALU_Op_r[0] ),
    .C(net143),
    .Y(_0778_));
 sky130_fd_sc_hd__or2_4 _3704_ (.A(_2855_),
    .B(net340),
    .X(_0779_));
 sky130_fd_sc_hd__nand2_1 _3705_ (.A(_2861_),
    .B(_0779_),
    .Y(_0780_));
 sky130_fd_sc_hd__o31a_2 _3706_ (.A1(_2861_),
    .A2(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ),
    .A3(_0778_),
    .B1(_0780_),
    .X(_0781_));
 sky130_fd_sc_hd__and2_1 _3707_ (.A(\z80.tv80s.i_tv80_core.Read_To_Reg_r[1] ),
    .B(\z80.tv80s.i_tv80_core.Read_To_Reg_r[2] ),
    .X(_0782_));
 sky130_fd_sc_hd__or3_1 _3708_ (.A(\z80.tv80s.i_tv80_core.Read_To_Reg_r[3] ),
    .B(_2875_),
    .C(_0782_),
    .X(_0783_));
 sky130_fd_sc_hd__or3b_1 _3709_ (.A(net873),
    .B(_0783_),
    .C_N(_0781_),
    .X(_0784_));
 sky130_fd_sc_hd__a31o_4 _3710_ (.A1(_0770_),
    .A2(_0776_),
    .A3(_0784_),
    .B1(net124),
    .X(_0785_));
 sky130_fd_sc_hd__o2111ai_4 _3711_ (.A1(net106),
    .A2(_0764_),
    .B1(_0768_),
    .C1(net122),
    .D1(net136),
    .Y(_0786_));
 sky130_fd_sc_hd__a211oi_4 _3712_ (.A1(_2856_),
    .A2(_0786_),
    .B1(_0762_),
    .C1(_0754_),
    .Y(_0787_));
 sky130_fd_sc_hd__a211o_1 _3713_ (.A1(_2856_),
    .A2(_0786_),
    .B1(_0762_),
    .C1(_0754_),
    .X(_0788_));
 sky130_fd_sc_hd__mux2_2 _3714_ (.A0(\z80.tv80s.i_tv80_core.XY_State[1] ),
    .A1(\z80.tv80s.i_tv80_core.RegAddrA_r[2] ),
    .S(_0788_),
    .X(_0789_));
 sky130_fd_sc_hd__a21oi_4 _3715_ (.A1(_2856_),
    .A2(_0786_),
    .B1(net103),
    .Y(_0790_));
 sky130_fd_sc_hd__a21o_1 _3716_ (.A1(_2856_),
    .A2(_0786_),
    .B1(net103),
    .X(_0791_));
 sky130_fd_sc_hd__nand2_2 _3717_ (.A(_0776_),
    .B(_0791_),
    .Y(_0792_));
 sky130_fd_sc_hd__a21o_1 _3718_ (.A1(_0776_),
    .A2(_0791_),
    .B1(\z80.tv80s.i_tv80_core.Alternate ),
    .X(_0793_));
 sky130_fd_sc_hd__o21a_4 _3719_ (.A1(_0789_),
    .A2(_0792_),
    .B1(_0793_),
    .X(_0794_));
 sky130_fd_sc_hd__o21ai_4 _3720_ (.A1(_0789_),
    .A2(_0792_),
    .B1(_0793_),
    .Y(_0795_));
 sky130_fd_sc_hd__a21o_1 _3721_ (.A1(\z80.tv80s.i_tv80_core.RegAddrA_r[1] ),
    .A2(_0775_),
    .B1(net89),
    .X(_0796_));
 sky130_fd_sc_hd__a211o_1 _3722_ (.A1(_2856_),
    .A2(_0786_),
    .B1(_0761_),
    .C1(net103),
    .X(_0797_));
 sky130_fd_sc_hd__o31ai_2 _3723_ (.A1(_0787_),
    .A2(_0790_),
    .A3(_0796_),
    .B1(_0797_),
    .Y(_0798_));
 sky130_fd_sc_hd__o31a_4 _3724_ (.A1(_0787_),
    .A2(_0790_),
    .A3(_0796_),
    .B1(_0797_),
    .X(_0799_));
 sky130_fd_sc_hd__o21a_1 _3725_ (.A1(\z80.tv80s.i_tv80_core.RegAddrA_r[0] ),
    .A2(_0774_),
    .B1(net86),
    .X(_0800_));
 sky130_fd_sc_hd__o21ai_2 _3726_ (.A1(\z80.tv80s.i_tv80_core.RegAddrA_r[0] ),
    .A2(_0774_),
    .B1(net86),
    .Y(_0801_));
 sky130_fd_sc_hd__a211oi_2 _3727_ (.A1(_2856_),
    .A2(_0786_),
    .B1(_0754_),
    .C1(net103),
    .Y(_0802_));
 sky130_fd_sc_hd__a211o_1 _3728_ (.A1(_2856_),
    .A2(_0786_),
    .B1(_0754_),
    .C1(net103),
    .X(_0803_));
 sky130_fd_sc_hd__a31o_1 _3729_ (.A1(_0788_),
    .A2(_0791_),
    .A3(_0801_),
    .B1(_0802_),
    .X(_0804_));
 sky130_fd_sc_hd__o31a_4 _3730_ (.A1(_0787_),
    .A2(_0790_),
    .A3(_0800_),
    .B1(_0803_),
    .X(_0805_));
 sky130_fd_sc_hd__and3_4 _3731_ (.A(_0795_),
    .B(_0799_),
    .C(net69),
    .X(_0806_));
 sky130_fd_sc_hd__or3_1 _3732_ (.A(_0794_),
    .B(net71),
    .C(net70),
    .X(_0807_));
 sky130_fd_sc_hd__or2_4 _3733_ (.A(_0785_),
    .B(_0807_),
    .X(_0808_));
 sky130_fd_sc_hd__o211a_2 _3734_ (.A1(net136),
    .A2(\z80.tv80s.i_tv80_core.ts[2] ),
    .B1(_0711_),
    .C1(_0769_),
    .X(_0809_));
 sky130_fd_sc_hd__inv_2 _3735_ (.A(net76),
    .Y(_0810_));
 sky130_fd_sc_hd__and4_2 _3736_ (.A(net166),
    .B(_2980_),
    .C(net97),
    .D(_0406_),
    .X(_0811_));
 sky130_fd_sc_hd__inv_4 _3737_ (.A(_0811_),
    .Y(_0812_));
 sky130_fd_sc_hd__and2_1 _3738_ (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ),
    .B(_0778_),
    .X(_0813_));
 sky130_fd_sc_hd__nand2_4 _3739_ (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ),
    .B(_0778_),
    .Y(_0814_));
 sky130_fd_sc_hd__and2_4 _3740_ (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[2] ),
    .B(_2863_),
    .X(_0815_));
 sky130_fd_sc_hd__xor2_2 _3741_ (.A(net143),
    .B(\z80.tv80s.i_tv80_core.BusB[0] ),
    .X(_0816_));
 sky130_fd_sc_hd__and2_1 _3742_ (.A(\z80.tv80s.i_tv80_core.BusA[0] ),
    .B(_0816_),
    .X(_0817_));
 sky130_fd_sc_hd__or2_1 _3743_ (.A(net143),
    .B(_0817_),
    .X(_0818_));
 sky130_fd_sc_hd__xor2_2 _3744_ (.A(\z80.tv80s.i_tv80_core.BusA[0] ),
    .B(_0816_),
    .X(_0819_));
 sky130_fd_sc_hd__and2b_1 _3745_ (.A_N(\z80.tv80s.i_tv80_core.ALU_Op_r[2] ),
    .B(\z80.tv80s.i_tv80_core.F[0] ),
    .X(_0820_));
 sky130_fd_sc_hd__nor2_1 _3746_ (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[0] ),
    .B(\z80.tv80s.i_tv80_core.ALU_Op_r[1] ),
    .Y(_0821_));
 sky130_fd_sc_hd__xor2_1 _3747_ (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[0] ),
    .B(net143),
    .X(_0822_));
 sky130_fd_sc_hd__mux2_1 _3748_ (.A0(net143),
    .A1(_0822_),
    .S(_0820_),
    .X(_0823_));
 sky130_fd_sc_hd__or2_1 _3749_ (.A(_0819_),
    .B(_0823_),
    .X(_0824_));
 sky130_fd_sc_hd__nand2_1 _3750_ (.A(_0819_),
    .B(_0823_),
    .Y(_0825_));
 sky130_fd_sc_hd__and2_2 _3751_ (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[2] ),
    .B(_0777_),
    .X(_0826_));
 sky130_fd_sc_hd__nand2_4 _3752_ (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[2] ),
    .B(_0777_),
    .Y(_0827_));
 sky130_fd_sc_hd__and3_2 _3753_ (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[2] ),
    .B(\z80.tv80s.i_tv80_core.ALU_Op_r[0] ),
    .C(net111),
    .X(_0828_));
 sky130_fd_sc_hd__a22o_1 _3754_ (.A1(_0815_),
    .A2(_0818_),
    .B1(_0819_),
    .B2(_0828_),
    .X(_0829_));
 sky130_fd_sc_hd__a31o_1 _3755_ (.A1(_0824_),
    .A2(_0825_),
    .A3(_0827_),
    .B1(_0829_),
    .X(_0830_));
 sky130_fd_sc_hd__o41a_1 _3756_ (.A1(net111),
    .A2(\z80.tv80s.i_tv80_core.BusA[0] ),
    .A3(\z80.tv80s.i_tv80_core.BusB[0] ),
    .A4(_0827_),
    .B1(_0830_),
    .X(_0831_));
 sky130_fd_sc_hd__and3b_1 _3757_ (.A_N(\z80.tv80s.i_tv80_core.ALU_Op_r[2] ),
    .B(net143),
    .C(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ),
    .X(_0832_));
 sky130_fd_sc_hd__or3_2 _3758_ (.A(_2862_),
    .B(\z80.tv80s.i_tv80_core.ALU_Op_r[2] ),
    .C(net111),
    .X(_0833_));
 sky130_fd_sc_hd__nor2_4 _3759_ (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[0] ),
    .B(_0833_),
    .Y(_0834_));
 sky130_fd_sc_hd__nor2_1 _3760_ (.A(net153),
    .B(_2899_),
    .Y(_0835_));
 sky130_fd_sc_hd__nand2_2 _3761_ (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[0] ),
    .B(_0832_),
    .Y(_0836_));
 sky130_fd_sc_hd__inv_2 _3762_ (.A(_0836_),
    .Y(_0837_));
 sky130_fd_sc_hd__o311a_1 _3763_ (.A1(net153),
    .A2(_2863_),
    .A3(_2899_),
    .B1(_0832_),
    .C1(\z80.tv80s.i_tv80_core.BusB[0] ),
    .X(_0838_));
 sky130_fd_sc_hd__and3b_4 _3764_ (.A_N(\z80.tv80s.i_tv80_core.ALU_Op_r[2] ),
    .B(_0821_),
    .C(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ),
    .X(_0839_));
 sky130_fd_sc_hd__a211o_1 _3765_ (.A1(net148),
    .A2(\z80.tv80s.i_tv80_core.F[0] ),
    .B1(net96),
    .C1(net153),
    .X(_0840_));
 sky130_fd_sc_hd__a21oi_1 _3766_ (.A1(net162),
    .A2(_2898_),
    .B1(_0840_),
    .Y(_0841_));
 sky130_fd_sc_hd__a21o_1 _3767_ (.A1(net154),
    .A2(_2865_),
    .B1(_0841_),
    .X(_0842_));
 sky130_fd_sc_hd__inv_2 _3768_ (.A(_0842_),
    .Y(_0843_));
 sky130_fd_sc_hd__and3b_4 _3769_ (.A_N(_0821_),
    .B(_0826_),
    .C(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ),
    .X(_0844_));
 sky130_fd_sc_hd__inv_2 _3770_ (.A(_0844_),
    .Y(_0845_));
 sky130_fd_sc_hd__mux2_1 _3771_ (.A0(\z80.tv80s.i_tv80_core.BusB[0] ),
    .A1(\z80.tv80s.i_tv80_core.BusB[4] ),
    .S(\z80.tv80s.i_tv80_core.ALU_Op_r[0] ),
    .X(_0846_));
 sky130_fd_sc_hd__nand2_1 _3772_ (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[2] ),
    .B(_0821_),
    .Y(_0847_));
 sky130_fd_sc_hd__nor2_2 _3773_ (.A(_2862_),
    .B(_0847_),
    .Y(_0848_));
 sky130_fd_sc_hd__or2_1 _3774_ (.A(_2862_),
    .B(_0847_),
    .X(_0849_));
 sky130_fd_sc_hd__a22o_1 _3775_ (.A1(_0844_),
    .A2(_0846_),
    .B1(_0848_),
    .B2(\z80.tv80s.i_tv80_core.BusA[0] ),
    .X(_0850_));
 sky130_fd_sc_hd__and4b_4 _3776_ (.A_N(\z80.tv80s.i_tv80_core.ALU_Op_r[2] ),
    .B(\z80.tv80s.i_tv80_core.ALU_Op_r[0] ),
    .C(net111),
    .D(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ),
    .X(_0851_));
 sky130_fd_sc_hd__a21o_1 _3777_ (.A1(\z80.tv80s.i_tv80_core.BusB[0] ),
    .A2(_0851_),
    .B1(_0834_),
    .X(_0852_));
 sky130_fd_sc_hd__a221o_1 _3778_ (.A1(_0839_),
    .A2(_0843_),
    .B1(_0852_),
    .B2(_0835_),
    .C1(_0850_),
    .X(_0853_));
 sky130_fd_sc_hd__a2111o_1 _3779_ (.A1(_0814_),
    .A2(_0831_),
    .B1(_0838_),
    .C1(_0853_),
    .D1(_2861_),
    .X(_0854_));
 sky130_fd_sc_hd__o211a_1 _3780_ (.A1(\z80.tv80s.i_tv80_core.Save_ALU_r ),
    .A2(\z80.tv80s.di_reg[0] ),
    .B1(_0812_),
    .C1(_0854_),
    .X(_0855_));
 sky130_fd_sc_hd__a21oi_4 _3781_ (.A1(net709),
    .A2(_0811_),
    .B1(_0855_),
    .Y(_0856_));
 sky130_fd_sc_hd__inv_2 _3782_ (.A(_0856_),
    .Y(_0857_));
 sky130_fd_sc_hd__o21ai_1 _3783_ (.A1(_0809_),
    .A2(_0856_),
    .B1(_0775_),
    .Y(_0858_));
 sky130_fd_sc_hd__nand2_1 _3784_ (.A(net152),
    .B(_0412_),
    .Y(_0859_));
 sky130_fd_sc_hd__or3_1 _3785_ (.A(\z80.tv80s.i_tv80_core.i_mcode.MCycle[3] ),
    .B(_2857_),
    .C(_0398_),
    .X(_0860_));
 sky130_fd_sc_hd__nor2_1 _3786_ (.A(net133),
    .B(_0860_),
    .Y(_0861_));
 sky130_fd_sc_hd__o21ai_1 _3787_ (.A1(_2945_),
    .A2(_0861_),
    .B1(net165),
    .Y(_0862_));
 sky130_fd_sc_hd__a31oi_4 _3788_ (.A1(_0747_),
    .A2(_0750_),
    .A3(_0859_),
    .B1(_0862_),
    .Y(_0863_));
 sky130_fd_sc_hd__a211o_1 _3789_ (.A1(_3041_),
    .A2(_0400_),
    .B1(_0767_),
    .C1(_3048_),
    .X(_0864_));
 sky130_fd_sc_hd__a21o_1 _3790_ (.A1(net152),
    .A2(_0398_),
    .B1(net136),
    .X(_0865_));
 sky130_fd_sc_hd__a31o_1 _3791_ (.A1(net106),
    .A2(_0864_),
    .A3(_0865_),
    .B1(_0863_),
    .X(_0866_));
 sky130_fd_sc_hd__inv_2 _3792_ (.A(net81),
    .Y(_0867_));
 sky130_fd_sc_hd__and3_4 _3793_ (.A(_0795_),
    .B(net71),
    .C(net70),
    .X(_0868_));
 sky130_fd_sc_hd__or3_1 _3794_ (.A(_0794_),
    .B(_0799_),
    .C(net69),
    .X(_0869_));
 sky130_fd_sc_hd__and3_4 _3795_ (.A(_0795_),
    .B(net71),
    .C(net69),
    .X(_0870_));
 sky130_fd_sc_hd__or3_1 _3796_ (.A(_0794_),
    .B(_0799_),
    .C(net70),
    .X(_0871_));
 sky130_fd_sc_hd__o22a_1 _3797_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][0] ),
    .A2(_0869_),
    .B1(_0871_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][0] ),
    .X(_0872_));
 sky130_fd_sc_hd__o211a_2 _3798_ (.A1(_0789_),
    .A2(_0792_),
    .B1(_0793_),
    .C1(_0798_),
    .X(_0873_));
 sky130_fd_sc_hd__and2_2 _3799_ (.A(net70),
    .B(_0873_),
    .X(_0874_));
 sky130_fd_sc_hd__nand2_2 _3800_ (.A(net70),
    .B(_0873_),
    .Y(_0875_));
 sky130_fd_sc_hd__and2_2 _3801_ (.A(net69),
    .B(_0873_),
    .X(_0876_));
 sky130_fd_sc_hd__nand2_2 _3802_ (.A(net69),
    .B(_0873_),
    .Y(_0877_));
 sky130_fd_sc_hd__o221a_1 _3803_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][0] ),
    .A2(_0875_),
    .B1(_0877_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][0] ),
    .C1(_0872_),
    .X(_0878_));
 sky130_fd_sc_hd__and3_4 _3804_ (.A(_0795_),
    .B(_0799_),
    .C(net70),
    .X(_0879_));
 sky130_fd_sc_hd__or3_1 _3805_ (.A(_0794_),
    .B(net71),
    .C(net69),
    .X(_0880_));
 sky130_fd_sc_hd__nor2_1 _3806_ (.A(_0795_),
    .B(net71),
    .Y(_0881_));
 sky130_fd_sc_hd__and3_4 _3807_ (.A(_0794_),
    .B(_0799_),
    .C(net70),
    .X(_0882_));
 sky130_fd_sc_hd__nand2_2 _3808_ (.A(net70),
    .B(_0881_),
    .Y(_0883_));
 sky130_fd_sc_hd__o22a_1 _3809_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][0] ),
    .A2(_0880_),
    .B1(_0883_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][0] ),
    .X(_0884_));
 sky130_fd_sc_hd__and3_4 _3810_ (.A(_0794_),
    .B(_0799_),
    .C(net69),
    .X(_0885_));
 sky130_fd_sc_hd__nand2_2 _3811_ (.A(net69),
    .B(_0881_),
    .Y(_0886_));
 sky130_fd_sc_hd__o221a_1 _3812_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][0] ),
    .A2(_0807_),
    .B1(_0886_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][0] ),
    .C1(_0884_),
    .X(_0887_));
 sky130_fd_sc_hd__nand2_2 _3813_ (.A(_0878_),
    .B(_0887_),
    .Y(_0888_));
 sky130_fd_sc_hd__inv_2 _3814_ (.A(_0888_),
    .Y(_0889_));
 sky130_fd_sc_hd__xnor2_1 _3815_ (.A(_0867_),
    .B(_0888_),
    .Y(_0890_));
 sky130_fd_sc_hd__and4_1 _3816_ (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][7] ),
    .B(_0795_),
    .C(net71),
    .D(net69),
    .X(_0891_));
 sky130_fd_sc_hd__and3_1 _3817_ (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][7] ),
    .B(net70),
    .C(_0873_),
    .X(_0892_));
 sky130_fd_sc_hd__and3_1 _3818_ (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][7] ),
    .B(net69),
    .C(_0873_),
    .X(_0893_));
 sky130_fd_sc_hd__a2111o_1 _3819_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][7] ),
    .A2(_0868_),
    .B1(_0891_),
    .C1(_0892_),
    .D1(_0893_),
    .X(_0894_));
 sky130_fd_sc_hd__a22o_1 _3820_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][7] ),
    .A2(_0879_),
    .B1(_0882_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][7] ),
    .X(_0895_));
 sky130_fd_sc_hd__a22o_1 _3821_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][7] ),
    .A2(_0806_),
    .B1(_0885_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][7] ),
    .X(_0896_));
 sky130_fd_sc_hd__or3_2 _3822_ (.A(_0894_),
    .B(_0895_),
    .C(_0896_),
    .X(_0897_));
 sky130_fd_sc_hd__xnor2_1 _3823_ (.A(_0867_),
    .B(_0897_),
    .Y(_0898_));
 sky130_fd_sc_hd__a22o_1 _3824_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][6] ),
    .A2(_0868_),
    .B1(_0870_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][6] ),
    .X(_0899_));
 sky130_fd_sc_hd__mux2_1 _3825_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][6] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][6] ),
    .S(net69),
    .X(_0900_));
 sky130_fd_sc_hd__mux2_1 _3826_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][6] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][6] ),
    .S(net69),
    .X(_0901_));
 sky130_fd_sc_hd__o21a_1 _3827_ (.A1(net71),
    .A2(_0901_),
    .B1(_0794_),
    .X(_0902_));
 sky130_fd_sc_hd__o21a_1 _3828_ (.A1(_0799_),
    .A2(_0900_),
    .B1(_0902_),
    .X(_0903_));
 sky130_fd_sc_hd__a22o_1 _3829_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][6] ),
    .A2(_0806_),
    .B1(_0879_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][6] ),
    .X(_0904_));
 sky130_fd_sc_hd__or3_2 _3830_ (.A(_0899_),
    .B(_0903_),
    .C(_0904_),
    .X(_0905_));
 sky130_fd_sc_hd__and2_1 _3831_ (.A(net80),
    .B(_0905_),
    .X(_0906_));
 sky130_fd_sc_hd__xnor2_1 _3832_ (.A(_0867_),
    .B(_0905_),
    .Y(_0907_));
 sky130_fd_sc_hd__and2_1 _3833_ (.A(_0898_),
    .B(_0907_),
    .X(_0908_));
 sky130_fd_sc_hd__a22o_1 _3834_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][5] ),
    .A2(_0874_),
    .B1(_0876_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][5] ),
    .X(_0909_));
 sky130_fd_sc_hd__a22o_1 _3835_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][5] ),
    .A2(_0868_),
    .B1(_0870_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][5] ),
    .X(_0910_));
 sky130_fd_sc_hd__a22o_1 _3836_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][5] ),
    .A2(_0879_),
    .B1(_0882_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][5] ),
    .X(_0911_));
 sky130_fd_sc_hd__a221o_1 _3837_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][5] ),
    .A2(_0806_),
    .B1(_0885_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][5] ),
    .C1(_0911_),
    .X(_0912_));
 sky130_fd_sc_hd__or3_2 _3838_ (.A(_0909_),
    .B(_0910_),
    .C(_0912_),
    .X(_0913_));
 sky130_fd_sc_hd__xnor2_1 _3839_ (.A(_0867_),
    .B(_0913_),
    .Y(_0914_));
 sky130_fd_sc_hd__a22o_1 _3840_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][4] ),
    .A2(_0868_),
    .B1(_0870_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][4] ),
    .X(_0915_));
 sky130_fd_sc_hd__mux2_1 _3841_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][4] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][4] ),
    .S(net69),
    .X(_0916_));
 sky130_fd_sc_hd__mux2_1 _3842_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][4] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][4] ),
    .S(net69),
    .X(_0917_));
 sky130_fd_sc_hd__o21a_1 _3843_ (.A1(net71),
    .A2(_0917_),
    .B1(_0794_),
    .X(_0918_));
 sky130_fd_sc_hd__o21a_1 _3844_ (.A1(_0799_),
    .A2(_0916_),
    .B1(_0918_),
    .X(_0919_));
 sky130_fd_sc_hd__a22o_1 _3845_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][4] ),
    .A2(_0806_),
    .B1(_0879_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][4] ),
    .X(_0920_));
 sky130_fd_sc_hd__or3_4 _3846_ (.A(_0915_),
    .B(_0919_),
    .C(_0920_),
    .X(_0921_));
 sky130_fd_sc_hd__xnor2_1 _3847_ (.A(_0867_),
    .B(_0921_),
    .Y(_0922_));
 sky130_fd_sc_hd__o311a_1 _3848_ (.A1(_0787_),
    .A2(_0790_),
    .A3(_0800_),
    .B1(_0803_),
    .C1(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][3] ),
    .X(_0923_));
 sky130_fd_sc_hd__a211o_1 _3849_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][3] ),
    .A2(net70),
    .B1(_0923_),
    .C1(_0799_),
    .X(_0924_));
 sky130_fd_sc_hd__o311a_1 _3850_ (.A1(_0787_),
    .A2(_0790_),
    .A3(_0800_),
    .B1(_0803_),
    .C1(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][3] ),
    .X(_0925_));
 sky130_fd_sc_hd__a211o_1 _3851_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][3] ),
    .A2(net70),
    .B1(_0925_),
    .C1(net71),
    .X(_0926_));
 sky130_fd_sc_hd__and3_1 _3852_ (.A(_0794_),
    .B(_0924_),
    .C(_0926_),
    .X(_0927_));
 sky130_fd_sc_hd__mux2_1 _3853_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][3] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][3] ),
    .S(_0805_),
    .X(_0928_));
 sky130_fd_sc_hd__mux2_1 _3854_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][3] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][3] ),
    .S(_0805_),
    .X(_0929_));
 sky130_fd_sc_hd__mux2_1 _3855_ (.A0(_0928_),
    .A1(_0929_),
    .S(_0799_),
    .X(_0930_));
 sky130_fd_sc_hd__a21o_1 _3856_ (.A1(_0795_),
    .A2(_0930_),
    .B1(_0927_),
    .X(_0931_));
 sky130_fd_sc_hd__and2_1 _3857_ (.A(net81),
    .B(_0931_),
    .X(_0932_));
 sky130_fd_sc_hd__nand2_1 _3858_ (.A(net81),
    .B(_0931_),
    .Y(_0933_));
 sky130_fd_sc_hd__nor2_1 _3859_ (.A(net81),
    .B(_0931_),
    .Y(_0934_));
 sky130_fd_sc_hd__mux2_1 _3860_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][2] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][2] ),
    .S(_0805_),
    .X(_0935_));
 sky130_fd_sc_hd__mux2_1 _3861_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][2] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][2] ),
    .S(_0805_),
    .X(_0936_));
 sky130_fd_sc_hd__mux2_1 _3862_ (.A0(_0935_),
    .A1(_0936_),
    .S(_0799_),
    .X(_0937_));
 sky130_fd_sc_hd__mux2_1 _3863_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][2] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][2] ),
    .S(net69),
    .X(_0938_));
 sky130_fd_sc_hd__nor2_1 _3864_ (.A(_0799_),
    .B(_0938_),
    .Y(_0939_));
 sky130_fd_sc_hd__mux2_1 _3865_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][2] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][2] ),
    .S(net69),
    .X(_0940_));
 sky130_fd_sc_hd__o21ai_1 _3866_ (.A1(net71),
    .A2(_0940_),
    .B1(_0794_),
    .Y(_0941_));
 sky130_fd_sc_hd__a2bb2o_2 _3867_ (.A1_N(_0939_),
    .A2_N(_0941_),
    .B1(_0795_),
    .B2(_0937_),
    .X(_0942_));
 sky130_fd_sc_hd__nand2_1 _3868_ (.A(net81),
    .B(_0942_),
    .Y(_0943_));
 sky130_fd_sc_hd__mux2_1 _3869_ (.A0(net379),
    .A1(net391),
    .S(net70),
    .X(_0944_));
 sky130_fd_sc_hd__a311o_1 _3870_ (.A1(_0788_),
    .A2(_0791_),
    .A3(_0801_),
    .B1(_0802_),
    .C1(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][1] ),
    .X(_0945_));
 sky130_fd_sc_hd__o211a_1 _3871_ (.A1(net486),
    .A2(_0805_),
    .B1(_0945_),
    .C1(_0799_),
    .X(_0946_));
 sky130_fd_sc_hd__a211o_1 _3872_ (.A1(_0798_),
    .A2(_0944_),
    .B1(_0946_),
    .C1(_0794_),
    .X(_0947_));
 sky130_fd_sc_hd__a311o_1 _3873_ (.A1(_0788_),
    .A2(_0791_),
    .A3(_0801_),
    .B1(_0802_),
    .C1(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][1] ),
    .X(_0948_));
 sky130_fd_sc_hd__mux2_1 _3874_ (.A0(net299),
    .A1(net283),
    .S(net70),
    .X(_0949_));
 sky130_fd_sc_hd__o211a_1 _3875_ (.A1(net303),
    .A2(_0805_),
    .B1(_0948_),
    .C1(_0798_),
    .X(_0950_));
 sky130_fd_sc_hd__a211o_1 _3876_ (.A1(_0799_),
    .A2(_0949_),
    .B1(_0950_),
    .C1(_0795_),
    .X(_0951_));
 sky130_fd_sc_hd__nand2_1 _3877_ (.A(_0947_),
    .B(_0951_),
    .Y(_0952_));
 sky130_fd_sc_hd__and3_1 _3878_ (.A(net81),
    .B(_0947_),
    .C(_0951_),
    .X(_0953_));
 sky130_fd_sc_hd__a21o_1 _3879_ (.A1(_0947_),
    .A2(_0951_),
    .B1(net81),
    .X(_0954_));
 sky130_fd_sc_hd__nand2b_1 _3880_ (.A_N(_0953_),
    .B(_0954_),
    .Y(_0955_));
 sky130_fd_sc_hd__mux2_1 _3881_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][0] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][0] ),
    .S(net70),
    .X(_0956_));
 sky130_fd_sc_hd__mux2_1 _3882_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][0] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][0] ),
    .S(net70),
    .X(_0957_));
 sky130_fd_sc_hd__mux2_1 _3883_ (.A0(_0956_),
    .A1(_0957_),
    .S(_0799_),
    .X(_0958_));
 sky130_fd_sc_hd__mux2_1 _3884_ (.A0(net346),
    .A1(net295),
    .S(net70),
    .X(_0959_));
 sky130_fd_sc_hd__nand2_1 _3885_ (.A(net71),
    .B(_0959_),
    .Y(_0960_));
 sky130_fd_sc_hd__mux2_1 _3886_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][0] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][0] ),
    .S(_0804_),
    .X(_0961_));
 sky130_fd_sc_hd__a21oi_1 _3887_ (.A1(_0799_),
    .A2(_0961_),
    .B1(_0794_),
    .Y(_0962_));
 sky130_fd_sc_hd__o2bb2a_2 _3888_ (.A1_N(_0960_),
    .A2_N(_0962_),
    .B1(_0795_),
    .B2(_0958_),
    .X(_0963_));
 sky130_fd_sc_hd__a2bb2o_1 _3889_ (.A1_N(_0795_),
    .A2_N(_0958_),
    .B1(_0960_),
    .B2(_0962_),
    .X(_0964_));
 sky130_fd_sc_hd__a21oi_1 _3890_ (.A1(_0954_),
    .A2(_0963_),
    .B1(_0953_),
    .Y(_0965_));
 sky130_fd_sc_hd__nor2_1 _3891_ (.A(net81),
    .B(_0942_),
    .Y(_0966_));
 sky130_fd_sc_hd__xnor2_1 _3892_ (.A(net81),
    .B(_0942_),
    .Y(_0967_));
 sky130_fd_sc_hd__or2_1 _3893_ (.A(_0965_),
    .B(_0967_),
    .X(_0968_));
 sky130_fd_sc_hd__nand2_1 _3894_ (.A(_0943_),
    .B(_0968_),
    .Y(_0969_));
 sky130_fd_sc_hd__o311a_1 _3895_ (.A1(_0934_),
    .A2(_0965_),
    .A3(_0967_),
    .B1(_0943_),
    .C1(_0933_),
    .X(_0970_));
 sky130_fd_sc_hd__and2b_1 _3896_ (.A_N(_0970_),
    .B(_0922_),
    .X(_0971_));
 sky130_fd_sc_hd__and2_1 _3897_ (.A(_0914_),
    .B(_0971_),
    .X(_0972_));
 sky130_fd_sc_hd__and3_1 _3898_ (.A(_0908_),
    .B(_0914_),
    .C(_0971_),
    .X(_0973_));
 sky130_fd_sc_hd__o21a_1 _3899_ (.A1(_0913_),
    .A2(_0921_),
    .B1(net80),
    .X(_0974_));
 sky130_fd_sc_hd__a221o_1 _3900_ (.A1(net80),
    .A2(_0897_),
    .B1(_0908_),
    .B2(_0974_),
    .C1(_0906_),
    .X(_0975_));
 sky130_fd_sc_hd__or2_1 _3901_ (.A(_0973_),
    .B(_0975_),
    .X(_0976_));
 sky130_fd_sc_hd__o21bai_2 _3902_ (.A1(_0973_),
    .A2(_0975_),
    .B1_N(_0890_),
    .Y(_0977_));
 sky130_fd_sc_hd__xnor2_1 _3903_ (.A(_0890_),
    .B(_0976_),
    .Y(_0978_));
 sky130_fd_sc_hd__a21o_1 _3904_ (.A1(net76),
    .A2(_0978_),
    .B1(_0858_),
    .X(_0979_));
 sky130_fd_sc_hd__o21a_1 _3905_ (.A1(net229),
    .A2(net85),
    .B1(net86),
    .X(_0980_));
 sky130_fd_sc_hd__nor2_4 _3906_ (.A(\z80.tv80s.i_tv80_core.RegAddrB_r[0] ),
    .B(net89),
    .Y(_0981_));
 sky130_fd_sc_hd__or2_1 _3907_ (.A(\z80.tv80s.i_tv80_core.Alternate ),
    .B(net86),
    .X(_0982_));
 sky130_fd_sc_hd__o21a_1 _3908_ (.A1(\z80.tv80s.i_tv80_core.RegAddrB_r[2] ),
    .A2(_0772_),
    .B1(_0982_),
    .X(_0983_));
 sky130_fd_sc_hd__o21ai_4 _3909_ (.A1(\z80.tv80s.i_tv80_core.RegAddrB_r[2] ),
    .A2(_0772_),
    .B1(_0982_),
    .Y(_0984_));
 sky130_fd_sc_hd__mux4_2 _3910_ (.A0(net496),
    .A1(net440),
    .A2(net383),
    .A3(net329),
    .S0(net83),
    .S1(net74),
    .X(_0985_));
 sky130_fd_sc_hd__a22o_2 _3911_ (.A1(_0979_),
    .A2(_0980_),
    .B1(_0985_),
    .B2(net89),
    .X(_0986_));
 sky130_fd_sc_hd__mux2_1 _3912_ (.A0(_0986_),
    .A1(net457),
    .S(_0808_),
    .X(_0040_));
 sky130_fd_sc_hd__and2b_1 _3913_ (.A_N(\z80.tv80s.i_tv80_core.BusB[1] ),
    .B(net143),
    .X(_0987_));
 sky130_fd_sc_hd__and2b_1 _3914_ (.A_N(net143),
    .B(\z80.tv80s.i_tv80_core.BusB[1] ),
    .X(_0988_));
 sky130_fd_sc_hd__o21ai_1 _3915_ (.A1(_0987_),
    .A2(_0988_),
    .B1(\z80.tv80s.i_tv80_core.BusA[1] ),
    .Y(_0989_));
 sky130_fd_sc_hd__nand2_1 _3916_ (.A(net111),
    .B(_0989_),
    .Y(_0990_));
 sky130_fd_sc_hd__or3_1 _3917_ (.A(\z80.tv80s.i_tv80_core.BusA[1] ),
    .B(_0987_),
    .C(_0988_),
    .X(_0991_));
 sky130_fd_sc_hd__and2_1 _3918_ (.A(_0989_),
    .B(_0991_),
    .X(_0992_));
 sky130_fd_sc_hd__a21o_1 _3919_ (.A1(_0819_),
    .A2(_0823_),
    .B1(_0817_),
    .X(_0993_));
 sky130_fd_sc_hd__or2_1 _3920_ (.A(_0992_),
    .B(_0993_),
    .X(_0994_));
 sky130_fd_sc_hd__nand2_1 _3921_ (.A(_0992_),
    .B(_0993_),
    .Y(_0995_));
 sky130_fd_sc_hd__a22o_1 _3922_ (.A1(_0815_),
    .A2(_0990_),
    .B1(_0992_),
    .B2(_0828_),
    .X(_0996_));
 sky130_fd_sc_hd__a31o_1 _3923_ (.A1(_0827_),
    .A2(_0994_),
    .A3(_0995_),
    .B1(_0996_),
    .X(_0997_));
 sky130_fd_sc_hd__o41a_2 _3924_ (.A1(net111),
    .A2(\z80.tv80s.i_tv80_core.BusA[1] ),
    .A3(\z80.tv80s.i_tv80_core.BusB[1] ),
    .A4(_0827_),
    .B1(_0997_),
    .X(_0998_));
 sky130_fd_sc_hd__mux2_1 _3925_ (.A0(\z80.tv80s.i_tv80_core.BusB[1] ),
    .A1(\z80.tv80s.i_tv80_core.BusB[5] ),
    .S(\z80.tv80s.i_tv80_core.ALU_Op_r[0] ),
    .X(_0999_));
 sky130_fd_sc_hd__mux2_1 _3926_ (.A0(\z80.tv80s.i_tv80_core.BusA[0] ),
    .A1(\z80.tv80s.i_tv80_core.BusA[2] ),
    .S(net153),
    .X(_1000_));
 sky130_fd_sc_hd__nor2_1 _3927_ (.A(net144),
    .B(_0469_),
    .Y(_1001_));
 sky130_fd_sc_hd__nor2_1 _3928_ (.A(_2867_),
    .B(_0833_),
    .Y(_1002_));
 sky130_fd_sc_hd__o31a_1 _3929_ (.A1(net144),
    .A2(_0469_),
    .A3(_0851_),
    .B1(\z80.tv80s.i_tv80_core.BusB[1] ),
    .X(_1003_));
 sky130_fd_sc_hd__o22a_1 _3930_ (.A1(_1001_),
    .A2(_1002_),
    .B1(_1003_),
    .B2(_0834_),
    .X(_1004_));
 sky130_fd_sc_hd__a221o_1 _3931_ (.A1(_0844_),
    .A2(_0999_),
    .B1(_1000_),
    .B2(_0839_),
    .C1(_1004_),
    .X(_1005_));
 sky130_fd_sc_hd__o21a_1 _3932_ (.A1(\z80.tv80s.i_tv80_core.BusA[1] ),
    .A2(\z80.tv80s.i_tv80_core.BusA[2] ),
    .B1(\z80.tv80s.i_tv80_core.BusA[3] ),
    .X(_1006_));
 sky130_fd_sc_hd__o21ai_1 _3933_ (.A1(\z80.tv80s.i_tv80_core.BusA[1] ),
    .A2(\z80.tv80s.i_tv80_core.BusA[2] ),
    .B1(\z80.tv80s.i_tv80_core.BusA[3] ),
    .Y(_1007_));
 sky130_fd_sc_hd__nor2_1 _3934_ (.A(\z80.tv80s.i_tv80_core.F[4] ),
    .B(_1006_),
    .Y(_1008_));
 sky130_fd_sc_hd__or2_1 _3935_ (.A(\z80.tv80s.i_tv80_core.BusA[3] ),
    .B(\z80.tv80s.i_tv80_core.F[4] ),
    .X(_1009_));
 sky130_fd_sc_hd__mux2_1 _3936_ (.A0(_1008_),
    .A1(_1009_),
    .S(\z80.tv80s.i_tv80_core.BusA[1] ),
    .X(_1010_));
 sky130_fd_sc_hd__a2bb2o_1 _3937_ (.A1_N(_0849_),
    .A2_N(_1010_),
    .B1(_0998_),
    .B2(_0814_),
    .X(_1011_));
 sky130_fd_sc_hd__nor2_1 _3938_ (.A(_1005_),
    .B(_1011_),
    .Y(_1012_));
 sky130_fd_sc_hd__mux2_1 _3939_ (.A0(_2871_),
    .A1(_1012_),
    .S(\z80.tv80s.i_tv80_core.Save_ALU_r ),
    .X(_1013_));
 sky130_fd_sc_hd__mux2_4 _3940_ (.A0(_2867_),
    .A1(_1013_),
    .S(_0812_),
    .X(_1014_));
 sky130_fd_sc_hd__inv_2 _3941_ (.A(_1014_),
    .Y(_1015_));
 sky130_fd_sc_hd__o21ai_1 _3942_ (.A1(_0809_),
    .A2(_1014_),
    .B1(_0775_),
    .Y(_1016_));
 sky130_fd_sc_hd__a22o_1 _3943_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][1] ),
    .A2(_0874_),
    .B1(_0876_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][1] ),
    .X(_1017_));
 sky130_fd_sc_hd__a22o_1 _3944_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][1] ),
    .A2(_0868_),
    .B1(_0870_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][1] ),
    .X(_1018_));
 sky130_fd_sc_hd__a22o_1 _3945_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][1] ),
    .A2(_0879_),
    .B1(_0882_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][1] ),
    .X(_1019_));
 sky130_fd_sc_hd__a221o_1 _3946_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][1] ),
    .A2(_0806_),
    .B1(_0885_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][1] ),
    .C1(_1019_),
    .X(_1020_));
 sky130_fd_sc_hd__or3_4 _3947_ (.A(_1017_),
    .B(_1018_),
    .C(_1020_),
    .X(_1021_));
 sky130_fd_sc_hd__xnor2_1 _3948_ (.A(net80),
    .B(_1021_),
    .Y(_1022_));
 sky130_fd_sc_hd__o21ai_1 _3949_ (.A1(_0867_),
    .A2(_0888_),
    .B1(_0977_),
    .Y(_1023_));
 sky130_fd_sc_hd__xnor2_1 _3950_ (.A(_1022_),
    .B(_1023_),
    .Y(_1024_));
 sky130_fd_sc_hd__a21o_1 _3951_ (.A1(net76),
    .A2(_1024_),
    .B1(_1016_),
    .X(_1025_));
 sky130_fd_sc_hd__o21a_1 _3952_ (.A1(net243),
    .A2(net85),
    .B1(net86),
    .X(_1026_));
 sky130_fd_sc_hd__mux4_1 _3953_ (.A0(net446),
    .A1(net311),
    .A2(net459),
    .A3(net381),
    .S0(net74),
    .S1(net83),
    .X(_1027_));
 sky130_fd_sc_hd__a22o_2 _3954_ (.A1(_1025_),
    .A2(_1026_),
    .B1(_1027_),
    .B2(net89),
    .X(_1028_));
 sky130_fd_sc_hd__mux2_1 _3955_ (.A0(_1028_),
    .A1(net452),
    .S(_0808_),
    .X(_0041_));
 sky130_fd_sc_hd__mux4_1 _3956_ (.A0(net361),
    .A1(net315),
    .A2(net427),
    .A3(net313),
    .S0(net74),
    .S1(net83),
    .X(_1029_));
 sky130_fd_sc_hd__a22o_1 _3957_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][2] ),
    .A2(_0874_),
    .B1(_0876_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][2] ),
    .X(_1030_));
 sky130_fd_sc_hd__a221o_1 _3958_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][2] ),
    .A2(_0868_),
    .B1(_0870_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][2] ),
    .C1(_1030_),
    .X(_1031_));
 sky130_fd_sc_hd__a22o_1 _3959_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][2] ),
    .A2(_0879_),
    .B1(_0882_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][2] ),
    .X(_1032_));
 sky130_fd_sc_hd__a221o_1 _3960_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][2] ),
    .A2(_0806_),
    .B1(_0885_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][2] ),
    .C1(_1032_),
    .X(_1033_));
 sky130_fd_sc_hd__or2_2 _3961_ (.A(_1031_),
    .B(_1033_),
    .X(_1034_));
 sky130_fd_sc_hd__xnor2_1 _3962_ (.A(net80),
    .B(_1034_),
    .Y(_1035_));
 sky130_fd_sc_hd__o21ai_1 _3963_ (.A1(_0889_),
    .A2(_1021_),
    .B1(net80),
    .Y(_1036_));
 sky130_fd_sc_hd__o21bai_1 _3964_ (.A1(net80),
    .A2(_1021_),
    .B1_N(_0977_),
    .Y(_1037_));
 sky130_fd_sc_hd__a21oi_1 _3965_ (.A1(_1036_),
    .A2(_1037_),
    .B1(_1035_),
    .Y(_1038_));
 sky130_fd_sc_hd__and3_1 _3966_ (.A(_1035_),
    .B(_1036_),
    .C(_1037_),
    .X(_1039_));
 sky130_fd_sc_hd__nor2_1 _3967_ (.A(_1038_),
    .B(_1039_),
    .Y(_1040_));
 sky130_fd_sc_hd__nor2_1 _3968_ (.A(net111),
    .B(\z80.tv80s.i_tv80_core.BusB[2] ),
    .Y(_1041_));
 sky130_fd_sc_hd__nor2_1 _3969_ (.A(net143),
    .B(_2868_),
    .Y(_1042_));
 sky130_fd_sc_hd__o21ai_1 _3970_ (.A1(_1041_),
    .A2(_1042_),
    .B1(\z80.tv80s.i_tv80_core.BusA[2] ),
    .Y(_1043_));
 sky130_fd_sc_hd__nand2_1 _3971_ (.A(net111),
    .B(_1043_),
    .Y(_1044_));
 sky130_fd_sc_hd__or3_1 _3972_ (.A(\z80.tv80s.i_tv80_core.BusA[2] ),
    .B(_1041_),
    .C(_1042_),
    .X(_1045_));
 sky130_fd_sc_hd__and2_1 _3973_ (.A(_1043_),
    .B(_1045_),
    .X(_1046_));
 sky130_fd_sc_hd__nand2_1 _3974_ (.A(_0989_),
    .B(_0995_),
    .Y(_1047_));
 sky130_fd_sc_hd__xnor2_1 _3975_ (.A(_1046_),
    .B(_1047_),
    .Y(_1048_));
 sky130_fd_sc_hd__a22o_1 _3976_ (.A1(_0815_),
    .A2(_1044_),
    .B1(_1046_),
    .B2(_0828_),
    .X(_1049_));
 sky130_fd_sc_hd__o21ba_1 _3977_ (.A1(_0826_),
    .A2(_1048_),
    .B1_N(_1049_),
    .X(_1050_));
 sky130_fd_sc_hd__a31o_1 _3978_ (.A1(_2866_),
    .A2(_0826_),
    .A3(_1041_),
    .B1(_1050_),
    .X(_1051_));
 sky130_fd_sc_hd__nand2_1 _3979_ (.A(_0814_),
    .B(_1051_),
    .Y(_1052_));
 sky130_fd_sc_hd__mux2_1 _3980_ (.A0(\z80.tv80s.i_tv80_core.F[1] ),
    .A1(_2865_),
    .S(_1008_),
    .X(_1053_));
 sky130_fd_sc_hd__xor2_1 _3981_ (.A(\z80.tv80s.i_tv80_core.BusA[1] ),
    .B(\z80.tv80s.i_tv80_core.BusA[2] ),
    .X(_1054_));
 sky130_fd_sc_hd__xnor2_2 _3982_ (.A(_1053_),
    .B(_1054_),
    .Y(_1055_));
 sky130_fd_sc_hd__mux2_1 _3983_ (.A0(\z80.tv80s.i_tv80_core.BusB[2] ),
    .A1(\z80.tv80s.i_tv80_core.BusB[6] ),
    .S(\z80.tv80s.i_tv80_core.ALU_Op_r[0] ),
    .X(_1056_));
 sky130_fd_sc_hd__mux2_1 _3984_ (.A0(\z80.tv80s.i_tv80_core.BusA[1] ),
    .A1(\z80.tv80s.i_tv80_core.BusA[3] ),
    .S(net154),
    .X(_1057_));
 sky130_fd_sc_hd__a221o_1 _3985_ (.A1(_0844_),
    .A2(_1056_),
    .B1(_1057_),
    .B2(_0839_),
    .C1(_0814_),
    .X(_1058_));
 sky130_fd_sc_hd__nor2_1 _3986_ (.A(net144),
    .B(_3029_),
    .Y(_1059_));
 sky130_fd_sc_hd__nor2_1 _3987_ (.A(_0836_),
    .B(_1059_),
    .Y(_1060_));
 sky130_fd_sc_hd__a211o_1 _3988_ (.A1(_0851_),
    .A2(_1059_),
    .B1(_1060_),
    .C1(_0834_),
    .X(_1061_));
 sky130_fd_sc_hd__a22o_1 _3989_ (.A1(_0848_),
    .A2(_1055_),
    .B1(_1061_),
    .B2(\z80.tv80s.i_tv80_core.BusB[2] ),
    .X(_1062_));
 sky130_fd_sc_hd__a211o_1 _3990_ (.A1(_0834_),
    .A2(_1059_),
    .B1(_1062_),
    .C1(_1058_),
    .X(_1063_));
 sky130_fd_sc_hd__and3_1 _3991_ (.A(\z80.tv80s.i_tv80_core.Save_ALU_r ),
    .B(_1052_),
    .C(_1063_),
    .X(_1064_));
 sky130_fd_sc_hd__a21oi_1 _3992_ (.A1(_2861_),
    .A2(\z80.tv80s.di_reg[2] ),
    .B1(_1064_),
    .Y(_1065_));
 sky130_fd_sc_hd__mux2_4 _3993_ (.A0(_2868_),
    .A1(_1065_),
    .S(_0812_),
    .X(_1066_));
 sky130_fd_sc_hd__inv_2 _3994_ (.A(_1066_),
    .Y(_1067_));
 sky130_fd_sc_hd__o21ai_1 _3995_ (.A1(net76),
    .A2(_1066_),
    .B1(_0775_),
    .Y(_1068_));
 sky130_fd_sc_hd__a21o_1 _3996_ (.A1(_0809_),
    .A2(_1040_),
    .B1(_1068_),
    .X(_1069_));
 sky130_fd_sc_hd__o21a_1 _3997_ (.A1(net237),
    .A2(net85),
    .B1(_1069_),
    .X(_1070_));
 sky130_fd_sc_hd__mux2_2 _3998_ (.A0(_1029_),
    .A1(_1070_),
    .S(net86),
    .X(_1071_));
 sky130_fd_sc_hd__mux2_1 _3999_ (.A0(_1071_),
    .A1(net507),
    .S(_0808_),
    .X(_0042_));
 sky130_fd_sc_hd__nor2_1 _4000_ (.A(net111),
    .B(\z80.tv80s.i_tv80_core.BusB[3] ),
    .Y(_1072_));
 sky130_fd_sc_hd__and2_1 _4001_ (.A(net111),
    .B(\z80.tv80s.i_tv80_core.BusB[3] ),
    .X(_1073_));
 sky130_fd_sc_hd__o21a_1 _4002_ (.A1(_1072_),
    .A2(_1073_),
    .B1(\z80.tv80s.i_tv80_core.BusA[3] ),
    .X(_1074_));
 sky130_fd_sc_hd__or2_1 _4003_ (.A(net143),
    .B(_1074_),
    .X(_1075_));
 sky130_fd_sc_hd__nor3_1 _4004_ (.A(\z80.tv80s.i_tv80_core.BusA[3] ),
    .B(_1072_),
    .C(_1073_),
    .Y(_1076_));
 sky130_fd_sc_hd__nor2_1 _4005_ (.A(_1074_),
    .B(_1076_),
    .Y(_1077_));
 sky130_fd_sc_hd__a21bo_1 _4006_ (.A1(_1046_),
    .A2(_1047_),
    .B1_N(_1043_),
    .X(_1078_));
 sky130_fd_sc_hd__or2_1 _4007_ (.A(_1077_),
    .B(_1078_),
    .X(_1079_));
 sky130_fd_sc_hd__a21oi_1 _4008_ (.A1(_1077_),
    .A2(_1078_),
    .B1(_0826_),
    .Y(_1080_));
 sky130_fd_sc_hd__a22o_1 _4009_ (.A1(_0815_),
    .A2(_1075_),
    .B1(_1077_),
    .B2(_0828_),
    .X(_1081_));
 sky130_fd_sc_hd__a21o_1 _4010_ (.A1(_1079_),
    .A2(_1080_),
    .B1(_1081_),
    .X(_1082_));
 sky130_fd_sc_hd__o41a_2 _4011_ (.A1(_2864_),
    .A2(\z80.tv80s.i_tv80_core.BusA[3] ),
    .A3(\z80.tv80s.i_tv80_core.BusB[3] ),
    .A4(_0827_),
    .B1(_1082_),
    .X(_1083_));
 sky130_fd_sc_hd__a21o_1 _4012_ (.A1(\z80.tv80s.i_tv80_core.BusA[1] ),
    .A2(\z80.tv80s.i_tv80_core.BusA[2] ),
    .B1(\z80.tv80s.i_tv80_core.BusA[3] ),
    .X(_1084_));
 sky130_fd_sc_hd__a31oi_1 _4013_ (.A1(\z80.tv80s.i_tv80_core.BusA[1] ),
    .A2(\z80.tv80s.i_tv80_core.BusA[2] ),
    .A3(\z80.tv80s.i_tv80_core.BusA[3] ),
    .B1(_1008_),
    .Y(_1085_));
 sky130_fd_sc_hd__or3_1 _4014_ (.A(\z80.tv80s.i_tv80_core.BusA[1] ),
    .B(\z80.tv80s.i_tv80_core.BusA[2] ),
    .C(\z80.tv80s.i_tv80_core.BusA[3] ),
    .X(_1086_));
 sky130_fd_sc_hd__a21o_1 _4015_ (.A1(_1007_),
    .A2(_1086_),
    .B1(\z80.tv80s.i_tv80_core.F[1] ),
    .X(_1087_));
 sky130_fd_sc_hd__nand2_1 _4016_ (.A(_1009_),
    .B(_1087_),
    .Y(_1088_));
 sky130_fd_sc_hd__a31o_1 _4017_ (.A1(\z80.tv80s.i_tv80_core.F[1] ),
    .A2(_1084_),
    .A3(_1085_),
    .B1(_1088_),
    .X(_1089_));
 sky130_fd_sc_hd__mux2_1 _4018_ (.A0(\z80.tv80s.i_tv80_core.BusB[3] ),
    .A1(\z80.tv80s.i_tv80_core.BusB[7] ),
    .S(\z80.tv80s.i_tv80_core.ALU_Op_r[0] ),
    .X(_1090_));
 sky130_fd_sc_hd__mux2_1 _4019_ (.A0(\z80.tv80s.i_tv80_core.BusA[2] ),
    .A1(\z80.tv80s.i_tv80_core.BusA[4] ),
    .S(net154),
    .X(_1091_));
 sky130_fd_sc_hd__and2_1 _4020_ (.A(_0839_),
    .B(_1091_),
    .X(_1092_));
 sky130_fd_sc_hd__mux2_1 _4021_ (.A0(_0837_),
    .A1(_0851_),
    .S(_0468_),
    .X(_1093_));
 sky130_fd_sc_hd__or2_1 _4022_ (.A(\z80.tv80s.i_tv80_core.BusB[3] ),
    .B(_0468_),
    .X(_1094_));
 sky130_fd_sc_hd__a2bb2o_1 _4023_ (.A1_N(_0849_),
    .A2_N(_1089_),
    .B1(_1090_),
    .B2(_0844_),
    .X(_1095_));
 sky130_fd_sc_hd__a221o_1 _4024_ (.A1(\z80.tv80s.i_tv80_core.BusB[3] ),
    .A2(_1093_),
    .B1(_1094_),
    .B2(_0834_),
    .C1(_1092_),
    .X(_1096_));
 sky130_fd_sc_hd__a211o_1 _4025_ (.A1(_0814_),
    .A2(_1083_),
    .B1(_1095_),
    .C1(_1096_),
    .X(_1097_));
 sky130_fd_sc_hd__mux2_1 _4026_ (.A0(\z80.tv80s.di_reg[3] ),
    .A1(_1097_),
    .S(\z80.tv80s.i_tv80_core.Save_ALU_r ),
    .X(_1098_));
 sky130_fd_sc_hd__and2_1 _4027_ (.A(net649),
    .B(_0811_),
    .X(_1099_));
 sky130_fd_sc_hd__a21oi_4 _4028_ (.A1(_0812_),
    .A2(_1098_),
    .B1(_1099_),
    .Y(_1100_));
 sky130_fd_sc_hd__inv_2 _4029_ (.A(_1100_),
    .Y(_1101_));
 sky130_fd_sc_hd__o21ai_1 _4030_ (.A1(_0809_),
    .A2(_1100_),
    .B1(_0775_),
    .Y(_1102_));
 sky130_fd_sc_hd__a22o_1 _4031_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][3] ),
    .A2(_0868_),
    .B1(_0870_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][3] ),
    .X(_1103_));
 sky130_fd_sc_hd__a221o_1 _4032_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][3] ),
    .A2(_0874_),
    .B1(_0876_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][3] ),
    .C1(_1103_),
    .X(_1104_));
 sky130_fd_sc_hd__a22o_1 _4033_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][3] ),
    .A2(_0879_),
    .B1(_0882_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][3] ),
    .X(_1105_));
 sky130_fd_sc_hd__a221o_1 _4034_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][3] ),
    .A2(_0806_),
    .B1(_0885_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][3] ),
    .C1(_1105_),
    .X(_1106_));
 sky130_fd_sc_hd__or2_2 _4035_ (.A(_1104_),
    .B(_1106_),
    .X(_1107_));
 sky130_fd_sc_hd__xnor2_1 _4036_ (.A(_0867_),
    .B(_1107_),
    .Y(_1108_));
 sky130_fd_sc_hd__a21o_1 _4037_ (.A1(net80),
    .A2(_1034_),
    .B1(_1038_),
    .X(_1109_));
 sky130_fd_sc_hd__xor2_1 _4038_ (.A(_1108_),
    .B(_1109_),
    .X(_1110_));
 sky130_fd_sc_hd__a21o_1 _4039_ (.A1(net76),
    .A2(_1110_),
    .B1(_1102_),
    .X(_1111_));
 sky130_fd_sc_hd__o21a_1 _4040_ (.A1(net235),
    .A2(net85),
    .B1(net86),
    .X(_1112_));
 sky130_fd_sc_hd__mux4_2 _4041_ (.A0(net367),
    .A1(net393),
    .A2(net385),
    .A3(net293),
    .S0(net74),
    .S1(net82),
    .X(_1113_));
 sky130_fd_sc_hd__a22o_2 _4042_ (.A1(_1111_),
    .A2(_1112_),
    .B1(_1113_),
    .B2(net89),
    .X(_1114_));
 sky130_fd_sc_hd__mux2_1 _4043_ (.A0(_1114_),
    .A1(net505),
    .S(_0808_),
    .X(_0043_));
 sky130_fd_sc_hd__o41a_1 _4044_ (.A1(_0889_),
    .A2(_1021_),
    .A3(_1034_),
    .A4(_1107_),
    .B1(net80),
    .X(_1115_));
 sky130_fd_sc_hd__or3b_1 _4045_ (.A(_1022_),
    .B(_1035_),
    .C_N(_1108_),
    .X(_1116_));
 sky130_fd_sc_hd__o21bai_2 _4046_ (.A1(_0977_),
    .A2(_1116_),
    .B1_N(_1115_),
    .Y(_1117_));
 sky130_fd_sc_hd__a22o_1 _4047_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][4] ),
    .A2(_0868_),
    .B1(_0870_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][4] ),
    .X(_1118_));
 sky130_fd_sc_hd__a221o_1 _4048_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][4] ),
    .A2(_0874_),
    .B1(_0876_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][4] ),
    .C1(_1118_),
    .X(_1119_));
 sky130_fd_sc_hd__a22o_1 _4049_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][4] ),
    .A2(_0879_),
    .B1(_0882_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][4] ),
    .X(_1120_));
 sky130_fd_sc_hd__a221o_1 _4050_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][4] ),
    .A2(_0806_),
    .B1(_0885_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][4] ),
    .C1(_1120_),
    .X(_1121_));
 sky130_fd_sc_hd__or2_2 _4051_ (.A(_1119_),
    .B(_1121_),
    .X(_1122_));
 sky130_fd_sc_hd__xnor2_1 _4052_ (.A(_0867_),
    .B(_1122_),
    .Y(_1123_));
 sky130_fd_sc_hd__xnor2_1 _4053_ (.A(_1117_),
    .B(_1123_),
    .Y(_1124_));
 sky130_fd_sc_hd__nand2_1 _4054_ (.A(\z80.tv80s.i_tv80_core.F[1] ),
    .B(\z80.tv80s.i_tv80_core.F[4] ),
    .Y(_1125_));
 sky130_fd_sc_hd__o22a_1 _4055_ (.A1(\z80.tv80s.i_tv80_core.F[1] ),
    .A2(_1007_),
    .B1(_1084_),
    .B2(_1125_),
    .X(_1126_));
 sky130_fd_sc_hd__xor2_2 _4056_ (.A(\z80.tv80s.i_tv80_core.BusA[4] ),
    .B(_1126_),
    .X(_1127_));
 sky130_fd_sc_hd__nor2_1 _4057_ (.A(_0849_),
    .B(_1127_),
    .Y(_1128_));
 sky130_fd_sc_hd__mux2_1 _4058_ (.A0(\z80.tv80s.i_tv80_core.BusA[3] ),
    .A1(\z80.tv80s.i_tv80_core.BusA[5] ),
    .S(net154),
    .X(_1129_));
 sky130_fd_sc_hd__nor2_1 _4059_ (.A(_2864_),
    .B(\z80.tv80s.i_tv80_core.BusB[4] ),
    .Y(_1130_));
 sky130_fd_sc_hd__or3b_1 _4060_ (.A(\z80.tv80s.i_tv80_core.BusA[4] ),
    .B(_0827_),
    .C_N(_1130_),
    .X(_1131_));
 sky130_fd_sc_hd__and2_1 _4061_ (.A(_2864_),
    .B(\z80.tv80s.i_tv80_core.BusB[4] ),
    .X(_1132_));
 sky130_fd_sc_hd__o21ai_1 _4062_ (.A1(_1130_),
    .A2(_1132_),
    .B1(\z80.tv80s.i_tv80_core.BusA[4] ),
    .Y(_1133_));
 sky130_fd_sc_hd__or3_1 _4063_ (.A(\z80.tv80s.i_tv80_core.BusA[4] ),
    .B(_1130_),
    .C(_1132_),
    .X(_1134_));
 sky130_fd_sc_hd__and2_1 _4064_ (.A(_1133_),
    .B(_1134_),
    .X(_1135_));
 sky130_fd_sc_hd__a21o_1 _4065_ (.A1(_1077_),
    .A2(_1078_),
    .B1(_1074_),
    .X(_1136_));
 sky130_fd_sc_hd__a21oi_1 _4066_ (.A1(_1135_),
    .A2(_1136_),
    .B1(_0826_),
    .Y(_1137_));
 sky130_fd_sc_hd__o21a_1 _4067_ (.A1(_1135_),
    .A2(_1136_),
    .B1(_1137_),
    .X(_1138_));
 sky130_fd_sc_hd__nand2_1 _4068_ (.A(net111),
    .B(_1133_),
    .Y(_1139_));
 sky130_fd_sc_hd__a221o_1 _4069_ (.A1(_0828_),
    .A2(_1135_),
    .B1(_1139_),
    .B2(_0815_),
    .C1(_1138_),
    .X(_1140_));
 sky130_fd_sc_hd__nand2_1 _4070_ (.A(_1131_),
    .B(_1140_),
    .Y(_1141_));
 sky130_fd_sc_hd__inv_2 _4071_ (.A(_1141_),
    .Y(_1142_));
 sky130_fd_sc_hd__a221o_1 _4072_ (.A1(_0471_),
    .A2(_0834_),
    .B1(_0839_),
    .B2(_1129_),
    .C1(_0814_),
    .X(_1143_));
 sky130_fd_sc_hd__nor2_1 _4073_ (.A(_0471_),
    .B(_0836_),
    .Y(_1144_));
 sky130_fd_sc_hd__a211o_1 _4074_ (.A1(_0471_),
    .A2(_0851_),
    .B1(_1144_),
    .C1(_0834_),
    .X(_1145_));
 sky130_fd_sc_hd__a221o_1 _4075_ (.A1(\z80.tv80s.i_tv80_core.BusA[4] ),
    .A2(_0844_),
    .B1(_1145_),
    .B2(\z80.tv80s.i_tv80_core.BusB[4] ),
    .C1(_1143_),
    .X(_1146_));
 sky130_fd_sc_hd__o22a_1 _4076_ (.A1(_0813_),
    .A2(_1142_),
    .B1(_1146_),
    .B2(_1128_),
    .X(_1147_));
 sky130_fd_sc_hd__mux2_1 _4077_ (.A0(\z80.tv80s.di_reg[4] ),
    .A1(_1147_),
    .S(\z80.tv80s.i_tv80_core.Save_ALU_r ),
    .X(_1148_));
 sky130_fd_sc_hd__and2_1 _4078_ (.A(net728),
    .B(_0811_),
    .X(_1149_));
 sky130_fd_sc_hd__a21oi_4 _4079_ (.A1(_0812_),
    .A2(_1148_),
    .B1(_1149_),
    .Y(_1150_));
 sky130_fd_sc_hd__inv_2 _4080_ (.A(_1150_),
    .Y(_1151_));
 sky130_fd_sc_hd__o21a_1 _4081_ (.A1(net76),
    .A2(_1150_),
    .B1(net85),
    .X(_1152_));
 sky130_fd_sc_hd__o21ai_1 _4082_ (.A1(_0810_),
    .A2(_1124_),
    .B1(_1152_),
    .Y(_1153_));
 sky130_fd_sc_hd__o21a_1 _4083_ (.A1(net245),
    .A2(net85),
    .B1(net86),
    .X(_1154_));
 sky130_fd_sc_hd__mux4_1 _4084_ (.A0(net433),
    .A1(net323),
    .A2(net424),
    .A3(net397),
    .S0(net74),
    .S1(net83),
    .X(_1155_));
 sky130_fd_sc_hd__a22o_2 _4085_ (.A1(_1153_),
    .A2(_1154_),
    .B1(_1155_),
    .B2(net89),
    .X(_1156_));
 sky130_fd_sc_hd__mux2_1 _4086_ (.A0(_1156_),
    .A1(net472),
    .S(_0808_),
    .X(_0044_));
 sky130_fd_sc_hd__and2_1 _4087_ (.A(net643),
    .B(_0811_),
    .X(_1157_));
 sky130_fd_sc_hd__nor2_1 _4088_ (.A(net111),
    .B(\z80.tv80s.i_tv80_core.BusB[5] ),
    .Y(_1158_));
 sky130_fd_sc_hd__and2_1 _4089_ (.A(net111),
    .B(\z80.tv80s.i_tv80_core.BusB[5] ),
    .X(_1159_));
 sky130_fd_sc_hd__o21a_1 _4090_ (.A1(_1158_),
    .A2(_1159_),
    .B1(\z80.tv80s.i_tv80_core.BusA[5] ),
    .X(_1160_));
 sky130_fd_sc_hd__nor3_1 _4091_ (.A(\z80.tv80s.i_tv80_core.BusA[5] ),
    .B(_1158_),
    .C(_1159_),
    .Y(_1161_));
 sky130_fd_sc_hd__nor2_1 _4092_ (.A(_1160_),
    .B(_1161_),
    .Y(_1162_));
 sky130_fd_sc_hd__a21bo_1 _4093_ (.A1(_1135_),
    .A2(_1136_),
    .B1_N(_1133_),
    .X(_1163_));
 sky130_fd_sc_hd__nand2_1 _4094_ (.A(_1162_),
    .B(_1163_),
    .Y(_1164_));
 sky130_fd_sc_hd__or2_1 _4095_ (.A(_1162_),
    .B(_1163_),
    .X(_1165_));
 sky130_fd_sc_hd__or2_1 _4096_ (.A(net143),
    .B(_1160_),
    .X(_1166_));
 sky130_fd_sc_hd__a22o_1 _4097_ (.A1(_0828_),
    .A2(_1162_),
    .B1(_1166_),
    .B2(_0815_),
    .X(_1167_));
 sky130_fd_sc_hd__a31o_1 _4098_ (.A1(_0827_),
    .A2(_1164_),
    .A3(_1165_),
    .B1(_1167_),
    .X(_1168_));
 sky130_fd_sc_hd__o41a_2 _4099_ (.A1(_2864_),
    .A2(\z80.tv80s.i_tv80_core.BusA[5] ),
    .A3(\z80.tv80s.i_tv80_core.BusB[5] ),
    .A4(_0827_),
    .B1(_1168_),
    .X(_1169_));
 sky130_fd_sc_hd__and2_1 _4100_ (.A(\z80.tv80s.i_tv80_core.BusA[4] ),
    .B(_1006_),
    .X(_1170_));
 sky130_fd_sc_hd__nor2_1 _4101_ (.A(\z80.tv80s.i_tv80_core.BusA[5] ),
    .B(_1170_),
    .Y(_1171_));
 sky130_fd_sc_hd__o31a_1 _4102_ (.A1(\z80.tv80s.i_tv80_core.BusA[5] ),
    .A2(\z80.tv80s.i_tv80_core.BusA[6] ),
    .A3(_1170_),
    .B1(net162),
    .X(_1172_));
 sky130_fd_sc_hd__nor2_1 _4103_ (.A(\z80.tv80s.i_tv80_core.F[0] ),
    .B(_1172_),
    .Y(_1173_));
 sky130_fd_sc_hd__or2_4 _4104_ (.A(\z80.tv80s.i_tv80_core.F[0] ),
    .B(_1172_),
    .X(_1174_));
 sky130_fd_sc_hd__and3_1 _4105_ (.A(\z80.tv80s.i_tv80_core.BusA[4] ),
    .B(\z80.tv80s.i_tv80_core.BusA[5] ),
    .C(_1006_),
    .X(_1175_));
 sky130_fd_sc_hd__or2_1 _4106_ (.A(_1171_),
    .B(_1175_),
    .X(_1176_));
 sky130_fd_sc_hd__or3_1 _4107_ (.A(\z80.tv80s.i_tv80_core.BusA[4] ),
    .B(_1008_),
    .C(_1084_),
    .X(_1177_));
 sky130_fd_sc_hd__or2_1 _4108_ (.A(\z80.tv80s.i_tv80_core.BusA[5] ),
    .B(_1177_),
    .X(_1178_));
 sky130_fd_sc_hd__xor2_1 _4109_ (.A(\z80.tv80s.i_tv80_core.BusA[5] ),
    .B(_1177_),
    .X(_1179_));
 sky130_fd_sc_hd__mux2_1 _4110_ (.A0(_1176_),
    .A1(_1179_),
    .S(\z80.tv80s.i_tv80_core.F[1] ),
    .X(_1180_));
 sky130_fd_sc_hd__xnor2_2 _4111_ (.A(_1174_),
    .B(_1180_),
    .Y(_1181_));
 sky130_fd_sc_hd__inv_2 _4112_ (.A(_1181_),
    .Y(_1182_));
 sky130_fd_sc_hd__a22o_1 _4113_ (.A1(\z80.tv80s.i_tv80_core.BusA[5] ),
    .A2(_0844_),
    .B1(_0848_),
    .B2(_1181_),
    .X(_1183_));
 sky130_fd_sc_hd__mux2_1 _4114_ (.A0(\z80.tv80s.i_tv80_core.BusA[4] ),
    .A1(\z80.tv80s.i_tv80_core.BusA[6] ),
    .S(net154),
    .X(_1184_));
 sky130_fd_sc_hd__and2_1 _4115_ (.A(_0839_),
    .B(_1184_),
    .X(_1185_));
 sky130_fd_sc_hd__nor2_1 _4116_ (.A(_0470_),
    .B(_0836_),
    .Y(_1186_));
 sky130_fd_sc_hd__a211o_1 _4117_ (.A1(_0470_),
    .A2(_0851_),
    .B1(_1186_),
    .C1(_0834_),
    .X(_1187_));
 sky130_fd_sc_hd__a221o_1 _4118_ (.A1(_0470_),
    .A2(_0834_),
    .B1(_1187_),
    .B2(\z80.tv80s.i_tv80_core.BusB[5] ),
    .C1(_1185_),
    .X(_1188_));
 sky130_fd_sc_hd__a211o_1 _4119_ (.A1(_0814_),
    .A2(_1169_),
    .B1(_1183_),
    .C1(_1188_),
    .X(_1189_));
 sky130_fd_sc_hd__mux2_1 _4120_ (.A0(\z80.tv80s.di_reg[5] ),
    .A1(_1189_),
    .S(\z80.tv80s.i_tv80_core.Save_ALU_r ),
    .X(_1190_));
 sky130_fd_sc_hd__a21oi_4 _4121_ (.A1(_0812_),
    .A2(_1190_),
    .B1(_1157_),
    .Y(_1191_));
 sky130_fd_sc_hd__inv_2 _4122_ (.A(_1191_),
    .Y(_1192_));
 sky130_fd_sc_hd__o21ai_1 _4123_ (.A1(net76),
    .A2(_1191_),
    .B1(net85),
    .Y(_1193_));
 sky130_fd_sc_hd__a22o_1 _4124_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][5] ),
    .A2(_0868_),
    .B1(_0870_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][5] ),
    .X(_1194_));
 sky130_fd_sc_hd__a221o_1 _4125_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][5] ),
    .A2(_0874_),
    .B1(_0876_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][5] ),
    .C1(_1194_),
    .X(_1195_));
 sky130_fd_sc_hd__a22o_1 _4126_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][5] ),
    .A2(_0879_),
    .B1(_0882_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][5] ),
    .X(_1196_));
 sky130_fd_sc_hd__a221o_1 _4127_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][5] ),
    .A2(_0806_),
    .B1(_0885_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][5] ),
    .C1(_1196_),
    .X(_1197_));
 sky130_fd_sc_hd__or2_2 _4128_ (.A(_1195_),
    .B(_1197_),
    .X(_1198_));
 sky130_fd_sc_hd__nand2_1 _4129_ (.A(net80),
    .B(_1198_),
    .Y(_1199_));
 sky130_fd_sc_hd__inv_2 _4130_ (.A(_1199_),
    .Y(_1200_));
 sky130_fd_sc_hd__nor2_1 _4131_ (.A(net80),
    .B(_1198_),
    .Y(_1201_));
 sky130_fd_sc_hd__nor2_1 _4132_ (.A(_1200_),
    .B(_1201_),
    .Y(_1202_));
 sky130_fd_sc_hd__a22oi_2 _4133_ (.A1(net80),
    .A2(_1122_),
    .B1(_1123_),
    .B2(_1117_),
    .Y(_1203_));
 sky130_fd_sc_hd__xnor2_1 _4134_ (.A(_1202_),
    .B(_1203_),
    .Y(_1204_));
 sky130_fd_sc_hd__a21o_1 _4135_ (.A1(net76),
    .A2(_1204_),
    .B1(_1193_),
    .X(_1205_));
 sky130_fd_sc_hd__o21a_1 _4136_ (.A1(net241),
    .A2(net85),
    .B1(net86),
    .X(_1206_));
 sky130_fd_sc_hd__mux4_1 _4137_ (.A0(net410),
    .A1(net401),
    .A2(net428),
    .A3(net325),
    .S0(net74),
    .S1(net82),
    .X(_1207_));
 sky130_fd_sc_hd__a22o_2 _4138_ (.A1(_1205_),
    .A2(_1206_),
    .B1(_1207_),
    .B2(net89),
    .X(_1208_));
 sky130_fd_sc_hd__mux2_1 _4139_ (.A0(_1208_),
    .A1(net443),
    .S(_0808_),
    .X(_0045_));
 sky130_fd_sc_hd__a22o_1 _4140_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][6] ),
    .A2(_0868_),
    .B1(_0870_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][6] ),
    .X(_1209_));
 sky130_fd_sc_hd__a221o_1 _4141_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][6] ),
    .A2(_0874_),
    .B1(_0876_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][6] ),
    .C1(_1209_),
    .X(_1210_));
 sky130_fd_sc_hd__a22o_1 _4142_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][6] ),
    .A2(_0879_),
    .B1(_0882_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][6] ),
    .X(_1211_));
 sky130_fd_sc_hd__a221o_1 _4143_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][6] ),
    .A2(_0806_),
    .B1(_0885_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][6] ),
    .C1(_1211_),
    .X(_1212_));
 sky130_fd_sc_hd__or2_2 _4144_ (.A(_1210_),
    .B(_1212_),
    .X(_1213_));
 sky130_fd_sc_hd__and2_1 _4145_ (.A(net80),
    .B(_1213_),
    .X(_1214_));
 sky130_fd_sc_hd__nor2_1 _4146_ (.A(net80),
    .B(_1213_),
    .Y(_1215_));
 sky130_fd_sc_hd__nor2_1 _4147_ (.A(_1214_),
    .B(_1215_),
    .Y(_1216_));
 sky130_fd_sc_hd__o21ai_1 _4148_ (.A1(_1201_),
    .A2(_1203_),
    .B1(_1199_),
    .Y(_1217_));
 sky130_fd_sc_hd__xor2_1 _4149_ (.A(_1216_),
    .B(_1217_),
    .X(_1218_));
 sky130_fd_sc_hd__xor2_1 _4150_ (.A(net143),
    .B(\z80.tv80s.i_tv80_core.BusB[6] ),
    .X(_1219_));
 sky130_fd_sc_hd__and2_1 _4151_ (.A(\z80.tv80s.i_tv80_core.BusA[6] ),
    .B(_1219_),
    .X(_1220_));
 sky130_fd_sc_hd__nor2_1 _4152_ (.A(\z80.tv80s.i_tv80_core.BusA[6] ),
    .B(_1219_),
    .Y(_1221_));
 sky130_fd_sc_hd__nor2_1 _4153_ (.A(_1220_),
    .B(_1221_),
    .Y(_1222_));
 sky130_fd_sc_hd__a21o_1 _4154_ (.A1(_1162_),
    .A2(_1163_),
    .B1(_1160_),
    .X(_1223_));
 sky130_fd_sc_hd__xnor2_1 _4155_ (.A(_1222_),
    .B(_1223_),
    .Y(_1224_));
 sky130_fd_sc_hd__nor2_1 _4156_ (.A(_0826_),
    .B(_1224_),
    .Y(_1225_));
 sky130_fd_sc_hd__or2_1 _4157_ (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[1] ),
    .B(_1220_),
    .X(_1226_));
 sky130_fd_sc_hd__a221o_1 _4158_ (.A1(_0828_),
    .A2(_1222_),
    .B1(_1226_),
    .B2(_0815_),
    .C1(_1225_),
    .X(_1227_));
 sky130_fd_sc_hd__o41a_2 _4159_ (.A1(net111),
    .A2(\z80.tv80s.i_tv80_core.BusA[6] ),
    .A3(\z80.tv80s.i_tv80_core.BusB[6] ),
    .A4(_0827_),
    .B1(_1227_),
    .X(_1228_));
 sky130_fd_sc_hd__xnor2_1 _4160_ (.A(\z80.tv80s.i_tv80_core.BusA[6] ),
    .B(_1175_),
    .Y(_1229_));
 sky130_fd_sc_hd__a21o_1 _4161_ (.A1(_1174_),
    .A2(_1176_),
    .B1(_1229_),
    .X(_1230_));
 sky130_fd_sc_hd__nand2_1 _4162_ (.A(_1176_),
    .B(_1229_),
    .Y(_1231_));
 sky130_fd_sc_hd__o21ai_1 _4163_ (.A1(_1173_),
    .A2(_1231_),
    .B1(_1230_),
    .Y(_1232_));
 sky130_fd_sc_hd__xor2_1 _4164_ (.A(\z80.tv80s.i_tv80_core.BusA[6] ),
    .B(_1178_),
    .X(_1233_));
 sky130_fd_sc_hd__nor2_1 _4165_ (.A(_1173_),
    .B(_1179_),
    .Y(_1234_));
 sky130_fd_sc_hd__xnor2_1 _4166_ (.A(_1233_),
    .B(_1234_),
    .Y(_1235_));
 sky130_fd_sc_hd__mux2_2 _4167_ (.A0(_1232_),
    .A1(_1235_),
    .S(\z80.tv80s.i_tv80_core.F[1] ),
    .X(_1236_));
 sky130_fd_sc_hd__nor2_1 _4168_ (.A(_0405_),
    .B(_0836_),
    .Y(_1237_));
 sky130_fd_sc_hd__mux2_1 _4169_ (.A0(\z80.tv80s.i_tv80_core.BusA[5] ),
    .A1(net162),
    .S(net154),
    .X(_1238_));
 sky130_fd_sc_hd__a221o_1 _4170_ (.A1(\z80.tv80s.i_tv80_core.BusA[6] ),
    .A2(_0844_),
    .B1(_1238_),
    .B2(_0839_),
    .C1(_0814_),
    .X(_1239_));
 sky130_fd_sc_hd__a211o_1 _4171_ (.A1(_0405_),
    .A2(_0851_),
    .B1(_1237_),
    .C1(_0834_),
    .X(_1240_));
 sky130_fd_sc_hd__a22o_1 _4172_ (.A1(_0405_),
    .A2(_0834_),
    .B1(_1240_),
    .B2(\z80.tv80s.i_tv80_core.BusB[6] ),
    .X(_1241_));
 sky130_fd_sc_hd__a211o_1 _4173_ (.A1(_0848_),
    .A2(_1236_),
    .B1(_1239_),
    .C1(_1241_),
    .X(_1242_));
 sky130_fd_sc_hd__o211a_1 _4174_ (.A1(_0813_),
    .A2(_1228_),
    .B1(_1242_),
    .C1(\z80.tv80s.i_tv80_core.Save_ALU_r ),
    .X(_1243_));
 sky130_fd_sc_hd__a21oi_1 _4175_ (.A1(_2861_),
    .A2(\z80.tv80s.di_reg[6] ),
    .B1(_1243_),
    .Y(_1244_));
 sky130_fd_sc_hd__mux2_4 _4176_ (.A0(_2869_),
    .A1(_1244_),
    .S(_0812_),
    .X(_1245_));
 sky130_fd_sc_hd__inv_2 _4177_ (.A(_1245_),
    .Y(_1246_));
 sky130_fd_sc_hd__nor2_1 _4178_ (.A(net76),
    .B(_1245_),
    .Y(_1247_));
 sky130_fd_sc_hd__a211o_1 _4179_ (.A1(net76),
    .A2(_1218_),
    .B1(_1247_),
    .C1(_0774_),
    .X(_1248_));
 sky130_fd_sc_hd__o21a_1 _4180_ (.A1(net227),
    .A2(net85),
    .B1(net86),
    .X(_1249_));
 sky130_fd_sc_hd__mux4_2 _4181_ (.A0(net358),
    .A1(net334),
    .A2(net348),
    .A3(net336),
    .S0(net74),
    .S1(net82),
    .X(_1250_));
 sky130_fd_sc_hd__a22o_2 _4182_ (.A1(_1248_),
    .A2(_1249_),
    .B1(_1250_),
    .B2(net89),
    .X(_1251_));
 sky130_fd_sc_hd__mux2_1 _4183_ (.A0(_1251_),
    .A1(net437),
    .S(_0808_),
    .X(_0046_));
 sky130_fd_sc_hd__a21o_1 _4184_ (.A1(_1216_),
    .A2(_1217_),
    .B1(_1214_),
    .X(_1252_));
 sky130_fd_sc_hd__a22o_1 _4185_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][7] ),
    .A2(_0874_),
    .B1(_0876_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][7] ),
    .X(_1253_));
 sky130_fd_sc_hd__a221o_1 _4186_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][7] ),
    .A2(_0868_),
    .B1(_0870_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][7] ),
    .C1(_1253_),
    .X(_1254_));
 sky130_fd_sc_hd__a22o_1 _4187_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][7] ),
    .A2(_0879_),
    .B1(_0882_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][7] ),
    .X(_1255_));
 sky130_fd_sc_hd__a221o_1 _4188_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][7] ),
    .A2(_0806_),
    .B1(_0885_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][7] ),
    .C1(_1255_),
    .X(_1256_));
 sky130_fd_sc_hd__or2_1 _4189_ (.A(_1254_),
    .B(_1256_),
    .X(_1257_));
 sky130_fd_sc_hd__xnor2_1 _4190_ (.A(net80),
    .B(_1257_),
    .Y(_1258_));
 sky130_fd_sc_hd__xnor2_1 _4191_ (.A(_1252_),
    .B(_1258_),
    .Y(_1259_));
 sky130_fd_sc_hd__a21o_1 _4192_ (.A1(_1222_),
    .A2(_1223_),
    .B1(_1220_),
    .X(_1260_));
 sky130_fd_sc_hd__xor2_1 _4193_ (.A(net162),
    .B(_1260_),
    .X(_1261_));
 sky130_fd_sc_hd__xor2_1 _4194_ (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[1] ),
    .B(\z80.tv80s.i_tv80_core.BusB[7] ),
    .X(_1262_));
 sky130_fd_sc_hd__or2_1 _4195_ (.A(_1261_),
    .B(_1262_),
    .X(_1263_));
 sky130_fd_sc_hd__nand2_1 _4196_ (.A(_1261_),
    .B(_1262_),
    .Y(_1264_));
 sky130_fd_sc_hd__or2_1 _4197_ (.A(net162),
    .B(\z80.tv80s.i_tv80_core.BusB[7] ),
    .X(_1265_));
 sky130_fd_sc_hd__nand2_1 _4198_ (.A(net162),
    .B(\z80.tv80s.i_tv80_core.BusB[7] ),
    .Y(_1266_));
 sky130_fd_sc_hd__nand2_1 _4199_ (.A(_2864_),
    .B(_1266_),
    .Y(_1267_));
 sky130_fd_sc_hd__a32o_1 _4200_ (.A1(_0828_),
    .A2(_1265_),
    .A3(_1266_),
    .B1(_1267_),
    .B2(_0815_),
    .X(_1268_));
 sky130_fd_sc_hd__a31o_1 _4201_ (.A1(_0827_),
    .A2(_1263_),
    .A3(_1264_),
    .B1(_1268_),
    .X(_1269_));
 sky130_fd_sc_hd__o41a_2 _4202_ (.A1(net111),
    .A2(net162),
    .A3(\z80.tv80s.i_tv80_core.BusB[7] ),
    .A4(_0827_),
    .B1(_1269_),
    .X(_1270_));
 sky130_fd_sc_hd__nand2_1 _4203_ (.A(_1174_),
    .B(_1231_),
    .Y(_1271_));
 sky130_fd_sc_hd__xor2_1 _4204_ (.A(net162),
    .B(\z80.tv80s.i_tv80_core.BusA[6] ),
    .X(_1272_));
 sky130_fd_sc_hd__mux2_1 _4205_ (.A0(net162),
    .A1(_1272_),
    .S(_1175_),
    .X(_1273_));
 sky130_fd_sc_hd__xnor2_1 _4206_ (.A(_1271_),
    .B(_1273_),
    .Y(_1274_));
 sky130_fd_sc_hd__or3_1 _4207_ (.A(net162),
    .B(\z80.tv80s.i_tv80_core.BusA[6] ),
    .C(_1178_),
    .X(_1275_));
 sky130_fd_sc_hd__o21ai_1 _4208_ (.A1(\z80.tv80s.i_tv80_core.BusA[6] ),
    .A2(_1178_),
    .B1(\z80.tv80s.i_tv80_core.BusA[7] ),
    .Y(_1276_));
 sky130_fd_sc_hd__nand2_1 _4209_ (.A(_1275_),
    .B(_1276_),
    .Y(_1277_));
 sky130_fd_sc_hd__nor2_1 _4210_ (.A(_1179_),
    .B(_1233_),
    .Y(_1278_));
 sky130_fd_sc_hd__nor2_1 _4211_ (.A(_1277_),
    .B(_1278_),
    .Y(_1279_));
 sky130_fd_sc_hd__or2_1 _4212_ (.A(_1173_),
    .B(_1278_),
    .X(_1280_));
 sky130_fd_sc_hd__a22o_1 _4213_ (.A1(_1174_),
    .A2(_1279_),
    .B1(_1280_),
    .B2(_1277_),
    .X(_1281_));
 sky130_fd_sc_hd__mux2_1 _4214_ (.A0(_1274_),
    .A1(_1281_),
    .S(\z80.tv80s.i_tv80_core.F[1] ),
    .X(_1282_));
 sky130_fd_sc_hd__a22oi_1 _4215_ (.A1(\z80.tv80s.i_tv80_core.BusA[7] ),
    .A2(_0844_),
    .B1(_0848_),
    .B2(_1282_),
    .Y(_1283_));
 sky130_fd_sc_hd__inv_2 _4216_ (.A(_1283_),
    .Y(_1284_));
 sky130_fd_sc_hd__and2_1 _4217_ (.A(net153),
    .B(\z80.tv80s.i_tv80_core.BusA[0] ),
    .X(_1285_));
 sky130_fd_sc_hd__a22o_1 _4218_ (.A1(net120),
    .A2(\z80.tv80s.i_tv80_core.BusA[6] ),
    .B1(_2898_),
    .B2(_1285_),
    .X(_1286_));
 sky130_fd_sc_hd__a221o_2 _4219_ (.A1(\z80.tv80s.i_tv80_core.F[0] ),
    .A2(_0468_),
    .B1(_0470_),
    .B2(net162),
    .C1(_1286_),
    .X(_1287_));
 sky130_fd_sc_hd__or2_1 _4220_ (.A(\z80.tv80s.i_tv80_core.BusB[7] ),
    .B(_0474_),
    .X(_1288_));
 sky130_fd_sc_hd__o211a_1 _4221_ (.A1(_2863_),
    .A2(_0475_),
    .B1(_0832_),
    .C1(_1288_),
    .X(_1289_));
 sky130_fd_sc_hd__and2_1 _4222_ (.A(\z80.tv80s.i_tv80_core.BusB[7] ),
    .B(_0474_),
    .X(_1290_));
 sky130_fd_sc_hd__and2_1 _4223_ (.A(_0851_),
    .B(_1290_),
    .X(_1291_));
 sky130_fd_sc_hd__a211o_1 _4224_ (.A1(_0839_),
    .A2(_1287_),
    .B1(_1289_),
    .C1(_1291_),
    .X(_1292_));
 sky130_fd_sc_hd__a211o_1 _4225_ (.A1(_0814_),
    .A2(_1270_),
    .B1(_1284_),
    .C1(_1292_),
    .X(_1293_));
 sky130_fd_sc_hd__mux2_1 _4226_ (.A0(\z80.tv80s.di_reg[7] ),
    .A1(_1293_),
    .S(net877),
    .X(_1294_));
 sky130_fd_sc_hd__mux2_4 _4227_ (.A0(net639),
    .A1(_1294_),
    .S(_0812_),
    .X(_1295_));
 sky130_fd_sc_hd__a21o_1 _4228_ (.A1(_0810_),
    .A2(_1295_),
    .B1(_0774_),
    .X(_1296_));
 sky130_fd_sc_hd__a21o_1 _4229_ (.A1(net76),
    .A2(_1259_),
    .B1(_1296_),
    .X(_1297_));
 sky130_fd_sc_hd__o21a_1 _4230_ (.A1(net231),
    .A2(net85),
    .B1(net86),
    .X(_1298_));
 sky130_fd_sc_hd__and2_4 _4231_ (.A(\z80.tv80s.i_tv80_core.RegAddrB_r[1] ),
    .B(net86),
    .X(_1299_));
 sky130_fd_sc_hd__nand2_4 _4232_ (.A(\z80.tv80s.i_tv80_core.RegAddrB_r[1] ),
    .B(net86),
    .Y(_1300_));
 sky130_fd_sc_hd__or3_1 _4233_ (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][7] ),
    .B(net142),
    .C(net89),
    .X(_1301_));
 sky130_fd_sc_hd__o211a_1 _4234_ (.A1(net341),
    .A2(net82),
    .B1(net74),
    .C1(_1301_),
    .X(_1302_));
 sky130_fd_sc_hd__mux2_1 _4235_ (.A0(net387),
    .A1(net373),
    .S(net83),
    .X(_1303_));
 sky130_fd_sc_hd__o221a_1 _4236_ (.A1(net403),
    .A2(net142),
    .B1(net83),
    .B2(net365),
    .C1(net75),
    .X(_1304_));
 sky130_fd_sc_hd__o221a_1 _4237_ (.A1(net462),
    .A2(net142),
    .B1(net83),
    .B2(net454),
    .C1(net73),
    .X(_1305_));
 sky130_fd_sc_hd__a211o_1 _4238_ (.A1(net73),
    .A2(_1303_),
    .B1(_1302_),
    .C1(_1299_),
    .X(_1306_));
 sky130_fd_sc_hd__o31a_1 _4239_ (.A1(_1300_),
    .A2(_1304_),
    .A3(_1305_),
    .B1(_1306_),
    .X(_1307_));
 sky130_fd_sc_hd__a22o_2 _4240_ (.A1(_1297_),
    .A2(_1298_),
    .B1(_1307_),
    .B2(net89),
    .X(_1308_));
 sky130_fd_sc_hd__mux2_1 _4241_ (.A0(_1308_),
    .A1(net454),
    .S(_0808_),
    .X(_0047_));
 sky130_fd_sc_hd__nand2_1 _4242_ (.A(net132),
    .B(_0406_),
    .Y(_1309_));
 sky130_fd_sc_hd__a31o_1 _4243_ (.A1(net109),
    .A2(_0407_),
    .A3(_1309_),
    .B1(net118),
    .X(_1310_));
 sky130_fd_sc_hd__inv_2 _4244_ (.A(_1310_),
    .Y(_1311_));
 sky130_fd_sc_hd__o21a_1 _4245_ (.A1(net97),
    .A2(_0461_),
    .B1(_2971_),
    .X(_1312_));
 sky130_fd_sc_hd__nor2_1 _4246_ (.A(_2930_),
    .B(_0477_),
    .Y(_1313_));
 sky130_fd_sc_hd__or2_1 _4247_ (.A(_2933_),
    .B(_1313_),
    .X(_1314_));
 sky130_fd_sc_hd__and3_1 _4248_ (.A(\z80.tv80s.i_tv80_core.i_mcode.MCycle[1] ),
    .B(_2896_),
    .C(_2982_),
    .X(_1315_));
 sky130_fd_sc_hd__or2_1 _4249_ (.A(_1314_),
    .B(_1315_),
    .X(_1316_));
 sky130_fd_sc_hd__or2_1 _4250_ (.A(_1312_),
    .B(_1316_),
    .X(_1317_));
 sky130_fd_sc_hd__nor2_1 _4251_ (.A(_0406_),
    .B(_0461_),
    .Y(_1318_));
 sky130_fd_sc_hd__or3b_1 _4252_ (.A(_2912_),
    .B(_2947_),
    .C_N(_0705_),
    .X(_1319_));
 sky130_fd_sc_hd__nor2_1 _4253_ (.A(_0434_),
    .B(_1318_),
    .Y(_1320_));
 sky130_fd_sc_hd__o32a_1 _4254_ (.A1(net137),
    .A2(_0397_),
    .A3(_0427_),
    .B1(_0430_),
    .B2(_1309_),
    .X(_1321_));
 sky130_fd_sc_hd__inv_2 _4255_ (.A(_1321_),
    .Y(_1322_));
 sky130_fd_sc_hd__o31a_1 _4256_ (.A1(net109),
    .A2(_1320_),
    .A3(_1322_),
    .B1(net148),
    .X(_1323_));
 sky130_fd_sc_hd__a311o_1 _4257_ (.A1(_2965_),
    .A2(_3001_),
    .A3(_0398_),
    .B1(_1317_),
    .C1(_1323_),
    .X(_1324_));
 sky130_fd_sc_hd__a221o_1 _4258_ (.A1(net159),
    .A2(net163),
    .B1(_1311_),
    .B2(_1324_),
    .C1(net106),
    .X(_1325_));
 sky130_fd_sc_hd__and3b_1 _4259_ (.A_N(_2907_),
    .B(net109),
    .C(_2849_),
    .X(_1326_));
 sky130_fd_sc_hd__or3_1 _4260_ (.A(net135),
    .B(_2907_),
    .C(net108),
    .X(_1327_));
 sky130_fd_sc_hd__nor2_1 _4261_ (.A(_1309_),
    .B(_1327_),
    .Y(_1328_));
 sky130_fd_sc_hd__nand2b_1 _4262_ (.A_N(_2999_),
    .B(_0760_),
    .Y(_1329_));
 sky130_fd_sc_hd__or2_1 _4263_ (.A(_0388_),
    .B(_0558_),
    .X(_1330_));
 sky130_fd_sc_hd__and3_2 _4264_ (.A(net152),
    .B(_0390_),
    .C(_0659_),
    .X(_1331_));
 sky130_fd_sc_hd__a221o_1 _4265_ (.A1(net147),
    .A2(_1328_),
    .B1(_1331_),
    .B2(_3001_),
    .C1(_1330_),
    .X(_1332_));
 sky130_fd_sc_hd__o21ai_4 _4266_ (.A1(_1329_),
    .A2(_1332_),
    .B1(_1325_),
    .Y(_1333_));
 sky130_fd_sc_hd__nor2_1 _4267_ (.A(net137),
    .B(_0427_),
    .Y(_1334_));
 sky130_fd_sc_hd__nor2_1 _4268_ (.A(net149),
    .B(_2848_),
    .Y(_1335_));
 sky130_fd_sc_hd__o21a_1 _4269_ (.A1(_0512_),
    .A2(_1335_),
    .B1(_1334_),
    .X(_1336_));
 sky130_fd_sc_hd__o21a_1 _4270_ (.A1(_1320_),
    .A2(_1336_),
    .B1(net146),
    .X(_1337_));
 sky130_fd_sc_hd__o21a_1 _4271_ (.A1(net131),
    .A2(_0553_),
    .B1(_0488_),
    .X(_1338_));
 sky130_fd_sc_hd__a31o_1 _4272_ (.A1(net152),
    .A2(_2962_),
    .A3(_0659_),
    .B1(_1338_),
    .X(_1339_));
 sky130_fd_sc_hd__and2_1 _4273_ (.A(net145),
    .B(_3029_),
    .X(_1340_));
 sky130_fd_sc_hd__a311o_1 _4274_ (.A1(net132),
    .A2(_0429_),
    .A3(_1340_),
    .B1(_0684_),
    .C1(net109),
    .X(_1341_));
 sky130_fd_sc_hd__a311o_1 _4275_ (.A1(_2934_),
    .A2(_2965_),
    .A3(_0398_),
    .B1(_1317_),
    .C1(_1341_),
    .X(_1342_));
 sky130_fd_sc_hd__or2_1 _4276_ (.A(net132),
    .B(net97),
    .X(_1343_));
 sky130_fd_sc_hd__a21o_1 _4277_ (.A1(_1340_),
    .A2(_1343_),
    .B1(net108),
    .X(_1344_));
 sky130_fd_sc_hd__o311a_1 _4278_ (.A1(_1337_),
    .A2(_1339_),
    .A3(_1342_),
    .B1(_1344_),
    .C1(net166),
    .X(_1345_));
 sky130_fd_sc_hd__a211o_1 _4279_ (.A1(net157),
    .A2(net163),
    .B1(net106),
    .C1(_1345_),
    .X(_1346_));
 sky130_fd_sc_hd__a32o_1 _4280_ (.A1(net132),
    .A2(_1326_),
    .A3(_1340_),
    .B1(_1331_),
    .B2(_2934_),
    .X(_1347_));
 sky130_fd_sc_hd__or4b_2 _4281_ (.A(_0678_),
    .B(_1330_),
    .C(_1347_),
    .D_N(_0760_),
    .X(_1348_));
 sky130_fd_sc_hd__nand2_4 _4282_ (.A(_1346_),
    .B(_1348_),
    .Y(_1349_));
 sky130_fd_sc_hd__inv_2 _4283_ (.A(_1349_),
    .Y(_1350_));
 sky130_fd_sc_hd__or3_1 _4284_ (.A(\z80.tv80s.i_tv80_core.XY_Ind ),
    .B(_0500_),
    .C(_1349_),
    .X(_1351_));
 sky130_fd_sc_hd__nand2b_1 _4285_ (.A_N(_1351_),
    .B(_1333_),
    .Y(_1352_));
 sky130_fd_sc_hd__mux2_1 _4286_ (.A0(\z80.tv80s.i_tv80_core.XY_State[1] ),
    .A1(\z80.tv80s.i_tv80_core.Alternate ),
    .S(_1352_),
    .X(_1353_));
 sky130_fd_sc_hd__mux2_1 _4287_ (.A0(net225),
    .A1(_1353_),
    .S(net113),
    .X(_0048_));
 sky130_fd_sc_hd__and2_1 _4288_ (.A(_2998_),
    .B(net107),
    .X(_1354_));
 sky130_fd_sc_hd__and3_4 _4289_ (.A(net154),
    .B(_2998_),
    .C(net107),
    .X(_1355_));
 sky130_fd_sc_hd__and3_2 _4290_ (.A(_2846_),
    .B(net122),
    .C(_1355_),
    .X(_1356_));
 sky130_fd_sc_hd__or3b_4 _4291_ (.A(net147),
    .B(_2854_),
    .C_N(_1355_),
    .X(_1357_));
 sky130_fd_sc_hd__and3_1 _4292_ (.A(net137),
    .B(net558),
    .C(_0603_),
    .X(_1358_));
 sky130_fd_sc_hd__o21ai_1 _4293_ (.A1(net558),
    .A2(_0607_),
    .B1(_1357_),
    .Y(_1359_));
 sky130_fd_sc_hd__a2bb2o_1 _4294_ (.A1_N(_1358_),
    .A2_N(_1359_),
    .B1(\z80.tv80s.i_tv80_core.ACC[0] ),
    .B2(_1356_),
    .X(_1360_));
 sky130_fd_sc_hd__mux2_1 _4295_ (.A0(net558),
    .A1(_1360_),
    .S(net115),
    .X(_0049_));
 sky130_fd_sc_hd__or2_1 _4296_ (.A(net615),
    .B(_1358_),
    .X(_1361_));
 sky130_fd_sc_hd__a21oi_1 _4297_ (.A1(net615),
    .A2(_1358_),
    .B1(_1356_),
    .Y(_1362_));
 sky130_fd_sc_hd__a22o_1 _4298_ (.A1(\z80.tv80s.i_tv80_core.ACC[1] ),
    .A2(_1356_),
    .B1(_1361_),
    .B2(_1362_),
    .X(_1363_));
 sky130_fd_sc_hd__mux2_1 _4299_ (.A0(net615),
    .A1(_1363_),
    .S(net115),
    .X(_0050_));
 sky130_fd_sc_hd__nor2_1 _4300_ (.A(net128),
    .B(_1362_),
    .Y(_1364_));
 sky130_fd_sc_hd__mux2_1 _4301_ (.A0(\z80.tv80s.i_tv80_core.ACC[2] ),
    .A1(_2877_),
    .S(_1357_),
    .X(_1365_));
 sky130_fd_sc_hd__mux2_1 _4302_ (.A0(net544),
    .A1(_1365_),
    .S(_1364_),
    .X(_0051_));
 sky130_fd_sc_hd__and3_1 _4303_ (.A(net558),
    .B(\z80.tv80s.i_tv80_core.R[1] ),
    .C(net544),
    .X(_1366_));
 sky130_fd_sc_hd__a31o_1 _4304_ (.A1(net137),
    .A2(_0603_),
    .A3(_1366_),
    .B1(net527),
    .X(_1367_));
 sky130_fd_sc_hd__nand4_1 _4305_ (.A(net527),
    .B(net102),
    .C(_0603_),
    .D(_1366_),
    .Y(_1368_));
 sky130_fd_sc_hd__a21o_1 _4306_ (.A1(_1357_),
    .A2(_1368_),
    .B1(net128),
    .X(_1369_));
 sky130_fd_sc_hd__a22o_1 _4307_ (.A1(\z80.tv80s.i_tv80_core.ACC[3] ),
    .A2(_1356_),
    .B1(_1367_),
    .B2(_1369_),
    .X(_1370_));
 sky130_fd_sc_hd__o21a_1 _4308_ (.A1(net117),
    .A2(net527),
    .B1(_1370_),
    .X(_0052_));
 sky130_fd_sc_hd__nor2_1 _4309_ (.A(net613),
    .B(_1368_),
    .Y(_1371_));
 sky130_fd_sc_hd__mux2_1 _4310_ (.A0(\z80.tv80s.i_tv80_core.ACC[4] ),
    .A1(_1371_),
    .S(_1357_),
    .X(_1372_));
 sky130_fd_sc_hd__a22o_1 _4311_ (.A1(net613),
    .A2(_1369_),
    .B1(_1372_),
    .B2(net117),
    .X(_0053_));
 sky130_fd_sc_hd__and4_1 _4312_ (.A(net527),
    .B(net613),
    .C(_0603_),
    .D(_1366_),
    .X(_1373_));
 sky130_fd_sc_hd__and3_1 _4313_ (.A(net137),
    .B(net564),
    .C(_1373_),
    .X(_1374_));
 sky130_fd_sc_hd__a21oi_1 _4314_ (.A1(net137),
    .A2(_1373_),
    .B1(net564),
    .Y(_1375_));
 sky130_fd_sc_hd__or3_1 _4315_ (.A(_1356_),
    .B(_1374_),
    .C(_1375_),
    .X(_1376_));
 sky130_fd_sc_hd__o21ai_1 _4316_ (.A1(_2879_),
    .A2(_1357_),
    .B1(_1376_),
    .Y(_1377_));
 sky130_fd_sc_hd__mux2_1 _4317_ (.A0(net564),
    .A1(_1377_),
    .S(net115),
    .X(_0054_));
 sky130_fd_sc_hd__a31o_1 _4318_ (.A1(net137),
    .A2(net564),
    .A3(_1373_),
    .B1(net684),
    .X(_1378_));
 sky130_fd_sc_hd__and4_1 _4319_ (.A(net115),
    .B(net564),
    .C(net102),
    .D(_1373_),
    .X(_1379_));
 sky130_fd_sc_hd__nand2_1 _4320_ (.A(net684),
    .B(_1379_),
    .Y(_1380_));
 sky130_fd_sc_hd__a21o_1 _4321_ (.A1(_1378_),
    .A2(_1380_),
    .B1(_1356_),
    .X(_1381_));
 sky130_fd_sc_hd__nand2_1 _4322_ (.A(net117),
    .B(_1356_),
    .Y(_1382_));
 sky130_fd_sc_hd__o221a_1 _4323_ (.A1(net117),
    .A2(net684),
    .B1(_1382_),
    .B2(\z80.tv80s.i_tv80_core.ACC[6] ),
    .C1(_1381_),
    .X(_0055_));
 sky130_fd_sc_hd__or2_1 _4324_ (.A(net651),
    .B(net163),
    .X(_1383_));
 sky130_fd_sc_hd__nor3_2 _4325_ (.A(_2849_),
    .B(_2918_),
    .C(net108),
    .Y(_1384_));
 sky130_fd_sc_hd__o21ai_1 _4326_ (.A1(_0450_),
    .A2(_0666_),
    .B1(_0679_),
    .Y(_1385_));
 sky130_fd_sc_hd__a21o_1 _4327_ (.A1(_2847_),
    .A2(_1385_),
    .B1(_1384_),
    .X(_1386_));
 sky130_fd_sc_hd__or2_1 _4328_ (.A(_0558_),
    .B(_1329_),
    .X(_1387_));
 sky130_fd_sc_hd__a221o_1 _4329_ (.A1(_3041_),
    .A2(_0401_),
    .B1(_1386_),
    .B2(net147),
    .C1(_1387_),
    .X(_1388_));
 sky130_fd_sc_hd__a22o_1 _4330_ (.A1(_0401_),
    .A2(_0422_),
    .B1(_0684_),
    .B2(_2847_),
    .X(_1389_));
 sky130_fd_sc_hd__and3_1 _4331_ (.A(net120),
    .B(_2847_),
    .C(_3026_),
    .X(_1390_));
 sky130_fd_sc_hd__and3_1 _4332_ (.A(_3026_),
    .B(_0405_),
    .C(_0512_),
    .X(_1391_));
 sky130_fd_sc_hd__a221o_1 _4333_ (.A1(_0429_),
    .A2(_0432_),
    .B1(_1390_),
    .B2(net135),
    .C1(_1391_),
    .X(_1392_));
 sky130_fd_sc_hd__a21o_1 _4334_ (.A1(\z80.tv80s.i_tv80_core.i_mcode.MCycle[0] ),
    .A2(_3021_),
    .B1(_1320_),
    .X(_1393_));
 sky130_fd_sc_hd__and3_1 _4335_ (.A(net120),
    .B(net131),
    .C(_2912_),
    .X(_1394_));
 sky130_fd_sc_hd__a211o_1 _4336_ (.A1(net159),
    .A2(_1312_),
    .B1(_1392_),
    .C1(_1394_),
    .X(_1395_));
 sky130_fd_sc_hd__a211o_1 _4337_ (.A1(net147),
    .A2(_1389_),
    .B1(_1395_),
    .C1(net109),
    .X(_1396_));
 sky130_fd_sc_hd__or2_1 _4338_ (.A(net135),
    .B(_0406_),
    .X(_1397_));
 sky130_fd_sc_hd__a31o_1 _4339_ (.A1(net159),
    .A2(net97),
    .A3(_1397_),
    .B1(net108),
    .X(_1398_));
 sky130_fd_sc_hd__o311a_1 _4340_ (.A1(_1315_),
    .A2(_1393_),
    .A3(_1396_),
    .B1(_1398_),
    .C1(net165),
    .X(_1399_));
 sky130_fd_sc_hd__a21oi_1 _4341_ (.A1(net106),
    .A2(_1388_),
    .B1(_1399_),
    .Y(_1400_));
 sky130_fd_sc_hd__a2bb2o_4 _4342_ (.A1_N(net651),
    .A2_N(_1400_),
    .B1(_1383_),
    .B2(net159),
    .X(_1401_));
 sky130_fd_sc_hd__a2111o_1 _4343_ (.A1(_2934_),
    .A2(_0684_),
    .B1(_0749_),
    .C1(_1338_),
    .D1(_1394_),
    .X(_1402_));
 sky130_fd_sc_hd__nand2_1 _4344_ (.A(_3032_),
    .B(_0661_),
    .Y(_1403_));
 sky130_fd_sc_hd__o211a_1 _4345_ (.A1(net135),
    .A2(_1335_),
    .B1(_0422_),
    .C1(net146),
    .X(_1404_));
 sky130_fd_sc_hd__a221o_1 _4346_ (.A1(_2948_),
    .A2(_0401_),
    .B1(_1312_),
    .B2(net157),
    .C1(_1315_),
    .X(_1405_));
 sky130_fd_sc_hd__a41o_1 _4347_ (.A1(net157),
    .A2(_2891_),
    .A3(net109),
    .A4(_1397_),
    .B1(_1404_),
    .X(_1406_));
 sky130_fd_sc_hd__a2111o_1 _4348_ (.A1(_0449_),
    .A2(_1403_),
    .B1(_1405_),
    .C1(_1406_),
    .D1(_1392_),
    .X(_1407_));
 sky130_fd_sc_hd__o31a_1 _4349_ (.A1(_0746_),
    .A2(_1402_),
    .A3(_1407_),
    .B1(net165),
    .X(_1408_));
 sky130_fd_sc_hd__a22o_1 _4350_ (.A1(_3041_),
    .A2(_0461_),
    .B1(_1384_),
    .B2(net146),
    .X(_1409_));
 sky130_fd_sc_hd__a211o_1 _4351_ (.A1(_2934_),
    .A2(_1385_),
    .B1(_1387_),
    .C1(_1409_),
    .X(_1410_));
 sky130_fd_sc_hd__a21oi_1 _4352_ (.A1(net106),
    .A2(_1410_),
    .B1(_1408_),
    .Y(_1411_));
 sky130_fd_sc_hd__a2bb2o_2 _4353_ (.A1_N(\z80.tv80s.i_tv80_core.i_mcode.MCycle[6] ),
    .A2_N(_1411_),
    .B1(_1383_),
    .B2(net157),
    .X(_1412_));
 sky130_fd_sc_hd__or4b_1 _4354_ (.A(net534),
    .B(_0500_),
    .C(_1401_),
    .D_N(_1412_),
    .X(_1413_));
 sky130_fd_sc_hd__mux2_1 _4355_ (.A0(\z80.tv80s.i_tv80_core.XY_State[1] ),
    .A1(net473),
    .S(_1413_),
    .X(_1414_));
 sky130_fd_sc_hd__mux2_1 _4356_ (.A0(net552),
    .A1(_1414_),
    .S(net113),
    .X(_0056_));
 sky130_fd_sc_hd__and3_2 _4357_ (.A(net165),
    .B(_2920_),
    .C(_2921_),
    .X(_1415_));
 sky130_fd_sc_hd__nand2_8 _4358_ (.A(net165),
    .B(_2923_),
    .Y(_1416_));
 sky130_fd_sc_hd__and3_2 _4359_ (.A(net165),
    .B(_2920_),
    .C(_2936_),
    .X(_1417_));
 sky130_fd_sc_hd__nand2_2 _4360_ (.A(net166),
    .B(_2938_),
    .Y(_1418_));
 sky130_fd_sc_hd__or2_1 _4361_ (.A(_1415_),
    .B(_1417_),
    .X(_1419_));
 sky130_fd_sc_hd__a21oi_1 _4362_ (.A1(net103),
    .A2(_1419_),
    .B1(net609),
    .Y(_1420_));
 sky130_fd_sc_hd__or2_1 _4363_ (.A(net609),
    .B(_1419_),
    .X(_1421_));
 sky130_fd_sc_hd__a22o_1 _4364_ (.A1(net473),
    .A2(_1420_),
    .B1(_1421_),
    .B2(net566),
    .X(_1422_));
 sky130_fd_sc_hd__mux2_1 _4365_ (.A0(net597),
    .A1(_1422_),
    .S(net113),
    .X(_0057_));
 sky130_fd_sc_hd__or2_1 _4366_ (.A(net123),
    .B(_1421_),
    .X(_1423_));
 sky130_fd_sc_hd__o22a_1 _4367_ (.A1(net113),
    .A2(net168),
    .B1(_0496_),
    .B2(_1423_),
    .X(_0058_));
 sky130_fd_sc_hd__nor2_4 _4368_ (.A(_0785_),
    .B(_0883_),
    .Y(_1424_));
 sky130_fd_sc_hd__mux2_1 _4369_ (.A0(net503),
    .A1(_0986_),
    .S(_1424_),
    .X(_0059_));
 sky130_fd_sc_hd__mux2_1 _4370_ (.A0(net415),
    .A1(_1028_),
    .S(_1424_),
    .X(_0060_));
 sky130_fd_sc_hd__mux2_1 _4371_ (.A0(net477),
    .A1(_1071_),
    .S(_1424_),
    .X(_0061_));
 sky130_fd_sc_hd__mux2_1 _4372_ (.A0(net394),
    .A1(_1114_),
    .S(_1424_),
    .X(_0062_));
 sky130_fd_sc_hd__mux2_1 _4373_ (.A0(net321),
    .A1(_1156_),
    .S(_1424_),
    .X(_0063_));
 sky130_fd_sc_hd__mux2_1 _4374_ (.A0(net354),
    .A1(_1208_),
    .S(_1424_),
    .X(_0064_));
 sky130_fd_sc_hd__mux2_1 _4375_ (.A0(net331),
    .A1(_1251_),
    .S(_1424_),
    .X(_0065_));
 sky130_fd_sc_hd__mux2_1 _4376_ (.A0(net403),
    .A1(_1308_),
    .S(_1424_),
    .X(_0066_));
 sky130_fd_sc_hd__nor2_4 _4377_ (.A(_0785_),
    .B(_0877_),
    .Y(_1425_));
 sky130_fd_sc_hd__mux2_1 _4378_ (.A0(net383),
    .A1(_0986_),
    .S(_1425_),
    .X(_0067_));
 sky130_fd_sc_hd__mux2_1 _4379_ (.A0(net311),
    .A1(_1028_),
    .S(_1425_),
    .X(_0068_));
 sky130_fd_sc_hd__mux2_1 _4380_ (.A0(net315),
    .A1(_1071_),
    .S(_1425_),
    .X(_0069_));
 sky130_fd_sc_hd__mux2_1 _4381_ (.A0(net393),
    .A1(_1114_),
    .S(_1425_),
    .X(_0070_));
 sky130_fd_sc_hd__mux2_1 _4382_ (.A0(net323),
    .A1(_1156_),
    .S(_1425_),
    .X(_0071_));
 sky130_fd_sc_hd__mux2_1 _4383_ (.A0(net401),
    .A1(_1208_),
    .S(_1425_),
    .X(_0072_));
 sky130_fd_sc_hd__mux2_1 _4384_ (.A0(net334),
    .A1(_1251_),
    .S(_1425_),
    .X(_0073_));
 sky130_fd_sc_hd__mux2_1 _4385_ (.A0(net341),
    .A1(_1308_),
    .S(_1425_),
    .X(_0074_));
 sky130_fd_sc_hd__nor2_1 _4386_ (.A(_3051_),
    .B(_0462_),
    .Y(_1426_));
 sky130_fd_sc_hd__a22o_1 _4387_ (.A1(net166),
    .A2(_1320_),
    .B1(_1426_),
    .B2(net107),
    .X(_1427_));
 sky130_fd_sc_hd__mux2_1 _4388_ (.A0(net526),
    .A1(_1427_),
    .S(net115),
    .X(_0075_));
 sky130_fd_sc_hd__nor2_4 _4389_ (.A(_0785_),
    .B(_0875_),
    .Y(_1428_));
 sky130_fd_sc_hd__mux2_1 _4390_ (.A0(net329),
    .A1(_0986_),
    .S(_1428_),
    .X(_0076_));
 sky130_fd_sc_hd__mux2_1 _4391_ (.A0(net381),
    .A1(_1028_),
    .S(_1428_),
    .X(_0077_));
 sky130_fd_sc_hd__mux2_1 _4392_ (.A0(net313),
    .A1(_1071_),
    .S(_1428_),
    .X(_0078_));
 sky130_fd_sc_hd__mux2_1 _4393_ (.A0(net293),
    .A1(_1114_),
    .S(_1428_),
    .X(_0079_));
 sky130_fd_sc_hd__mux2_1 _4394_ (.A0(net397),
    .A1(_1156_),
    .S(_1428_),
    .X(_0080_));
 sky130_fd_sc_hd__mux2_1 _4395_ (.A0(net325),
    .A1(_1208_),
    .S(_1428_),
    .X(_0081_));
 sky130_fd_sc_hd__mux2_1 _4396_ (.A0(net336),
    .A1(_1251_),
    .S(_1428_),
    .X(_0082_));
 sky130_fd_sc_hd__mux2_1 _4397_ (.A0(net359),
    .A1(_1308_),
    .S(_1428_),
    .X(_0083_));
 sky130_fd_sc_hd__or3b_2 _4398_ (.A(_2873_),
    .B(_0783_),
    .C_N(_0781_),
    .X(_1429_));
 sky130_fd_sc_hd__a31o_4 _4399_ (.A1(_0770_),
    .A2(_0776_),
    .A3(_1429_),
    .B1(net124),
    .X(_1430_));
 sky130_fd_sc_hd__nor2_4 _4400_ (.A(_0883_),
    .B(_1430_),
    .Y(_1431_));
 sky130_fd_sc_hd__nor2_1 _4401_ (.A(_0810_),
    .B(_0963_),
    .Y(_1432_));
 sky130_fd_sc_hd__o221a_1 _4402_ (.A1(\z80.tv80s.i_tv80_core.RegBusA_r[0] ),
    .A2(net85),
    .B1(_0858_),
    .B2(_1432_),
    .C1(_0773_),
    .X(_1433_));
 sky130_fd_sc_hd__mux4_1 _4403_ (.A0(net346),
    .A1(net295),
    .A2(net275),
    .A3(net277),
    .S0(net84),
    .S1(net75),
    .X(_1434_));
 sky130_fd_sc_hd__a21o_2 _4404_ (.A1(_0772_),
    .A2(_1434_),
    .B1(_1433_),
    .X(_1435_));
 sky130_fd_sc_hd__mux2_1 _4405_ (.A0(net285),
    .A1(_1435_),
    .S(_1431_),
    .X(_0084_));
 sky130_fd_sc_hd__or3_1 _4406_ (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][1] ),
    .B(net142),
    .C(_0772_),
    .X(_1436_));
 sky130_fd_sc_hd__o211a_1 _4407_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][1] ),
    .A2(_0981_),
    .B1(net75),
    .C1(_1436_),
    .X(_1437_));
 sky130_fd_sc_hd__mux2_1 _4408_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][1] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][1] ),
    .S(_0981_),
    .X(_1438_));
 sky130_fd_sc_hd__o221a_1 _4409_ (.A1(net283),
    .A2(net142),
    .B1(net84),
    .B2(net299),
    .C1(net75),
    .X(_1439_));
 sky130_fd_sc_hd__o221a_1 _4410_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][1] ),
    .A2(net142),
    .B1(net84),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][1] ),
    .C1(net73),
    .X(_1440_));
 sky130_fd_sc_hd__a211o_1 _4411_ (.A1(net73),
    .A2(_1438_),
    .B1(_1437_),
    .C1(_1299_),
    .X(_1441_));
 sky130_fd_sc_hd__o31a_1 _4412_ (.A1(_1300_),
    .A2(_1439_),
    .A3(_1440_),
    .B1(_1441_),
    .X(_1442_));
 sky130_fd_sc_hd__xnor2_1 _4413_ (.A(_0955_),
    .B(_0964_),
    .Y(_1443_));
 sky130_fd_sc_hd__nor2_1 _4414_ (.A(_0810_),
    .B(_1443_),
    .Y(_1444_));
 sky130_fd_sc_hd__o221a_1 _4415_ (.A1(\z80.tv80s.i_tv80_core.RegBusA_r[1] ),
    .A2(net85),
    .B1(_1016_),
    .B2(_1444_),
    .C1(_0773_),
    .X(_1445_));
 sky130_fd_sc_hd__a21o_2 _4416_ (.A1(net89),
    .A2(_1442_),
    .B1(_1445_),
    .X(_1446_));
 sky130_fd_sc_hd__mux2_1 _4417_ (.A0(net283),
    .A1(_1446_),
    .S(_1431_),
    .X(_0085_));
 sky130_fd_sc_hd__or3_1 _4418_ (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][2] ),
    .B(\z80.tv80s.i_tv80_core.RegAddrB_r[0] ),
    .C(_0772_),
    .X(_1447_));
 sky130_fd_sc_hd__o211a_1 _4419_ (.A1(net409),
    .A2(_0981_),
    .B1(net75),
    .C1(_1447_),
    .X(_1448_));
 sky130_fd_sc_hd__mux2_1 _4420_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][2] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][2] ),
    .S(net84),
    .X(_1449_));
 sky130_fd_sc_hd__o221a_1 _4421_ (.A1(net345),
    .A2(\z80.tv80s.i_tv80_core.RegAddrB_r[0] ),
    .B1(_0981_),
    .B2(net484),
    .C1(net75),
    .X(_1450_));
 sky130_fd_sc_hd__o221a_1 _4422_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][2] ),
    .A2(\z80.tv80s.i_tv80_core.RegAddrB_r[0] ),
    .B1(net84),
    .B2(net492),
    .C1(net73),
    .X(_1451_));
 sky130_fd_sc_hd__a211o_1 _4423_ (.A1(net73),
    .A2(_1449_),
    .B1(_1448_),
    .C1(_1299_),
    .X(_1452_));
 sky130_fd_sc_hd__o31a_1 _4424_ (.A1(_1300_),
    .A2(_1450_),
    .A3(_1451_),
    .B1(_1452_),
    .X(_1453_));
 sky130_fd_sc_hd__nand2_1 _4425_ (.A(_0965_),
    .B(_0967_),
    .Y(_1454_));
 sky130_fd_sc_hd__a31o_1 _4426_ (.A1(net76),
    .A2(_0968_),
    .A3(_1454_),
    .B1(_1068_),
    .X(_1455_));
 sky130_fd_sc_hd__o21a_1 _4427_ (.A1(net249),
    .A2(_0775_),
    .B1(_0773_),
    .X(_1456_));
 sky130_fd_sc_hd__a22o_2 _4428_ (.A1(net89),
    .A2(_1453_),
    .B1(_1455_),
    .B2(_1456_),
    .X(_1457_));
 sky130_fd_sc_hd__mux2_1 _4429_ (.A0(net345),
    .A1(_1457_),
    .S(_1431_),
    .X(_0086_));
 sky130_fd_sc_hd__nor2_1 _4430_ (.A(_0932_),
    .B(_0934_),
    .Y(_1458_));
 sky130_fd_sc_hd__xnor2_1 _4431_ (.A(_0969_),
    .B(_1458_),
    .Y(_1459_));
 sky130_fd_sc_hd__o21bai_1 _4432_ (.A1(_0810_),
    .A2(_1459_),
    .B1_N(_1102_),
    .Y(_1460_));
 sky130_fd_sc_hd__o21a_1 _4433_ (.A1(net253),
    .A2(_0775_),
    .B1(_0773_),
    .X(_1461_));
 sky130_fd_sc_hd__mux4_1 _4434_ (.A0(net423),
    .A1(net301),
    .A2(net343),
    .A3(net371),
    .S0(net75),
    .S1(net84),
    .X(_1462_));
 sky130_fd_sc_hd__a22o_2 _4435_ (.A1(_1460_),
    .A2(_1461_),
    .B1(_1462_),
    .B2(net89),
    .X(_1463_));
 sky130_fd_sc_hd__mux2_1 _4436_ (.A0(net338),
    .A1(_1463_),
    .S(_1431_),
    .X(_0087_));
 sky130_fd_sc_hd__xnor2_1 _4437_ (.A(_0922_),
    .B(_0970_),
    .Y(_1464_));
 sky130_fd_sc_hd__nand2_1 _4438_ (.A(net76),
    .B(_1464_),
    .Y(_1465_));
 sky130_fd_sc_hd__o2bb2a_1 _4439_ (.A1_N(_1152_),
    .A2_N(_1465_),
    .B1(net223),
    .B2(net85),
    .X(_1466_));
 sky130_fd_sc_hd__mux4_2 _4440_ (.A0(net469),
    .A1(net431),
    .A2(net417),
    .A3(net305),
    .S0(net74),
    .S1(net82),
    .X(_1467_));
 sky130_fd_sc_hd__mux2_2 _4441_ (.A0(_1466_),
    .A1(_1467_),
    .S(net89),
    .X(_1468_));
 sky130_fd_sc_hd__mux2_1 _4442_ (.A0(net491),
    .A1(_1468_),
    .S(_1431_),
    .X(_0088_));
 sky130_fd_sc_hd__a21oi_1 _4443_ (.A1(net80),
    .A2(_0921_),
    .B1(_0971_),
    .Y(_1469_));
 sky130_fd_sc_hd__xnor2_1 _4444_ (.A(_0914_),
    .B(_1469_),
    .Y(_1470_));
 sky130_fd_sc_hd__a21o_1 _4445_ (.A1(net76),
    .A2(_1470_),
    .B1(_1193_),
    .X(_1471_));
 sky130_fd_sc_hd__o21a_1 _4446_ (.A1(net247),
    .A2(net85),
    .B1(net86),
    .X(_1472_));
 sky130_fd_sc_hd__mux4_1 _4447_ (.A0(net287),
    .A1(net396),
    .A2(net319),
    .A3(net352),
    .S0(net74),
    .S1(net82),
    .X(_1473_));
 sky130_fd_sc_hd__a22o_2 _4448_ (.A1(_1471_),
    .A2(_1472_),
    .B1(_1473_),
    .B2(net89),
    .X(_1474_));
 sky130_fd_sc_hd__mux2_1 _4449_ (.A0(net483),
    .A1(_1474_),
    .S(_1431_),
    .X(_0089_));
 sky130_fd_sc_hd__o21a_1 _4450_ (.A1(_0972_),
    .A2(_0974_),
    .B1(_0907_),
    .X(_1475_));
 sky130_fd_sc_hd__nor3_1 _4451_ (.A(_0907_),
    .B(_0972_),
    .C(_0974_),
    .Y(_1476_));
 sky130_fd_sc_hd__nor2_1 _4452_ (.A(_1475_),
    .B(_1476_),
    .Y(_1477_));
 sky130_fd_sc_hd__a211o_1 _4453_ (.A1(net76),
    .A2(_1477_),
    .B1(_1247_),
    .C1(_0774_),
    .X(_1478_));
 sky130_fd_sc_hd__o21a_1 _4454_ (.A1(net251),
    .A2(net85),
    .B1(net86),
    .X(_1479_));
 sky130_fd_sc_hd__mux4_1 _4455_ (.A0(net309),
    .A1(net273),
    .A2(net333),
    .A3(net271),
    .S0(net75),
    .S1(net84),
    .X(_1480_));
 sky130_fd_sc_hd__a22o_2 _4456_ (.A1(_1478_),
    .A2(_1479_),
    .B1(_1480_),
    .B2(net89),
    .X(_1481_));
 sky130_fd_sc_hd__mux2_1 _4457_ (.A0(net317),
    .A1(_1481_),
    .S(_1431_),
    .X(_0090_));
 sky130_fd_sc_hd__mux4_1 _4458_ (.A0(net504),
    .A1(net435),
    .A2(net475),
    .A3(net281),
    .S0(net75),
    .S1(net84),
    .X(_1482_));
 sky130_fd_sc_hd__nor2_1 _4459_ (.A(_0906_),
    .B(_1475_),
    .Y(_1483_));
 sky130_fd_sc_hd__xnor2_1 _4460_ (.A(_0898_),
    .B(_1483_),
    .Y(_1484_));
 sky130_fd_sc_hd__a21o_1 _4461_ (.A1(net76),
    .A2(_1484_),
    .B1(_1296_),
    .X(_1485_));
 sky130_fd_sc_hd__o21a_1 _4462_ (.A1(net233),
    .A2(net85),
    .B1(_1485_),
    .X(_1486_));
 sky130_fd_sc_hd__mux2_2 _4463_ (.A0(_1482_),
    .A1(_1486_),
    .S(net86),
    .X(_1487_));
 sky130_fd_sc_hd__mux2_1 _4464_ (.A0(net480),
    .A1(_1487_),
    .S(_1431_),
    .X(_0091_));
 sky130_fd_sc_hd__nor2_4 _4465_ (.A(_0785_),
    .B(_0886_),
    .Y(_1488_));
 sky130_fd_sc_hd__mux2_1 _4466_ (.A0(net488),
    .A1(_0986_),
    .S(_1488_),
    .X(_0092_));
 sky130_fd_sc_hd__mux2_1 _4467_ (.A0(net356),
    .A1(_1028_),
    .S(_1488_),
    .X(_0093_));
 sky130_fd_sc_hd__mux2_1 _4468_ (.A0(net434),
    .A1(_1071_),
    .S(_1488_),
    .X(_0094_));
 sky130_fd_sc_hd__mux2_1 _4469_ (.A0(net456),
    .A1(_1114_),
    .S(_1488_),
    .X(_0095_));
 sky130_fd_sc_hd__mux2_1 _4470_ (.A0(net377),
    .A1(_1156_),
    .S(_1488_),
    .X(_0096_));
 sky130_fd_sc_hd__mux2_1 _4471_ (.A0(net407),
    .A1(_1208_),
    .S(_1488_),
    .X(_0097_));
 sky130_fd_sc_hd__mux2_1 _4472_ (.A0(net327),
    .A1(_1251_),
    .S(_1488_),
    .X(_0098_));
 sky130_fd_sc_hd__mux2_1 _4473_ (.A0(net365),
    .A1(_1308_),
    .S(_1488_),
    .X(_0099_));
 sky130_fd_sc_hd__nor2_4 _4474_ (.A(_0877_),
    .B(_1430_),
    .Y(_1489_));
 sky130_fd_sc_hd__mux2_1 _4475_ (.A0(net275),
    .A1(_1435_),
    .S(_1489_),
    .X(_0100_));
 sky130_fd_sc_hd__mux2_1 _4476_ (.A0(net419),
    .A1(_1446_),
    .S(_1489_),
    .X(_0101_));
 sky130_fd_sc_hd__mux2_1 _4477_ (.A0(net409),
    .A1(_1457_),
    .S(_1489_),
    .X(_0102_));
 sky130_fd_sc_hd__mux2_1 _4478_ (.A0(net301),
    .A1(_1463_),
    .S(_1489_),
    .X(_0103_));
 sky130_fd_sc_hd__mux2_1 _4479_ (.A0(net431),
    .A1(_1468_),
    .S(_1489_),
    .X(_0104_));
 sky130_fd_sc_hd__mux2_1 _4480_ (.A0(net396),
    .A1(_1474_),
    .S(_1489_),
    .X(_0105_));
 sky130_fd_sc_hd__mux2_1 _4481_ (.A0(net273),
    .A1(_1481_),
    .S(_1489_),
    .X(_0106_));
 sky130_fd_sc_hd__mux2_1 _4482_ (.A0(net435),
    .A1(_1487_),
    .S(_1489_),
    .X(_0107_));
 sky130_fd_sc_hd__or2_4 _4483_ (.A(_0785_),
    .B(_0871_),
    .X(_1490_));
 sky130_fd_sc_hd__mux2_1 _4484_ (.A0(_0986_),
    .A1(net496),
    .S(_1490_),
    .X(_0108_));
 sky130_fd_sc_hd__mux2_1 _4485_ (.A0(_1028_),
    .A1(net446),
    .S(_1490_),
    .X(_0109_));
 sky130_fd_sc_hd__mux2_1 _4486_ (.A0(_1071_),
    .A1(net361),
    .S(_1490_),
    .X(_0110_));
 sky130_fd_sc_hd__mux2_1 _4487_ (.A0(_1114_),
    .A1(net367),
    .S(_1490_),
    .X(_0111_));
 sky130_fd_sc_hd__mux2_1 _4488_ (.A0(_1156_),
    .A1(net433),
    .S(_1490_),
    .X(_0112_));
 sky130_fd_sc_hd__mux2_1 _4489_ (.A0(_1208_),
    .A1(net410),
    .S(_1490_),
    .X(_0113_));
 sky130_fd_sc_hd__mux2_1 _4490_ (.A0(_1251_),
    .A1(net358),
    .S(_1490_),
    .X(_0114_));
 sky130_fd_sc_hd__mux2_1 _4491_ (.A0(_1308_),
    .A1(net387),
    .S(_1490_),
    .X(_0115_));
 sky130_fd_sc_hd__or2_4 _4492_ (.A(_0869_),
    .B(_1430_),
    .X(_1491_));
 sky130_fd_sc_hd__mux2_1 _4493_ (.A0(_1435_),
    .A1(net295),
    .S(_1491_),
    .X(_0116_));
 sky130_fd_sc_hd__mux2_1 _4494_ (.A0(_1446_),
    .A1(net391),
    .S(_1491_),
    .X(_0117_));
 sky130_fd_sc_hd__mux2_1 _4495_ (.A0(_1457_),
    .A1(net350),
    .S(_1491_),
    .X(_0118_));
 sky130_fd_sc_hd__mux2_1 _4496_ (.A0(_1463_),
    .A1(net343),
    .S(_1491_),
    .X(_0119_));
 sky130_fd_sc_hd__mux2_1 _4497_ (.A0(_1468_),
    .A1(net417),
    .S(_1491_),
    .X(_0120_));
 sky130_fd_sc_hd__mux2_1 _4498_ (.A0(_1474_),
    .A1(net319),
    .S(_1491_),
    .X(_0121_));
 sky130_fd_sc_hd__mux2_1 _4499_ (.A0(_1481_),
    .A1(net333),
    .S(_1491_),
    .X(_0122_));
 sky130_fd_sc_hd__mux2_1 _4500_ (.A0(_1487_),
    .A1(net475),
    .S(_1491_),
    .X(_0123_));
 sky130_fd_sc_hd__or2_4 _4501_ (.A(_0871_),
    .B(_1430_),
    .X(_1492_));
 sky130_fd_sc_hd__mux2_1 _4502_ (.A0(_1435_),
    .A1(net346),
    .S(_1492_),
    .X(_0124_));
 sky130_fd_sc_hd__mux2_1 _4503_ (.A0(_1446_),
    .A1(net379),
    .S(_1492_),
    .X(_0125_));
 sky130_fd_sc_hd__mux2_1 _4504_ (.A0(_1457_),
    .A1(net444),
    .S(_1492_),
    .X(_0126_));
 sky130_fd_sc_hd__mux2_1 _4505_ (.A0(_1463_),
    .A1(net423),
    .S(_1492_),
    .X(_0127_));
 sky130_fd_sc_hd__mux2_1 _4506_ (.A0(_1468_),
    .A1(net469),
    .S(_1492_),
    .X(_0128_));
 sky130_fd_sc_hd__mux2_1 _4507_ (.A0(_1474_),
    .A1(net287),
    .S(_1492_),
    .X(_0129_));
 sky130_fd_sc_hd__mux2_1 _4508_ (.A0(_1481_),
    .A1(net309),
    .S(_1492_),
    .X(_0130_));
 sky130_fd_sc_hd__mux2_1 _4509_ (.A0(_1487_),
    .A1(net504),
    .S(_1492_),
    .X(_0131_));
 sky130_fd_sc_hd__or2_4 _4510_ (.A(_0785_),
    .B(_0880_),
    .X(_1493_));
 sky130_fd_sc_hd__mux2_1 _4511_ (.A0(_0986_),
    .A1(net511),
    .S(_1493_),
    .X(_0132_));
 sky130_fd_sc_hd__mux2_1 _4512_ (.A0(_1028_),
    .A1(net438),
    .S(_1493_),
    .X(_0133_));
 sky130_fd_sc_hd__mux2_1 _4513_ (.A0(_1071_),
    .A1(net529),
    .S(_1493_),
    .X(_0134_));
 sky130_fd_sc_hd__mux2_1 _4514_ (.A0(_1114_),
    .A1(net414),
    .S(_1493_),
    .X(_0135_));
 sky130_fd_sc_hd__mux2_1 _4515_ (.A0(_1156_),
    .A1(net517),
    .S(_1493_),
    .X(_0136_));
 sky130_fd_sc_hd__mux2_1 _4516_ (.A0(_1208_),
    .A1(net442),
    .S(_1493_),
    .X(_0137_));
 sky130_fd_sc_hd__mux2_1 _4517_ (.A0(_1251_),
    .A1(net460),
    .S(_1493_),
    .X(_0138_));
 sky130_fd_sc_hd__mux2_1 _4518_ (.A0(_1308_),
    .A1(net462),
    .S(_1493_),
    .X(_0139_));
 sky130_fd_sc_hd__or2_4 _4519_ (.A(_0807_),
    .B(_1430_),
    .X(_1494_));
 sky130_fd_sc_hd__mux2_1 _4520_ (.A0(_1435_),
    .A1(net369),
    .S(_1494_),
    .X(_0140_));
 sky130_fd_sc_hd__mux2_1 _4521_ (.A0(_1446_),
    .A1(net512),
    .S(_1494_),
    .X(_0141_));
 sky130_fd_sc_hd__mux2_1 _4522_ (.A0(_1457_),
    .A1(net492),
    .S(_1494_),
    .X(_0142_));
 sky130_fd_sc_hd__mux2_1 _4523_ (.A0(_1463_),
    .A1(net421),
    .S(_1494_),
    .X(_0143_));
 sky130_fd_sc_hd__mux2_1 _4524_ (.A0(_1468_),
    .A1(net482),
    .S(_1494_),
    .X(_0144_));
 sky130_fd_sc_hd__mux2_1 _4525_ (.A0(_1474_),
    .A1(net490),
    .S(_1494_),
    .X(_0145_));
 sky130_fd_sc_hd__mux2_1 _4526_ (.A0(_1481_),
    .A1(net448),
    .S(_1494_),
    .X(_0146_));
 sky130_fd_sc_hd__mux2_1 _4527_ (.A0(_1487_),
    .A1(net510),
    .S(_1494_),
    .X(_0147_));
 sky130_fd_sc_hd__nor2_4 _4528_ (.A(_0875_),
    .B(_1430_),
    .Y(_1495_));
 sky130_fd_sc_hd__mux2_1 _4529_ (.A0(net277),
    .A1(_1435_),
    .S(_1495_),
    .X(_0148_));
 sky130_fd_sc_hd__mux2_1 _4530_ (.A0(net303),
    .A1(_1446_),
    .S(_1495_),
    .X(_0149_));
 sky130_fd_sc_hd__mux2_1 _4531_ (.A0(net289),
    .A1(_1457_),
    .S(_1495_),
    .X(_0150_));
 sky130_fd_sc_hd__mux2_1 _4532_ (.A0(net371),
    .A1(_1463_),
    .S(_1495_),
    .X(_0151_));
 sky130_fd_sc_hd__mux2_1 _4533_ (.A0(net305),
    .A1(_1468_),
    .S(_1495_),
    .X(_0152_));
 sky130_fd_sc_hd__mux2_1 _4534_ (.A0(net352),
    .A1(_1474_),
    .S(_1495_),
    .X(_0153_));
 sky130_fd_sc_hd__mux2_1 _4535_ (.A0(net271),
    .A1(_1481_),
    .S(_1495_),
    .X(_0154_));
 sky130_fd_sc_hd__mux2_1 _4536_ (.A0(net281),
    .A1(_1487_),
    .S(_1495_),
    .X(_0155_));
 sky130_fd_sc_hd__nor2_4 _4537_ (.A(_0886_),
    .B(_1430_),
    .Y(_1496_));
 sky130_fd_sc_hd__mux2_1 _4538_ (.A0(net307),
    .A1(_1435_),
    .S(_1496_),
    .X(_0156_));
 sky130_fd_sc_hd__mux2_1 _4539_ (.A0(net299),
    .A1(_1446_),
    .S(_1496_),
    .X(_0157_));
 sky130_fd_sc_hd__mux2_1 _4540_ (.A0(net484),
    .A1(_1457_),
    .S(_1496_),
    .X(_0158_));
 sky130_fd_sc_hd__mux2_1 _4541_ (.A0(net426),
    .A1(_1463_),
    .S(_1496_),
    .X(_0159_));
 sky130_fd_sc_hd__mux2_1 _4542_ (.A0(net506),
    .A1(_1468_),
    .S(_1496_),
    .X(_0160_));
 sky130_fd_sc_hd__mux2_1 _4543_ (.A0(net485),
    .A1(_1474_),
    .S(_1496_),
    .X(_0161_));
 sky130_fd_sc_hd__mux2_1 _4544_ (.A0(net291),
    .A1(_1481_),
    .S(_1496_),
    .X(_0162_));
 sky130_fd_sc_hd__mux2_1 _4545_ (.A0(net497),
    .A1(_1487_),
    .S(_1496_),
    .X(_0163_));
 sky130_fd_sc_hd__or2_4 _4546_ (.A(_0785_),
    .B(_0869_),
    .X(_1497_));
 sky130_fd_sc_hd__mux2_1 _4547_ (.A0(_0986_),
    .A1(net440),
    .S(_1497_),
    .X(_0164_));
 sky130_fd_sc_hd__mux2_1 _4548_ (.A0(_1028_),
    .A1(net459),
    .S(_1497_),
    .X(_0165_));
 sky130_fd_sc_hd__mux2_1 _4549_ (.A0(_1071_),
    .A1(net427),
    .S(_1497_),
    .X(_0166_));
 sky130_fd_sc_hd__mux2_1 _4550_ (.A0(_1114_),
    .A1(net385),
    .S(_1497_),
    .X(_0167_));
 sky130_fd_sc_hd__mux2_1 _4551_ (.A0(_1156_),
    .A1(net424),
    .S(_1497_),
    .X(_0168_));
 sky130_fd_sc_hd__mux2_1 _4552_ (.A0(_1208_),
    .A1(net428),
    .S(_1497_),
    .X(_0169_));
 sky130_fd_sc_hd__mux2_1 _4553_ (.A0(_1251_),
    .A1(net348),
    .S(_1497_),
    .X(_0170_));
 sky130_fd_sc_hd__mux2_1 _4554_ (.A0(_1308_),
    .A1(net373),
    .S(_1497_),
    .X(_0171_));
 sky130_fd_sc_hd__nand2_2 _4555_ (.A(\z80.tv80s.i_tv80_core.ISet[0] ),
    .B(_2952_),
    .Y(_1498_));
 sky130_fd_sc_hd__and4_4 _4556_ (.A(\z80.tv80s.i_tv80_core.ISet[0] ),
    .B(net116),
    .C(_2952_),
    .D(net94),
    .X(_1499_));
 sky130_fd_sc_hd__nor4_1 _4557_ (.A(net118),
    .B(net110),
    .C(_2899_),
    .D(_2951_),
    .Y(_1500_));
 sky130_fd_sc_hd__inv_2 _4558_ (.A(net92),
    .Y(_1501_));
 sky130_fd_sc_hd__nor2_2 _4559_ (.A(net102),
    .B(_1501_),
    .Y(_1502_));
 sky130_fd_sc_hd__mux2_1 _4560_ (.A0(net686),
    .A1(\z80.tv80s.i_tv80_core.ACC[0] ),
    .S(_1499_),
    .X(_0172_));
 sky130_fd_sc_hd__mux2_1 _4561_ (.A0(net656),
    .A1(\z80.tv80s.i_tv80_core.ACC[1] ),
    .S(_1499_),
    .X(_0173_));
 sky130_fd_sc_hd__mux2_1 _4562_ (.A0(net682),
    .A1(\z80.tv80s.i_tv80_core.ACC[2] ),
    .S(_1499_),
    .X(_0174_));
 sky130_fd_sc_hd__mux2_1 _4563_ (.A0(net696),
    .A1(\z80.tv80s.i_tv80_core.ACC[3] ),
    .S(_1499_),
    .X(_0175_));
 sky130_fd_sc_hd__mux2_1 _4564_ (.A0(net678),
    .A1(\z80.tv80s.i_tv80_core.ACC[4] ),
    .S(_1499_),
    .X(_0176_));
 sky130_fd_sc_hd__mux2_1 _4565_ (.A0(net674),
    .A1(\z80.tv80s.i_tv80_core.ACC[5] ),
    .S(_1499_),
    .X(_0177_));
 sky130_fd_sc_hd__mux2_1 _4566_ (.A0(net658),
    .A1(\z80.tv80s.i_tv80_core.ACC[6] ),
    .S(_1499_),
    .X(_0178_));
 sky130_fd_sc_hd__mux2_1 _4567_ (.A0(net654),
    .A1(\z80.tv80s.i_tv80_core.ACC[7] ),
    .S(_1499_),
    .X(_0179_));
 sky130_fd_sc_hd__mux2_1 _4568_ (.A0(net734),
    .A1(\z80.tv80s.i_tv80_core.F[0] ),
    .S(_1499_),
    .X(_0180_));
 sky130_fd_sc_hd__mux2_1 _4569_ (.A0(net747),
    .A1(\z80.tv80s.i_tv80_core.F[1] ),
    .S(_1499_),
    .X(_0181_));
 sky130_fd_sc_hd__mux2_1 _4570_ (.A0(net668),
    .A1(\z80.tv80s.i_tv80_core.F[2] ),
    .S(_1499_),
    .X(_0182_));
 sky130_fd_sc_hd__mux2_1 _4571_ (.A0(net730),
    .A1(\z80.tv80s.i_tv80_core.F[3] ),
    .S(_1499_),
    .X(_0183_));
 sky130_fd_sc_hd__mux2_1 _4572_ (.A0(net670),
    .A1(\z80.tv80s.i_tv80_core.F[4] ),
    .S(_1499_),
    .X(_0184_));
 sky130_fd_sc_hd__mux2_1 _4573_ (.A0(net705),
    .A1(\z80.tv80s.i_tv80_core.F[5] ),
    .S(_1499_),
    .X(_0185_));
 sky130_fd_sc_hd__mux2_1 _4574_ (.A0(net701),
    .A1(\z80.tv80s.i_tv80_core.F[6] ),
    .S(_1499_),
    .X(_0186_));
 sky130_fd_sc_hd__mux2_1 _4575_ (.A0(net666),
    .A1(\z80.tv80s.i_tv80_core.F[7] ),
    .S(_1499_),
    .X(_0187_));
 sky130_fd_sc_hd__a21o_1 _4576_ (.A1(net96),
    .A2(_1331_),
    .B1(_2999_),
    .X(_1503_));
 sky130_fd_sc_hd__and3_1 _4577_ (.A(_2965_),
    .B(net96),
    .C(_0398_),
    .X(_1504_));
 sky130_fd_sc_hd__a31o_1 _4578_ (.A1(net132),
    .A2(net96),
    .A3(_1334_),
    .B1(_1504_),
    .X(_1505_));
 sky130_fd_sc_hd__a22oi_2 _4579_ (.A1(net107),
    .A2(_1503_),
    .B1(_1505_),
    .B2(\z80.tv80s.i_tv80_core.ISet[0] ),
    .Y(_1506_));
 sky130_fd_sc_hd__a22o_1 _4580_ (.A1(net107),
    .A2(_1503_),
    .B1(_1505_),
    .B2(\z80.tv80s.i_tv80_core.ISet[0] ),
    .X(_1507_));
 sky130_fd_sc_hd__a21oi_1 _4581_ (.A1(_1333_),
    .A2(_1349_),
    .B1(_1506_),
    .Y(_1508_));
 sky130_fd_sc_hd__nor2_2 _4582_ (.A(net125),
    .B(_1508_),
    .Y(_1509_));
 sky130_fd_sc_hd__a31o_1 _4583_ (.A1(net147),
    .A2(net146),
    .A3(net130),
    .B1(net131),
    .X(_1510_));
 sky130_fd_sc_hd__a21bo_1 _4584_ (.A1(net132),
    .A2(net96),
    .B1_N(_1510_),
    .X(_1511_));
 sky130_fd_sc_hd__inv_2 _4585_ (.A(_1511_),
    .Y(_1512_));
 sky130_fd_sc_hd__a221o_1 _4586_ (.A1(_1334_),
    .A2(_1510_),
    .B1(_1512_),
    .B2(_2965_),
    .C1(net109),
    .X(_1513_));
 sky130_fd_sc_hd__o21a_1 _4587_ (.A1(_2920_),
    .A2(_0642_),
    .B1(_2885_),
    .X(_1514_));
 sky130_fd_sc_hd__or2_1 _4588_ (.A(_0488_),
    .B(_1514_),
    .X(_1515_));
 sky130_fd_sc_hd__o21ai_1 _4589_ (.A1(_2963_),
    .A2(_0554_),
    .B1(_0434_),
    .Y(_1516_));
 sky130_fd_sc_hd__a22o_1 _4590_ (.A1(net132),
    .A2(_1515_),
    .B1(_1516_),
    .B2(net150),
    .X(_1517_));
 sky130_fd_sc_hd__a21o_1 _4591_ (.A1(net152),
    .A2(_1343_),
    .B1(_2981_),
    .X(_1518_));
 sky130_fd_sc_hd__o311a_2 _4592_ (.A1(_1317_),
    .A2(_1513_),
    .A3(_1517_),
    .B1(_1518_),
    .C1(net166),
    .X(_1519_));
 sky130_fd_sc_hd__a211o_1 _4593_ (.A1(net152),
    .A2(_1326_),
    .B1(_0448_),
    .C1(_2991_),
    .X(_1520_));
 sky130_fd_sc_hd__nand2_1 _4594_ (.A(\z80.tv80s.i_tv80_core.i_mcode.MCycle[3] ),
    .B(net96),
    .Y(_1521_));
 sky130_fd_sc_hd__or2_1 _4595_ (.A(\z80.tv80s.i_tv80_core.i_mcode.MCycle[3] ),
    .B(net96),
    .X(_1522_));
 sky130_fd_sc_hd__a32o_1 _4596_ (.A1(_1331_),
    .A2(_1521_),
    .A3(_1522_),
    .B1(_1520_),
    .B2(net132),
    .X(_1523_));
 sky130_fd_sc_hd__o21a_1 _4597_ (.A1(_0558_),
    .A2(_1523_),
    .B1(net106),
    .X(_1524_));
 sky130_fd_sc_hd__a211oi_4 _4598_ (.A1(net161),
    .A2(net163),
    .B1(_1519_),
    .C1(_1524_),
    .Y(_1525_));
 sky130_fd_sc_hd__a211o_2 _4599_ (.A1(net161),
    .A2(net163),
    .B1(_1519_),
    .C1(_1524_),
    .X(_1526_));
 sky130_fd_sc_hd__nand2_1 _4600_ (.A(_0888_),
    .B(_1525_),
    .Y(_1527_));
 sky130_fd_sc_hd__nor2_1 _4601_ (.A(_1333_),
    .B(_1349_),
    .Y(_1528_));
 sky130_fd_sc_hd__nor2_2 _4602_ (.A(_1507_),
    .B(_1528_),
    .Y(_1529_));
 sky130_fd_sc_hd__o211a_1 _4603_ (.A1(_0963_),
    .A2(_1525_),
    .B1(_1527_),
    .C1(_1529_),
    .X(_1530_));
 sky130_fd_sc_hd__and4_2 _4604_ (.A(_1333_),
    .B(_1349_),
    .C(_1507_),
    .D(_1525_),
    .X(_1531_));
 sky130_fd_sc_hd__and4_2 _4605_ (.A(_1333_),
    .B(_1349_),
    .C(_1507_),
    .D(_1526_),
    .X(_1532_));
 sky130_fd_sc_hd__and2_2 _4606_ (.A(_1525_),
    .B(_1528_),
    .X(_1533_));
 sky130_fd_sc_hd__and2_2 _4607_ (.A(_1526_),
    .B(_1528_),
    .X(_1534_));
 sky130_fd_sc_hd__a221o_1 _4608_ (.A1(\z80.tv80s.di_reg[0] ),
    .A2(_1533_),
    .B1(_1534_),
    .B2(\z80.tv80s.i_tv80_core.ACC[0] ),
    .C1(_1530_),
    .X(_1535_));
 sky130_fd_sc_hd__a221o_1 _4609_ (.A1(net637),
    .A2(_1531_),
    .B1(_1532_),
    .B2(net664),
    .C1(_1535_),
    .X(_1536_));
 sky130_fd_sc_hd__a22o_1 _4610_ (.A1(net125),
    .A2(net672),
    .B1(_1509_),
    .B2(_1536_),
    .X(_0188_));
 sky130_fd_sc_hd__nand2_1 _4611_ (.A(_0952_),
    .B(_1526_),
    .Y(_1537_));
 sky130_fd_sc_hd__o211a_1 _4612_ (.A1(_1021_),
    .A2(_1526_),
    .B1(_1529_),
    .C1(_1537_),
    .X(_1538_));
 sky130_fd_sc_hd__a221o_1 _4613_ (.A1(\z80.tv80s.di_reg[1] ),
    .A2(_1533_),
    .B1(_1534_),
    .B2(\z80.tv80s.i_tv80_core.ACC[1] ),
    .C1(_1538_),
    .X(_1539_));
 sky130_fd_sc_hd__a221o_1 _4614_ (.A1(net680),
    .A2(_1531_),
    .B1(_1532_),
    .B2(net740),
    .C1(_1539_),
    .X(_1540_));
 sky130_fd_sc_hd__a22o_1 _4615_ (.A1(net126),
    .A2(net784),
    .B1(_1509_),
    .B2(_1540_),
    .X(_0189_));
 sky130_fd_sc_hd__mux2_1 _4616_ (.A0(_0942_),
    .A1(_1034_),
    .S(_1525_),
    .X(_1541_));
 sky130_fd_sc_hd__a22o_1 _4617_ (.A1(\z80.tv80s.di_reg[2] ),
    .A2(_1533_),
    .B1(_1534_),
    .B2(\z80.tv80s.i_tv80_core.ACC[2] ),
    .X(_1542_));
 sky130_fd_sc_hd__a221o_1 _4618_ (.A1(net713),
    .A2(_1531_),
    .B1(_1532_),
    .B2(net583),
    .C1(_1542_),
    .X(_1543_));
 sky130_fd_sc_hd__a21o_1 _4619_ (.A1(_1529_),
    .A2(_1541_),
    .B1(_1543_),
    .X(_1544_));
 sky130_fd_sc_hd__a22o_1 _4620_ (.A1(net126),
    .A2(net749),
    .B1(_1509_),
    .B2(_1544_),
    .X(_0190_));
 sky130_fd_sc_hd__mux2_1 _4621_ (.A0(_0931_),
    .A1(_1107_),
    .S(_1525_),
    .X(_1545_));
 sky130_fd_sc_hd__a22o_1 _4622_ (.A1(\z80.tv80s.di_reg[3] ),
    .A2(_1533_),
    .B1(_1534_),
    .B2(\z80.tv80s.i_tv80_core.ACC[3] ),
    .X(_1546_));
 sky130_fd_sc_hd__a221o_1 _4623_ (.A1(\z80.tv80s.i_tv80_core.SP[3] ),
    .A2(_1531_),
    .B1(_1532_),
    .B2(\z80.tv80s.i_tv80_core.SP[11] ),
    .C1(_1546_),
    .X(_1547_));
 sky130_fd_sc_hd__a21o_1 _4624_ (.A1(_1529_),
    .A2(_1545_),
    .B1(_1547_),
    .X(_1548_));
 sky130_fd_sc_hd__a22o_1 _4625_ (.A1(net125),
    .A2(net690),
    .B1(_1509_),
    .B2(_1548_),
    .X(_0191_));
 sky130_fd_sc_hd__mux2_1 _4626_ (.A0(_0921_),
    .A1(_1122_),
    .S(_1525_),
    .X(_1549_));
 sky130_fd_sc_hd__a22o_1 _4627_ (.A1(\z80.tv80s.di_reg[4] ),
    .A2(_1533_),
    .B1(_1534_),
    .B2(\z80.tv80s.i_tv80_core.ACC[4] ),
    .X(_1550_));
 sky130_fd_sc_hd__a221o_1 _4628_ (.A1(net662),
    .A2(_1531_),
    .B1(_1532_),
    .B2(\z80.tv80s.i_tv80_core.SP[12] ),
    .C1(_1550_),
    .X(_1551_));
 sky130_fd_sc_hd__a21o_1 _4629_ (.A1(_1529_),
    .A2(_1549_),
    .B1(_1551_),
    .X(_1552_));
 sky130_fd_sc_hd__a22o_1 _4630_ (.A1(net126),
    .A2(net707),
    .B1(_1509_),
    .B2(_1552_),
    .X(_0192_));
 sky130_fd_sc_hd__mux2_1 _4631_ (.A0(_0913_),
    .A1(_1198_),
    .S(_1525_),
    .X(_1553_));
 sky130_fd_sc_hd__a22o_1 _4632_ (.A1(\z80.tv80s.di_reg[5] ),
    .A2(_1533_),
    .B1(_1534_),
    .B2(\z80.tv80s.i_tv80_core.ACC[5] ),
    .X(_1554_));
 sky130_fd_sc_hd__a221o_1 _4633_ (.A1(net718),
    .A2(_1531_),
    .B1(_1532_),
    .B2(net688),
    .C1(_1554_),
    .X(_1555_));
 sky130_fd_sc_hd__a21o_1 _4634_ (.A1(_1529_),
    .A2(_1553_),
    .B1(_1555_),
    .X(_1556_));
 sky130_fd_sc_hd__a22o_1 _4635_ (.A1(net126),
    .A2(net726),
    .B1(_1509_),
    .B2(_1556_),
    .X(_0193_));
 sky130_fd_sc_hd__or2_1 _4636_ (.A(_0905_),
    .B(_1525_),
    .X(_1557_));
 sky130_fd_sc_hd__o211a_1 _4637_ (.A1(_1213_),
    .A2(_1526_),
    .B1(_1529_),
    .C1(_1557_),
    .X(_1558_));
 sky130_fd_sc_hd__a221o_1 _4638_ (.A1(\z80.tv80s.di_reg[6] ),
    .A2(_1533_),
    .B1(_1534_),
    .B2(\z80.tv80s.i_tv80_core.ACC[6] ),
    .C1(_1558_),
    .X(_1559_));
 sky130_fd_sc_hd__a221o_1 _4639_ (.A1(net660),
    .A2(_1531_),
    .B1(_1532_),
    .B2(\z80.tv80s.i_tv80_core.SP[14] ),
    .C1(_1559_),
    .X(_1560_));
 sky130_fd_sc_hd__a22o_1 _4640_ (.A1(net126),
    .A2(net768),
    .B1(_1509_),
    .B2(_1560_),
    .X(_0194_));
 sky130_fd_sc_hd__or2_1 _4641_ (.A(_0897_),
    .B(_1525_),
    .X(_1561_));
 sky130_fd_sc_hd__o211a_1 _4642_ (.A1(_1257_),
    .A2(_1526_),
    .B1(_1529_),
    .C1(_1561_),
    .X(_1562_));
 sky130_fd_sc_hd__a221o_1 _4643_ (.A1(net848),
    .A2(_1533_),
    .B1(_1534_),
    .B2(net849),
    .C1(_1562_),
    .X(_1563_));
 sky130_fd_sc_hd__a221o_1 _4644_ (.A1(net798),
    .A2(_1531_),
    .B1(_1532_),
    .B2(net814),
    .C1(_1563_),
    .X(_1564_));
 sky130_fd_sc_hd__a22o_1 _4645_ (.A1(net126),
    .A2(net162),
    .B1(_1509_),
    .B2(_1564_),
    .X(_0195_));
 sky130_fd_sc_hd__and2b_1 _4646_ (.A_N(net14),
    .B(\z80.tv80s.i_tv80_core.Oldnmi_n ),
    .X(_1565_));
 sky130_fd_sc_hd__o21ba_1 _4647_ (.A1(net518),
    .A2(_1565_),
    .B1_N(net621),
    .X(_0196_));
 sky130_fd_sc_hd__a211o_1 _4648_ (.A1(net778),
    .A2(net585),
    .B1(net711),
    .C1(net621),
    .X(_1566_));
 sky130_fd_sc_hd__nand2_2 _4649_ (.A(net101),
    .B(_1566_),
    .Y(_1567_));
 sky130_fd_sc_hd__and2_1 _4650_ (.A(net13),
    .B(_1567_),
    .X(_1568_));
 sky130_fd_sc_hd__a21o_1 _4651_ (.A1(net129),
    .A2(net163),
    .B1(net101),
    .X(_1569_));
 sky130_fd_sc_hd__and3_4 _4652_ (.A(net113),
    .B(_0603_),
    .C(_1569_),
    .X(_1570_));
 sky130_fd_sc_hd__nand2_1 _4653_ (.A(net778),
    .B(net269),
    .Y(_1571_));
 sky130_fd_sc_hd__o21ai_4 _4654_ (.A1(net94),
    .A2(_1571_),
    .B1(_1570_),
    .Y(_1572_));
 sky130_fd_sc_hd__o22a_1 _4655_ (.A1(net160),
    .A2(_1570_),
    .B1(_1572_),
    .B2(_1568_),
    .X(_0197_));
 sky130_fd_sc_hd__and2_1 _4656_ (.A(net12),
    .B(_1567_),
    .X(_1573_));
 sky130_fd_sc_hd__o22a_1 _4657_ (.A1(net159),
    .A2(_1570_),
    .B1(_1572_),
    .B2(_1573_),
    .X(_0198_));
 sky130_fd_sc_hd__and2_1 _4658_ (.A(net10),
    .B(_1567_),
    .X(_1574_));
 sky130_fd_sc_hd__o22a_1 _4659_ (.A1(net156),
    .A2(_1570_),
    .B1(_1572_),
    .B2(_1574_),
    .X(_0199_));
 sky130_fd_sc_hd__and2_1 _4660_ (.A(net7),
    .B(_1567_),
    .X(_1575_));
 sky130_fd_sc_hd__o22a_1 _4661_ (.A1(net153),
    .A2(_1570_),
    .B1(_1572_),
    .B2(_1575_),
    .X(_0200_));
 sky130_fd_sc_hd__and2_1 _4662_ (.A(net6),
    .B(_1567_),
    .X(_1576_));
 sky130_fd_sc_hd__o22a_1 _4663_ (.A1(net148),
    .A2(_1570_),
    .B1(_1572_),
    .B2(_1576_),
    .X(_0201_));
 sky130_fd_sc_hd__and2_1 _4664_ (.A(net8),
    .B(_1567_),
    .X(_1577_));
 sky130_fd_sc_hd__o22a_1 _4665_ (.A1(net144),
    .A2(_1570_),
    .B1(_1572_),
    .B2(_1577_),
    .X(_0202_));
 sky130_fd_sc_hd__and2_1 _4666_ (.A(net9),
    .B(_1567_),
    .X(_1578_));
 sky130_fd_sc_hd__o22a_1 _4667_ (.A1(net835),
    .A2(_1570_),
    .B1(_1572_),
    .B2(_1578_),
    .X(_0203_));
 sky130_fd_sc_hd__and2_1 _4668_ (.A(net11),
    .B(_1567_),
    .X(_1579_));
 sky130_fd_sc_hd__o22a_1 _4669_ (.A1(net845),
    .A2(_1570_),
    .B1(_1572_),
    .B2(_1579_),
    .X(_0204_));
 sky130_fd_sc_hd__and4_2 _4670_ (.A(_2874_),
    .B(net720),
    .C(_0781_),
    .D(_0782_),
    .X(_1580_));
 sky130_fd_sc_hd__nand2_8 _4671_ (.A(_2873_),
    .B(_1580_),
    .Y(_1581_));
 sky130_fd_sc_hd__a21oi_4 _4672_ (.A1(_0779_),
    .A2(_1581_),
    .B1(net127),
    .Y(_1582_));
 sky130_fd_sc_hd__nor2_1 _4673_ (.A(_0856_),
    .B(_1581_),
    .Y(_1583_));
 sky130_fd_sc_hd__nor2_1 _4674_ (.A(net105),
    .B(_0554_),
    .Y(_1584_));
 sky130_fd_sc_hd__or3_4 _4675_ (.A(net152),
    .B(net105),
    .C(_0667_),
    .X(_1585_));
 sky130_fd_sc_hd__and2_4 _4676_ (.A(_0676_),
    .B(_1584_),
    .X(_1586_));
 sky130_fd_sc_hd__mux2_1 _4677_ (.A0(\z80.tv80s.i_tv80_core.BusB[0] ),
    .A1(\z80.tv80s.i_tv80_core.BusA[0] ),
    .S(_1586_),
    .X(_1587_));
 sky130_fd_sc_hd__mux2_1 _4678_ (.A0(\z80.tv80s.i_tv80_core.BusB[4] ),
    .A1(_1587_),
    .S(_1585_),
    .X(_1588_));
 sky130_fd_sc_hd__o21a_1 _4679_ (.A1(_0779_),
    .A2(_1588_),
    .B1(_1581_),
    .X(_1589_));
 sky130_fd_sc_hd__o32a_1 _4680_ (.A1(net127),
    .A2(_1583_),
    .A3(_1589_),
    .B1(net530),
    .B2(_1582_),
    .X(_0205_));
 sky130_fd_sc_hd__nor2_1 _4681_ (.A(_1014_),
    .B(_1581_),
    .Y(_1590_));
 sky130_fd_sc_hd__mux2_1 _4682_ (.A0(\z80.tv80s.i_tv80_core.BusB[1] ),
    .A1(\z80.tv80s.i_tv80_core.BusA[1] ),
    .S(_1586_),
    .X(_1591_));
 sky130_fd_sc_hd__mux2_1 _4683_ (.A0(\z80.tv80s.i_tv80_core.BusB[5] ),
    .A1(_1591_),
    .S(_1585_),
    .X(_1592_));
 sky130_fd_sc_hd__o21a_1 _4684_ (.A1(_0779_),
    .A2(_1592_),
    .B1(_1581_),
    .X(_1593_));
 sky130_fd_sc_hd__o32a_1 _4685_ (.A1(net127),
    .A2(_1590_),
    .A3(_1593_),
    .B1(net554),
    .B2(_1582_),
    .X(_0206_));
 sky130_fd_sc_hd__mux2_1 _4686_ (.A0(\z80.tv80s.i_tv80_core.BusB[2] ),
    .A1(\z80.tv80s.i_tv80_core.BusA[2] ),
    .S(_1586_),
    .X(_1594_));
 sky130_fd_sc_hd__mux2_1 _4687_ (.A0(\z80.tv80s.i_tv80_core.BusB[6] ),
    .A1(_1594_),
    .S(_1585_),
    .X(_1595_));
 sky130_fd_sc_hd__nor2_1 _4688_ (.A(_1066_),
    .B(_1581_),
    .Y(_1596_));
 sky130_fd_sc_hd__o21a_1 _4689_ (.A1(_0779_),
    .A2(_1595_),
    .B1(_1581_),
    .X(_1597_));
 sky130_fd_sc_hd__o32a_1 _4690_ (.A1(net127),
    .A2(_1596_),
    .A3(_1597_),
    .B1(net546),
    .B2(_1582_),
    .X(_0207_));
 sky130_fd_sc_hd__nor2_1 _4691_ (.A(_1100_),
    .B(_1581_),
    .Y(_1598_));
 sky130_fd_sc_hd__mux2_1 _4692_ (.A0(\z80.tv80s.i_tv80_core.BusB[3] ),
    .A1(\z80.tv80s.i_tv80_core.BusA[3] ),
    .S(_1586_),
    .X(_1599_));
 sky130_fd_sc_hd__mux2_1 _4693_ (.A0(\z80.tv80s.i_tv80_core.BusB[7] ),
    .A1(_1599_),
    .S(_1585_),
    .X(_1600_));
 sky130_fd_sc_hd__o21a_1 _4694_ (.A1(_0779_),
    .A2(_1600_),
    .B1(_1581_),
    .X(_1601_));
 sky130_fd_sc_hd__o32a_1 _4695_ (.A1(net127),
    .A2(_1598_),
    .A3(_1601_),
    .B1(net536),
    .B2(_1582_),
    .X(_0208_));
 sky130_fd_sc_hd__nor2_1 _4696_ (.A(_1150_),
    .B(_1581_),
    .Y(_1602_));
 sky130_fd_sc_hd__mux2_1 _4697_ (.A0(\z80.tv80s.i_tv80_core.BusB[4] ),
    .A1(\z80.tv80s.i_tv80_core.BusB[0] ),
    .S(_1586_),
    .X(_1603_));
 sky130_fd_sc_hd__mux2_1 _4698_ (.A0(\z80.tv80s.i_tv80_core.BusA[0] ),
    .A1(_1603_),
    .S(_1585_),
    .X(_1604_));
 sky130_fd_sc_hd__o21a_1 _4699_ (.A1(_0779_),
    .A2(_1604_),
    .B1(_1581_),
    .X(_1605_));
 sky130_fd_sc_hd__o32a_1 _4700_ (.A1(net127),
    .A2(_1602_),
    .A3(_1605_),
    .B1(net540),
    .B2(_1582_),
    .X(_0209_));
 sky130_fd_sc_hd__nor2_1 _4701_ (.A(_1191_),
    .B(_1581_),
    .Y(_1606_));
 sky130_fd_sc_hd__mux2_1 _4702_ (.A0(\z80.tv80s.i_tv80_core.BusB[5] ),
    .A1(\z80.tv80s.i_tv80_core.BusB[1] ),
    .S(_1586_),
    .X(_1607_));
 sky130_fd_sc_hd__mux2_1 _4703_ (.A0(\z80.tv80s.i_tv80_core.BusA[1] ),
    .A1(_1607_),
    .S(_1585_),
    .X(_1608_));
 sky130_fd_sc_hd__o21a_1 _4704_ (.A1(_0779_),
    .A2(_1608_),
    .B1(_1581_),
    .X(_1609_));
 sky130_fd_sc_hd__o32a_1 _4705_ (.A1(net127),
    .A2(_1606_),
    .A3(_1609_),
    .B1(net538),
    .B2(_1582_),
    .X(_0210_));
 sky130_fd_sc_hd__nor2_1 _4706_ (.A(_1245_),
    .B(_1581_),
    .Y(_1610_));
 sky130_fd_sc_hd__mux2_1 _4707_ (.A0(\z80.tv80s.i_tv80_core.BusB[6] ),
    .A1(\z80.tv80s.i_tv80_core.BusB[2] ),
    .S(_1586_),
    .X(_1611_));
 sky130_fd_sc_hd__mux2_1 _4708_ (.A0(\z80.tv80s.i_tv80_core.BusA[2] ),
    .A1(_1611_),
    .S(_1585_),
    .X(_1612_));
 sky130_fd_sc_hd__o21a_1 _4709_ (.A1(_0779_),
    .A2(_1612_),
    .B1(_1581_),
    .X(_1613_));
 sky130_fd_sc_hd__o32a_1 _4710_ (.A1(net127),
    .A2(_1610_),
    .A3(_1613_),
    .B1(net532),
    .B2(_1582_),
    .X(_0211_));
 sky130_fd_sc_hd__mux2_1 _4711_ (.A0(\z80.tv80s.i_tv80_core.BusB[7] ),
    .A1(\z80.tv80s.i_tv80_core.BusB[3] ),
    .S(_1586_),
    .X(_1614_));
 sky130_fd_sc_hd__mux2_1 _4712_ (.A0(\z80.tv80s.i_tv80_core.BusA[3] ),
    .A1(_1614_),
    .S(_1585_),
    .X(_1615_));
 sky130_fd_sc_hd__or2_1 _4713_ (.A(_0779_),
    .B(_1615_),
    .X(_1616_));
 sky130_fd_sc_hd__mux2_1 _4714_ (.A0(_1295_),
    .A1(_1616_),
    .S(_1581_),
    .X(_1617_));
 sky130_fd_sc_hd__o22a_1 _4715_ (.A1(net550),
    .A2(_1582_),
    .B1(_1617_),
    .B2(net127),
    .X(_0212_));
 sky130_fd_sc_hd__and4_2 _4716_ (.A(net154),
    .B(_2846_),
    .C(\z80.tv80s.i_tv80_core.ISet[0] ),
    .D(_2929_),
    .X(_1618_));
 sky130_fd_sc_hd__nand2_1 _4717_ (.A(_0577_),
    .B(_1618_),
    .Y(_1619_));
 sky130_fd_sc_hd__a21o_2 _4718_ (.A1(_1498_),
    .A2(_1619_),
    .B1(net102),
    .X(_1620_));
 sky130_fd_sc_hd__inv_2 _4719_ (.A(_1620_),
    .Y(_1621_));
 sky130_fd_sc_hd__or4_4 _4720_ (.A(net119),
    .B(_2930_),
    .C(_0469_),
    .D(net60),
    .X(_1622_));
 sky130_fd_sc_hd__o22a_1 _4721_ (.A1(net686),
    .A2(_1501_),
    .B1(_1622_),
    .B2(_2876_),
    .X(_1623_));
 sky130_fd_sc_hd__o22a_1 _4722_ (.A1(\z80.tv80s.i_tv80_core.ACC[0] ),
    .A2(_1621_),
    .B1(_1623_),
    .B2(net102),
    .X(_1624_));
 sky130_fd_sc_hd__or3b_1 _4723_ (.A(_2846_),
    .B(_2854_),
    .C_N(_1354_),
    .X(_1625_));
 sky130_fd_sc_hd__and3_4 _4724_ (.A(net147),
    .B(\z80.tv80s.i_tv80_core.ts[3] ),
    .C(_1354_),
    .X(_1626_));
 sky130_fd_sc_hd__nand2_4 _4725_ (.A(net633),
    .B(_1580_),
    .Y(_1627_));
 sky130_fd_sc_hd__mux2_1 _4726_ (.A0(net581),
    .A1(net558),
    .S(_1355_),
    .X(_1628_));
 sky130_fd_sc_hd__mux2_1 _4727_ (.A0(_1624_),
    .A1(_1628_),
    .S(_1626_),
    .X(_1629_));
 sky130_fd_sc_hd__mux2_1 _4728_ (.A0(_0857_),
    .A1(_1629_),
    .S(_1627_),
    .X(_1630_));
 sky130_fd_sc_hd__mux2_1 _4729_ (.A0(net852),
    .A1(_1630_),
    .S(net115),
    .X(_0213_));
 sky130_fd_sc_hd__a2bb2o_1 _4730_ (.A1_N(\z80.tv80s.i_tv80_core.ACC[1] ),
    .A2_N(_1622_),
    .B1(net91),
    .B2(net656),
    .X(_1631_));
 sky130_fd_sc_hd__a22o_1 _4731_ (.A1(\z80.tv80s.i_tv80_core.ACC[1] ),
    .A2(_1620_),
    .B1(_1631_),
    .B2(net94),
    .X(_1632_));
 sky130_fd_sc_hd__mux2_1 _4732_ (.A0(net676),
    .A1(net615),
    .S(_1355_),
    .X(_1633_));
 sky130_fd_sc_hd__mux2_1 _4733_ (.A0(_1632_),
    .A1(_1633_),
    .S(_1626_),
    .X(_1634_));
 sky130_fd_sc_hd__mux2_1 _4734_ (.A0(_1015_),
    .A1(_1634_),
    .S(_1627_),
    .X(_1635_));
 sky130_fd_sc_hd__mux2_1 _4735_ (.A0(net850),
    .A1(_1635_),
    .S(net115),
    .X(_0214_));
 sky130_fd_sc_hd__a2bb2o_1 _4736_ (.A1_N(\z80.tv80s.i_tv80_core.ACC[2] ),
    .A2_N(_1622_),
    .B1(net92),
    .B2(net682),
    .X(_1636_));
 sky130_fd_sc_hd__a22o_1 _4737_ (.A1(\z80.tv80s.i_tv80_core.ACC[2] ),
    .A2(_1620_),
    .B1(_1636_),
    .B2(net94),
    .X(_1637_));
 sky130_fd_sc_hd__mux2_1 _4738_ (.A0(net623),
    .A1(net544),
    .S(_1355_),
    .X(_1638_));
 sky130_fd_sc_hd__mux2_1 _4739_ (.A0(_1637_),
    .A1(_1638_),
    .S(_1626_),
    .X(_1639_));
 sky130_fd_sc_hd__mux2_1 _4740_ (.A0(_1067_),
    .A1(_1639_),
    .S(_1627_),
    .X(_1640_));
 sky130_fd_sc_hd__mux2_1 _4741_ (.A0(net855),
    .A1(_1640_),
    .S(net115),
    .X(_0215_));
 sky130_fd_sc_hd__a2bb2o_1 _4742_ (.A1_N(\z80.tv80s.i_tv80_core.ACC[3] ),
    .A2_N(_1622_),
    .B1(net91),
    .B2(net696),
    .X(_1641_));
 sky130_fd_sc_hd__a22o_1 _4743_ (.A1(\z80.tv80s.i_tv80_core.ACC[3] ),
    .A2(_1620_),
    .B1(_1641_),
    .B2(net94),
    .X(_1642_));
 sky130_fd_sc_hd__mux2_1 _4744_ (.A0(net627),
    .A1(net527),
    .S(_1355_),
    .X(_1643_));
 sky130_fd_sc_hd__mux2_1 _4745_ (.A0(_1642_),
    .A1(_1643_),
    .S(_1626_),
    .X(_1644_));
 sky130_fd_sc_hd__mux2_1 _4746_ (.A0(_1101_),
    .A1(_1644_),
    .S(_1627_),
    .X(_1645_));
 sky130_fd_sc_hd__mux2_1 _4747_ (.A0(net862),
    .A1(_1645_),
    .S(net115),
    .X(_0216_));
 sky130_fd_sc_hd__a2bb2o_1 _4748_ (.A1_N(\z80.tv80s.i_tv80_core.ACC[4] ),
    .A2_N(_1622_),
    .B1(net92),
    .B2(net678),
    .X(_1646_));
 sky130_fd_sc_hd__a22o_1 _4749_ (.A1(\z80.tv80s.i_tv80_core.ACC[4] ),
    .A2(_1620_),
    .B1(_1646_),
    .B2(net94),
    .X(_1647_));
 sky130_fd_sc_hd__mux2_1 _4750_ (.A0(net579),
    .A1(net613),
    .S(_1355_),
    .X(_1648_));
 sky130_fd_sc_hd__mux2_1 _4751_ (.A0(_1647_),
    .A1(_1648_),
    .S(_1626_),
    .X(_1649_));
 sky130_fd_sc_hd__mux2_1 _4752_ (.A0(_1151_),
    .A1(_1649_),
    .S(_1627_),
    .X(_1650_));
 sky130_fd_sc_hd__mux2_1 _4753_ (.A0(net851),
    .A1(_1650_),
    .S(net115),
    .X(_0217_));
 sky130_fd_sc_hd__a2bb2o_1 _4754_ (.A1_N(\z80.tv80s.i_tv80_core.ACC[5] ),
    .A2_N(_1622_),
    .B1(net91),
    .B2(net674),
    .X(_1651_));
 sky130_fd_sc_hd__a22o_1 _4755_ (.A1(\z80.tv80s.i_tv80_core.ACC[5] ),
    .A2(_1620_),
    .B1(_1651_),
    .B2(net94),
    .X(_1652_));
 sky130_fd_sc_hd__mux2_1 _4756_ (.A0(net722),
    .A1(net564),
    .S(_1355_),
    .X(_1653_));
 sky130_fd_sc_hd__mux2_1 _4757_ (.A0(_1652_),
    .A1(_1653_),
    .S(_1626_),
    .X(_1654_));
 sky130_fd_sc_hd__mux2_1 _4758_ (.A0(_1192_),
    .A1(_1654_),
    .S(_1627_),
    .X(_1655_));
 sky130_fd_sc_hd__mux2_1 _4759_ (.A0(net859),
    .A1(_1655_),
    .S(net115),
    .X(_0218_));
 sky130_fd_sc_hd__a2bb2o_1 _4760_ (.A1_N(\z80.tv80s.i_tv80_core.ACC[6] ),
    .A2_N(_1622_),
    .B1(net91),
    .B2(\z80.tv80s.i_tv80_core.Ap[6] ),
    .X(_1656_));
 sky130_fd_sc_hd__a22o_1 _4761_ (.A1(\z80.tv80s.i_tv80_core.ACC[6] ),
    .A2(_1620_),
    .B1(_1656_),
    .B2(net94),
    .X(_1657_));
 sky130_fd_sc_hd__mux2_1 _4762_ (.A0(net732),
    .A1(net684),
    .S(_1355_),
    .X(_1658_));
 sky130_fd_sc_hd__mux2_1 _4763_ (.A0(_1657_),
    .A1(_1658_),
    .S(_1626_),
    .X(_1659_));
 sky130_fd_sc_hd__mux2_1 _4764_ (.A0(_1246_),
    .A1(_1659_),
    .S(_1627_),
    .X(_1660_));
 sky130_fd_sc_hd__mux2_1 _4765_ (.A0(net857),
    .A1(_1660_),
    .S(net115),
    .X(_0219_));
 sky130_fd_sc_hd__a2bb2o_1 _4766_ (.A1_N(\z80.tv80s.i_tv80_core.ACC[7] ),
    .A2_N(_1622_),
    .B1(net91),
    .B2(net654),
    .X(_1661_));
 sky130_fd_sc_hd__a22o_1 _4767_ (.A1(\z80.tv80s.i_tv80_core.ACC[7] ),
    .A2(_1620_),
    .B1(_1661_),
    .B2(net94),
    .X(_1662_));
 sky130_fd_sc_hd__mux2_1 _4768_ (.A0(net792),
    .A1(net494),
    .S(_1355_),
    .X(_1663_));
 sky130_fd_sc_hd__mux2_1 _4769_ (.A0(_1662_),
    .A1(_1663_),
    .S(_1626_),
    .X(_1664_));
 sky130_fd_sc_hd__mux2_1 _4770_ (.A0(_1295_),
    .A1(_1664_),
    .S(_1627_),
    .X(_1665_));
 sky130_fd_sc_hd__mux2_1 _4771_ (.A0(net849),
    .A1(_1665_),
    .S(net115),
    .X(_0220_));
 sky130_fd_sc_hd__o21ai_2 _4772_ (.A1(_0577_),
    .A2(_0598_),
    .B1(_0605_),
    .Y(_1666_));
 sky130_fd_sc_hd__a22o_1 _4773_ (.A1(net130),
    .A2(_2917_),
    .B1(_0425_),
    .B2(_0652_),
    .X(_1667_));
 sky130_fd_sc_hd__a221oi_4 _4774_ (.A1(_0415_),
    .A2(_0514_),
    .B1(_0623_),
    .B2(_0861_),
    .C1(_1667_),
    .Y(_1668_));
 sky130_fd_sc_hd__o21a_4 _4775_ (.A1(net119),
    .A2(_1668_),
    .B1(_0728_),
    .X(_1669_));
 sky130_fd_sc_hd__o21ai_2 _4776_ (.A1(net119),
    .A2(_1668_),
    .B1(_0728_),
    .Y(_1670_));
 sky130_fd_sc_hd__mux4_1 _4777_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][0] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][0] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][0] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][0] ),
    .S0(net168),
    .S1(net139),
    .X(_1671_));
 sky130_fd_sc_hd__mux4_1 _4778_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][0] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][0] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][0] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][0] ),
    .S0(net168),
    .S1(net139),
    .X(_1672_));
 sky130_fd_sc_hd__mux2_4 _4779_ (.A0(_1672_),
    .A1(_1671_),
    .S(net597),
    .X(_1673_));
 sky130_fd_sc_hd__o21a_1 _4780_ (.A1(net88),
    .A2(_1673_),
    .B1(net79),
    .X(_1674_));
 sky130_fd_sc_hd__a2111o_1 _4781_ (.A1(_2899_),
    .A2(_2949_),
    .B1(_0416_),
    .C1(_0706_),
    .D1(_2912_),
    .X(_1675_));
 sky130_fd_sc_hd__and3_1 _4782_ (.A(net159),
    .B(net156),
    .C(\z80.tv80s.i_tv80_core.IR[7] ),
    .X(_1676_));
 sky130_fd_sc_hd__or4b_2 _4783_ (.A(net118),
    .B(_0653_),
    .C(_1675_),
    .D_N(_1676_),
    .X(_1677_));
 sky130_fd_sc_hd__or4_1 _4784_ (.A(_2948_),
    .B(_2949_),
    .C(_3022_),
    .D(_0433_),
    .X(_1678_));
 sky130_fd_sc_hd__or3_1 _4785_ (.A(_0419_),
    .B(_1319_),
    .C(_1678_),
    .X(_1679_));
 sky130_fd_sc_hd__or4_2 _4786_ (.A(net118),
    .B(_0699_),
    .C(_0860_),
    .D(_1679_),
    .X(_1680_));
 sky130_fd_sc_hd__nand2_2 _4787_ (.A(_1677_),
    .B(_1680_),
    .Y(_1681_));
 sky130_fd_sc_hd__and2_2 _4788_ (.A(\z80.tv80s.i_tv80_core.NMICycle ),
    .B(_0717_),
    .X(_1682_));
 sky130_fd_sc_hd__nor2_1 _4789_ (.A(net68),
    .B(_1682_),
    .Y(_1683_));
 sky130_fd_sc_hd__and3_2 _4790_ (.A(\z80.tv80s.i_tv80_core.i_mcode.MCycle[2] ),
    .B(\z80.tv80s.i_tv80_core.IntCycle ),
    .C(\z80.tv80s.i_tv80_core.IStatus[1] ),
    .X(_1684_));
 sky130_fd_sc_hd__nand3_2 _4791_ (.A(\z80.tv80s.i_tv80_core.i_mcode.MCycle[2] ),
    .B(\z80.tv80s.i_tv80_core.IntCycle ),
    .C(\z80.tv80s.i_tv80_core.IStatus[1] ),
    .Y(_1685_));
 sky130_fd_sc_hd__or3b_4 _4792_ (.A(_2894_),
    .B(_0458_),
    .C_N(_0496_),
    .X(_1686_));
 sky130_fd_sc_hd__inv_4 _4793_ (.A(_1686_),
    .Y(_1687_));
 sky130_fd_sc_hd__nor3b_2 _4794_ (.A(_0496_),
    .B(_0458_),
    .C_N(_0447_),
    .Y(_1688_));
 sky130_fd_sc_hd__or2_4 _4795_ (.A(_0447_),
    .B(_0496_),
    .X(_1689_));
 sky130_fd_sc_hd__clkinv_4 _4796_ (.A(_1689_),
    .Y(_1690_));
 sky130_fd_sc_hd__and3b_4 _4797_ (.A_N(_0496_),
    .B(_0447_),
    .C(_0458_),
    .X(_1691_));
 sky130_fd_sc_hd__a22o_1 _4798_ (.A1(_1673_),
    .A2(_1690_),
    .B1(_1691_),
    .B2(\z80.tv80s.di_reg[0] ),
    .X(_1692_));
 sky130_fd_sc_hd__a21o_1 _4799_ (.A1(\z80.tv80s.i_tv80_core.SP[0] ),
    .A2(_1688_),
    .B1(_1692_),
    .X(_1693_));
 sky130_fd_sc_hd__mux2_1 _4800_ (.A0(\z80.tv80s.i_tv80_core.TmpAddr[0] ),
    .A1(\z80.tv80s.i_tv80_core.PC[0] ),
    .S(_0502_),
    .X(_1694_));
 sky130_fd_sc_hd__mux2_1 _4801_ (.A0(_1673_),
    .A1(_1694_),
    .S(net103),
    .X(_1695_));
 sky130_fd_sc_hd__and4_4 _4802_ (.A(_2895_),
    .B(_0447_),
    .C(_0458_),
    .D(_0496_),
    .X(_1696_));
 sky130_fd_sc_hd__nor2_1 _4803_ (.A(_0703_),
    .B(_1675_),
    .Y(_1697_));
 sky130_fd_sc_hd__and4bb_1 _4804_ (.A_N(net118),
    .B_N(_0554_),
    .C(_0696_),
    .D(_2967_),
    .X(_1698_));
 sky130_fd_sc_hd__nor2_1 _4805_ (.A(_2947_),
    .B(_0697_),
    .Y(_1699_));
 sky130_fd_sc_hd__and4_1 _4806_ (.A(_0694_),
    .B(_1697_),
    .C(_1698_),
    .D(_1699_),
    .X(_1700_));
 sky130_fd_sc_hd__a21o_4 _4807_ (.A1(_0390_),
    .A2(_1584_),
    .B1(_1700_),
    .X(_1701_));
 sky130_fd_sc_hd__inv_2 _4808_ (.A(_1701_),
    .Y(_1702_));
 sky130_fd_sc_hd__nand2_1 _4809_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[0] ),
    .B(_1701_),
    .Y(_1703_));
 sky130_fd_sc_hd__or2_1 _4810_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[0] ),
    .B(_1701_),
    .X(_1704_));
 sky130_fd_sc_hd__a32o_1 _4811_ (.A1(_1696_),
    .A2(_1703_),
    .A3(_1704_),
    .B1(_1695_),
    .B2(net61),
    .X(_1705_));
 sky130_fd_sc_hd__a211o_1 _4812_ (.A1(\z80.tv80s.i_tv80_core.PC[0] ),
    .A2(_1687_),
    .B1(_1693_),
    .C1(_1705_),
    .X(_1706_));
 sky130_fd_sc_hd__mux2_1 _4813_ (.A0(\z80.tv80s.i_tv80_core.TmpAddr[0] ),
    .A1(_1706_),
    .S(net99),
    .X(_1707_));
 sky130_fd_sc_hd__a221o_1 _4814_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[0] ),
    .A2(net68),
    .B1(net66),
    .B2(_1707_),
    .C1(net90),
    .X(_1708_));
 sky130_fd_sc_hd__a221o_1 _4815_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[0] ),
    .A2(net78),
    .B1(_1674_),
    .B2(_1708_),
    .C1(net102),
    .X(_1709_));
 sky130_fd_sc_hd__o21ba_1 _4816_ (.A1(net558),
    .A2(net93),
    .B1_N(net59),
    .X(_1710_));
 sky130_fd_sc_hd__a22o_1 _4817_ (.A1(net569),
    .A2(net59),
    .B1(_1709_),
    .B2(_1710_),
    .X(_0221_));
 sky130_fd_sc_hd__a21o_1 _4818_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[1] ),
    .A2(_1684_),
    .B1(_1682_),
    .X(_1711_));
 sky130_fd_sc_hd__mux4_1 _4819_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][1] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][1] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][1] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][1] ),
    .S0(net168),
    .S1(net139),
    .X(_1712_));
 sky130_fd_sc_hd__nand2b_1 _4820_ (.A_N(_1712_),
    .B(net597),
    .Y(_1713_));
 sky130_fd_sc_hd__mux4_2 _4821_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][1] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][1] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][1] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][1] ),
    .S0(net168),
    .S1(net139),
    .X(_1714_));
 sky130_fd_sc_hd__o21a_1 _4822_ (.A1(net597),
    .A2(_1714_),
    .B1(_1713_),
    .X(_1715_));
 sky130_fd_sc_hd__o21ai_2 _4823_ (.A1(net169),
    .A2(_1714_),
    .B1(_1713_),
    .Y(_1716_));
 sky130_fd_sc_hd__nor2_1 _4824_ (.A(_1689_),
    .B(_1716_),
    .Y(_1717_));
 sky130_fd_sc_hd__a221o_1 _4825_ (.A1(\z80.tv80s.i_tv80_core.SP[1] ),
    .A2(_1688_),
    .B1(_1691_),
    .B2(\z80.tv80s.di_reg[1] ),
    .C1(_1717_),
    .X(_1718_));
 sky130_fd_sc_hd__mux2_1 _4826_ (.A0(\z80.tv80s.i_tv80_core.PC[1] ),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[1] ),
    .S(net140),
    .X(_1719_));
 sky130_fd_sc_hd__mux2_1 _4827_ (.A0(_1715_),
    .A1(_1719_),
    .S(net103),
    .X(_1720_));
 sky130_fd_sc_hd__and3_1 _4828_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[0] ),
    .B(\z80.tv80s.i_tv80_core.TmpAddr[1] ),
    .C(_1701_),
    .X(_1721_));
 sky130_fd_sc_hd__a21oi_1 _4829_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[0] ),
    .A2(_1701_),
    .B1(\z80.tv80s.i_tv80_core.TmpAddr[1] ),
    .Y(_1722_));
 sky130_fd_sc_hd__nor2_1 _4830_ (.A(_1721_),
    .B(_1722_),
    .Y(_1723_));
 sky130_fd_sc_hd__a22o_1 _4831_ (.A1(net61),
    .A2(_1720_),
    .B1(_1723_),
    .B2(_1696_),
    .X(_1724_));
 sky130_fd_sc_hd__a211o_1 _4832_ (.A1(\z80.tv80s.i_tv80_core.PC[1] ),
    .A2(_1687_),
    .B1(_1718_),
    .C1(_1724_),
    .X(_1725_));
 sky130_fd_sc_hd__a21o_1 _4833_ (.A1(net99),
    .A2(_1725_),
    .B1(_1711_),
    .X(_1726_));
 sky130_fd_sc_hd__mux2_1 _4834_ (.A0(_1726_),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[1] ),
    .S(net68),
    .X(_1727_));
 sky130_fd_sc_hd__nor2_1 _4835_ (.A(net88),
    .B(_1716_),
    .Y(_1728_));
 sky130_fd_sc_hd__a211o_1 _4836_ (.A1(net88),
    .A2(_1727_),
    .B1(_1728_),
    .C1(net78),
    .X(_1729_));
 sky130_fd_sc_hd__or2_1 _4837_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[1] ),
    .B(_1669_),
    .X(_1730_));
 sky130_fd_sc_hd__and2_1 _4838_ (.A(\z80.tv80s.i_tv80_core.R[1] ),
    .B(net102),
    .X(_1731_));
 sky130_fd_sc_hd__a31o_1 _4839_ (.A1(net94),
    .A2(_1729_),
    .A3(_1730_),
    .B1(_1731_),
    .X(_1732_));
 sky130_fd_sc_hd__mux2_1 _4840_ (.A0(_1732_),
    .A1(net587),
    .S(net59),
    .X(_0222_));
 sky130_fd_sc_hd__a21o_1 _4841_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[2] ),
    .A2(_1684_),
    .B1(_1682_),
    .X(_1733_));
 sky130_fd_sc_hd__mux4_1 _4842_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][2] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][2] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][2] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][2] ),
    .S0(net139),
    .S1(net168),
    .X(_1734_));
 sky130_fd_sc_hd__mux4_1 _4843_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][2] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][2] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][2] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][2] ),
    .S0(net139),
    .S1(net168),
    .X(_1735_));
 sky130_fd_sc_hd__mux2_2 _4844_ (.A0(_1735_),
    .A1(_1734_),
    .S(net169),
    .X(_1736_));
 sky130_fd_sc_hd__mux2_1 _4845_ (.A0(\z80.tv80s.i_tv80_core.PC[2] ),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[2] ),
    .S(net140),
    .X(_1737_));
 sky130_fd_sc_hd__mux2_1 _4846_ (.A0(_1736_),
    .A1(_1737_),
    .S(net103),
    .X(_1738_));
 sky130_fd_sc_hd__and2_1 _4847_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[2] ),
    .B(_1721_),
    .X(_1739_));
 sky130_fd_sc_hd__a221o_1 _4848_ (.A1(\z80.tv80s.i_tv80_core.SP[2] ),
    .A2(_1688_),
    .B1(_1690_),
    .B2(_1736_),
    .C1(_1687_),
    .X(_1740_));
 sky130_fd_sc_hd__o21ai_1 _4849_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[2] ),
    .A2(_1721_),
    .B1(_1696_),
    .Y(_1741_));
 sky130_fd_sc_hd__nor2_1 _4850_ (.A(_1739_),
    .B(_1741_),
    .Y(_1742_));
 sky130_fd_sc_hd__a22o_1 _4851_ (.A1(\z80.tv80s.di_reg[2] ),
    .A2(_1691_),
    .B1(_1738_),
    .B2(net61),
    .X(_1743_));
 sky130_fd_sc_hd__or3_1 _4852_ (.A(_1740_),
    .B(_1742_),
    .C(_1743_),
    .X(_1744_));
 sky130_fd_sc_hd__or2_1 _4853_ (.A(\z80.tv80s.i_tv80_core.PC[2] ),
    .B(_1686_),
    .X(_1745_));
 sky130_fd_sc_hd__a31o_1 _4854_ (.A1(net99),
    .A2(_1744_),
    .A3(_1745_),
    .B1(_1733_),
    .X(_1746_));
 sky130_fd_sc_hd__mux2_1 _4855_ (.A0(_1746_),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[2] ),
    .S(net68),
    .X(_1747_));
 sky130_fd_sc_hd__nand2_1 _4856_ (.A(net88),
    .B(_1747_),
    .Y(_1748_));
 sky130_fd_sc_hd__a21oi_1 _4857_ (.A1(_1417_),
    .A2(_1736_),
    .B1(_1670_),
    .Y(_1749_));
 sky130_fd_sc_hd__a221o_1 _4858_ (.A1(_2880_),
    .A2(net78),
    .B1(_1748_),
    .B2(_1749_),
    .C1(net102),
    .X(_1750_));
 sky130_fd_sc_hd__o21ai_1 _4859_ (.A1(_2877_),
    .A2(net94),
    .B1(_1750_),
    .Y(_1751_));
 sky130_fd_sc_hd__mux2_1 _4860_ (.A0(_1751_),
    .A1(net560),
    .S(net59),
    .X(_0223_));
 sky130_fd_sc_hd__mux4_1 _4861_ (.A0(net371),
    .A1(net301),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][3] ),
    .A3(net426),
    .S0(net139),
    .S1(net168),
    .X(_1752_));
 sky130_fd_sc_hd__mux4_1 _4862_ (.A0(net343),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][3] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][3] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][3] ),
    .S0(net139),
    .S1(net168),
    .X(_1753_));
 sky130_fd_sc_hd__mux2_2 _4863_ (.A0(_1753_),
    .A1(_1752_),
    .S(net169),
    .X(_1754_));
 sky130_fd_sc_hd__a21o_1 _4864_ (.A1(net90),
    .A2(_1754_),
    .B1(_1670_),
    .X(_1755_));
 sky130_fd_sc_hd__nand2_1 _4865_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[3] ),
    .B(_1739_),
    .Y(_1756_));
 sky130_fd_sc_hd__or2_1 _4866_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[3] ),
    .B(_1739_),
    .X(_1757_));
 sky130_fd_sc_hd__and3_1 _4867_ (.A(_1696_),
    .B(_1756_),
    .C(_1757_),
    .X(_1758_));
 sky130_fd_sc_hd__mux2_1 _4868_ (.A0(\z80.tv80s.i_tv80_core.PC[3] ),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[3] ),
    .S(net140),
    .X(_1759_));
 sky130_fd_sc_hd__mux2_1 _4869_ (.A0(_1754_),
    .A1(_1759_),
    .S(net103),
    .X(_1760_));
 sky130_fd_sc_hd__a221o_1 _4870_ (.A1(\z80.tv80s.i_tv80_core.SP[3] ),
    .A2(_1688_),
    .B1(_1690_),
    .B2(_1754_),
    .C1(_1687_),
    .X(_1761_));
 sky130_fd_sc_hd__a221o_1 _4871_ (.A1(\z80.tv80s.di_reg[3] ),
    .A2(_1691_),
    .B1(_1760_),
    .B2(_0498_),
    .C1(_1758_),
    .X(_1762_));
 sky130_fd_sc_hd__o22a_1 _4872_ (.A1(\z80.tv80s.i_tv80_core.PC[3] ),
    .A2(_1686_),
    .B1(_1761_),
    .B2(_1762_),
    .X(_1763_));
 sky130_fd_sc_hd__mux2_1 _4873_ (.A0(\z80.tv80s.i_tv80_core.TmpAddr[3] ),
    .A1(_1763_),
    .S(net99),
    .X(_1764_));
 sky130_fd_sc_hd__a22o_1 _4874_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[3] ),
    .A2(net68),
    .B1(net66),
    .B2(_1764_),
    .X(_1765_));
 sky130_fd_sc_hd__a21o_1 _4875_ (.A1(net88),
    .A2(_1765_),
    .B1(_1755_),
    .X(_1766_));
 sky130_fd_sc_hd__o21a_1 _4876_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[3] ),
    .A2(_1669_),
    .B1(net93),
    .X(_1767_));
 sky130_fd_sc_hd__a22o_1 _4877_ (.A1(net527),
    .A2(net102),
    .B1(_1766_),
    .B2(_1767_),
    .X(_1768_));
 sky130_fd_sc_hd__mux2_1 _4878_ (.A0(_1768_),
    .A1(net575),
    .S(net59),
    .X(_0224_));
 sky130_fd_sc_hd__mux4_1 _4879_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][4] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][4] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][4] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][4] ),
    .S0(net138),
    .S1(net167),
    .X(_1769_));
 sky130_fd_sc_hd__mux4_1 _4880_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][4] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][4] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][4] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][4] ),
    .S0(net138),
    .S1(net167),
    .X(_1770_));
 sky130_fd_sc_hd__mux2_4 _4881_ (.A0(_1770_),
    .A1(_1769_),
    .S(net169),
    .X(_1771_));
 sky130_fd_sc_hd__a21o_1 _4882_ (.A1(_1417_),
    .A2(_1771_),
    .B1(net78),
    .X(_1772_));
 sky130_fd_sc_hd__and3_1 _4883_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[3] ),
    .B(\z80.tv80s.i_tv80_core.TmpAddr[4] ),
    .C(_1739_),
    .X(_1773_));
 sky130_fd_sc_hd__a31o_1 _4884_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[2] ),
    .A2(\z80.tv80s.i_tv80_core.TmpAddr[3] ),
    .A3(_1721_),
    .B1(\z80.tv80s.i_tv80_core.TmpAddr[4] ),
    .X(_1774_));
 sky130_fd_sc_hd__and3b_1 _4885_ (.A_N(_1773_),
    .B(_1774_),
    .C(_1696_),
    .X(_1775_));
 sky130_fd_sc_hd__mux2_1 _4886_ (.A0(\z80.tv80s.i_tv80_core.PC[4] ),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[4] ),
    .S(net140),
    .X(_1776_));
 sky130_fd_sc_hd__mux2_1 _4887_ (.A0(_1771_),
    .A1(_1776_),
    .S(net103),
    .X(_1777_));
 sky130_fd_sc_hd__a221o_1 _4888_ (.A1(\z80.tv80s.i_tv80_core.SP[4] ),
    .A2(net62),
    .B1(_1690_),
    .B2(_1771_),
    .C1(_1687_),
    .X(_1778_));
 sky130_fd_sc_hd__a22o_1 _4889_ (.A1(\z80.tv80s.di_reg[4] ),
    .A2(_1691_),
    .B1(_1777_),
    .B2(net61),
    .X(_1779_));
 sky130_fd_sc_hd__or2_1 _4890_ (.A(\z80.tv80s.i_tv80_core.PC[4] ),
    .B(_1686_),
    .X(_1780_));
 sky130_fd_sc_hd__o31a_1 _4891_ (.A1(_1775_),
    .A2(_1778_),
    .A3(_1779_),
    .B1(_1780_),
    .X(_1781_));
 sky130_fd_sc_hd__mux2_1 _4892_ (.A0(\z80.tv80s.i_tv80_core.TmpAddr[4] ),
    .A1(_1781_),
    .S(net99),
    .X(_1782_));
 sky130_fd_sc_hd__a22o_1 _4893_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[4] ),
    .A2(_1681_),
    .B1(net66),
    .B2(_1782_),
    .X(_1783_));
 sky130_fd_sc_hd__a21o_1 _4894_ (.A1(net88),
    .A2(_1783_),
    .B1(_1772_),
    .X(_1784_));
 sky130_fd_sc_hd__o21a_1 _4895_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[4] ),
    .A2(_1669_),
    .B1(net93),
    .X(_1785_));
 sky130_fd_sc_hd__a22o_1 _4896_ (.A1(\z80.tv80s.i_tv80_core.R[4] ),
    .A2(net102),
    .B1(_1784_),
    .B2(_1785_),
    .X(_1786_));
 sky130_fd_sc_hd__mux2_1 _4897_ (.A0(_1786_),
    .A1(net591),
    .S(net59),
    .X(_0225_));
 sky130_fd_sc_hd__mux4_1 _4898_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][5] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][5] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][5] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][5] ),
    .S0(net138),
    .S1(net167),
    .X(_1787_));
 sky130_fd_sc_hd__mux4_1 _4899_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][5] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][5] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][5] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][5] ),
    .S0(net138),
    .S1(net167),
    .X(_1788_));
 sky130_fd_sc_hd__mux2_2 _4900_ (.A0(_1788_),
    .A1(_1787_),
    .S(net169),
    .X(_1789_));
 sky130_fd_sc_hd__nand2_1 _4901_ (.A(net90),
    .B(_1789_),
    .Y(_1790_));
 sky130_fd_sc_hd__a21o_1 _4902_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[5] ),
    .A2(_1684_),
    .B1(_1682_),
    .X(_1791_));
 sky130_fd_sc_hd__mux2_1 _4903_ (.A0(\z80.tv80s.i_tv80_core.PC[5] ),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[5] ),
    .S(net140),
    .X(_1792_));
 sky130_fd_sc_hd__mux2_1 _4904_ (.A0(_1789_),
    .A1(_1792_),
    .S(net103),
    .X(_1793_));
 sky130_fd_sc_hd__nand2_1 _4905_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[5] ),
    .B(_1773_),
    .Y(_1794_));
 sky130_fd_sc_hd__a221o_1 _4906_ (.A1(\z80.tv80s.i_tv80_core.SP[5] ),
    .A2(net62),
    .B1(_1690_),
    .B2(_1789_),
    .C1(_1687_),
    .X(_1795_));
 sky130_fd_sc_hd__o21a_1 _4907_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[5] ),
    .A2(_1773_),
    .B1(_1696_),
    .X(_1796_));
 sky130_fd_sc_hd__a22o_1 _4908_ (.A1(\z80.tv80s.di_reg[5] ),
    .A2(_1691_),
    .B1(_1793_),
    .B2(net61),
    .X(_1797_));
 sky130_fd_sc_hd__a211o_1 _4909_ (.A1(_1794_),
    .A2(_1796_),
    .B1(_1797_),
    .C1(_1795_),
    .X(_1798_));
 sky130_fd_sc_hd__or2_1 _4910_ (.A(\z80.tv80s.i_tv80_core.PC[5] ),
    .B(_1686_),
    .X(_1799_));
 sky130_fd_sc_hd__a31o_1 _4911_ (.A1(net98),
    .A2(_1798_),
    .A3(_1799_),
    .B1(_1791_),
    .X(_1800_));
 sky130_fd_sc_hd__mux2_1 _4912_ (.A0(_1800_),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[5] ),
    .S(net67),
    .X(_1801_));
 sky130_fd_sc_hd__a21bo_1 _4913_ (.A1(net88),
    .A2(_1801_),
    .B1_N(_1790_),
    .X(_1802_));
 sky130_fd_sc_hd__mux2_1 _4914_ (.A0(\z80.tv80s.i_tv80_core.TmpAddr[5] ),
    .A1(_1802_),
    .S(_1669_),
    .X(_1803_));
 sky130_fd_sc_hd__mux2_1 _4915_ (.A0(net564),
    .A1(_1803_),
    .S(net95),
    .X(_1804_));
 sky130_fd_sc_hd__mux2_1 _4916_ (.A0(_1804_),
    .A1(net571),
    .S(net59),
    .X(_0226_));
 sky130_fd_sc_hd__mux4_1 _4917_ (.A0(net271),
    .A1(net273),
    .A2(net317),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][6] ),
    .S0(\z80.tv80s.i_tv80_core.RegAddrC[0] ),
    .S1(\z80.tv80s.i_tv80_core.RegAddrC[1] ),
    .X(_1805_));
 sky130_fd_sc_hd__mux4_1 _4918_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][6] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][6] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][6] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][6] ),
    .S0(\z80.tv80s.i_tv80_core.RegAddrC[0] ),
    .S1(\z80.tv80s.i_tv80_core.RegAddrC[1] ),
    .X(_1806_));
 sky130_fd_sc_hd__mux2_2 _4919_ (.A0(_1806_),
    .A1(_1805_),
    .S(net597),
    .X(_1807_));
 sky130_fd_sc_hd__and2_1 _4920_ (.A(net90),
    .B(_1807_),
    .X(_1808_));
 sky130_fd_sc_hd__a21o_1 _4921_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[6] ),
    .A2(_1684_),
    .B1(_1682_),
    .X(_1809_));
 sky130_fd_sc_hd__and3_1 _4922_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[5] ),
    .B(\z80.tv80s.i_tv80_core.TmpAddr[6] ),
    .C(_1773_),
    .X(_1810_));
 sky130_fd_sc_hd__a21o_1 _4923_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[5] ),
    .A2(_1773_),
    .B1(\z80.tv80s.i_tv80_core.TmpAddr[6] ),
    .X(_1811_));
 sky130_fd_sc_hd__and3b_1 _4924_ (.A_N(_1810_),
    .B(_1811_),
    .C(_1696_),
    .X(_1812_));
 sky130_fd_sc_hd__mux2_1 _4925_ (.A0(\z80.tv80s.i_tv80_core.PC[6] ),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[6] ),
    .S(net140),
    .X(_1813_));
 sky130_fd_sc_hd__mux2_1 _4926_ (.A0(_1807_),
    .A1(_1813_),
    .S(net103),
    .X(_1814_));
 sky130_fd_sc_hd__a221o_1 _4927_ (.A1(\z80.tv80s.i_tv80_core.SP[6] ),
    .A2(net62),
    .B1(_1690_),
    .B2(_1807_),
    .C1(_1687_),
    .X(_1815_));
 sky130_fd_sc_hd__a22o_1 _4928_ (.A1(\z80.tv80s.di_reg[6] ),
    .A2(_1691_),
    .B1(_1814_),
    .B2(net61),
    .X(_1816_));
 sky130_fd_sc_hd__or3_1 _4929_ (.A(_1812_),
    .B(_1815_),
    .C(_1816_),
    .X(_1817_));
 sky130_fd_sc_hd__or2_1 _4930_ (.A(\z80.tv80s.i_tv80_core.PC[6] ),
    .B(_1686_),
    .X(_1818_));
 sky130_fd_sc_hd__a31o_1 _4931_ (.A1(net99),
    .A2(_1817_),
    .A3(_1818_),
    .B1(_1809_),
    .X(_1819_));
 sky130_fd_sc_hd__mux2_1 _4932_ (.A0(_1819_),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[6] ),
    .S(net68),
    .X(_1820_));
 sky130_fd_sc_hd__a21o_1 _4933_ (.A1(net88),
    .A2(_1820_),
    .B1(_1808_),
    .X(_1821_));
 sky130_fd_sc_hd__mux2_1 _4934_ (.A0(\z80.tv80s.i_tv80_core.TmpAddr[6] ),
    .A1(_1821_),
    .S(_1669_),
    .X(_1822_));
 sky130_fd_sc_hd__mux2_1 _4935_ (.A0(\z80.tv80s.i_tv80_core.R[6] ),
    .A1(_1822_),
    .S(net95),
    .X(_1823_));
 sky130_fd_sc_hd__mux2_1 _4936_ (.A0(_1823_),
    .A1(net601),
    .S(net59),
    .X(_0227_));
 sky130_fd_sc_hd__mux4_1 _4937_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][7] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][7] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][7] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][7] ),
    .S0(net139),
    .S1(net168),
    .X(_1824_));
 sky130_fd_sc_hd__nand2b_1 _4938_ (.A_N(_1824_),
    .B(net169),
    .Y(_1825_));
 sky130_fd_sc_hd__mux4_2 _4939_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][7] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][7] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][7] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][7] ),
    .S0(net139),
    .S1(net168),
    .X(_1826_));
 sky130_fd_sc_hd__o21ai_4 _4940_ (.A1(net169),
    .A2(_1826_),
    .B1(_1825_),
    .Y(_1827_));
 sky130_fd_sc_hd__inv_2 _4941_ (.A(_1827_),
    .Y(_1828_));
 sky130_fd_sc_hd__nand2_1 _4942_ (.A(net90),
    .B(_1828_),
    .Y(_1829_));
 sky130_fd_sc_hd__and4_1 _4943_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[4] ),
    .B(\z80.tv80s.i_tv80_core.TmpAddr[5] ),
    .C(\z80.tv80s.i_tv80_core.TmpAddr[6] ),
    .D(\z80.tv80s.i_tv80_core.TmpAddr[7] ),
    .X(_1830_));
 sky130_fd_sc_hd__and4_1 _4944_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[0] ),
    .B(\z80.tv80s.i_tv80_core.TmpAddr[1] ),
    .C(\z80.tv80s.i_tv80_core.TmpAddr[2] ),
    .D(\z80.tv80s.i_tv80_core.TmpAddr[3] ),
    .X(_1831_));
 sky130_fd_sc_hd__nand2_1 _4945_ (.A(_1830_),
    .B(_1831_),
    .Y(_1832_));
 sky130_fd_sc_hd__o221a_1 _4946_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[7] ),
    .A2(_1810_),
    .B1(_1832_),
    .B2(_1702_),
    .C1(_1696_),
    .X(_1833_));
 sky130_fd_sc_hd__mux2_1 _4947_ (.A0(\z80.tv80s.i_tv80_core.PC[7] ),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[7] ),
    .S(net140),
    .X(_1834_));
 sky130_fd_sc_hd__mux2_1 _4948_ (.A0(_1828_),
    .A1(_1834_),
    .S(net103),
    .X(_1835_));
 sky130_fd_sc_hd__nor2_1 _4949_ (.A(_1689_),
    .B(_1827_),
    .Y(_1836_));
 sky130_fd_sc_hd__a221o_1 _4950_ (.A1(\z80.tv80s.i_tv80_core.SP[7] ),
    .A2(net62),
    .B1(_1691_),
    .B2(\z80.tv80s.di_reg[7] ),
    .C1(_1836_),
    .X(_1837_));
 sky130_fd_sc_hd__a21o_1 _4951_ (.A1(net61),
    .A2(_1835_),
    .B1(_1837_),
    .X(_1838_));
 sky130_fd_sc_hd__a211o_1 _4952_ (.A1(\z80.tv80s.i_tv80_core.PC[7] ),
    .A2(_1687_),
    .B1(_1833_),
    .C1(_1838_),
    .X(_1839_));
 sky130_fd_sc_hd__mux2_1 _4953_ (.A0(\z80.tv80s.i_tv80_core.TmpAddr[7] ),
    .A1(_1839_),
    .S(net99),
    .X(_1840_));
 sky130_fd_sc_hd__a22o_1 _4954_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[7] ),
    .A2(net68),
    .B1(net66),
    .B2(_1840_),
    .X(_1841_));
 sky130_fd_sc_hd__a21bo_1 _4955_ (.A1(net87),
    .A2(_1841_),
    .B1_N(_1829_),
    .X(_1842_));
 sky130_fd_sc_hd__mux2_1 _4956_ (.A0(\z80.tv80s.i_tv80_core.TmpAddr[7] ),
    .A1(_1842_),
    .S(net79),
    .X(_1843_));
 sky130_fd_sc_hd__mux2_1 _4957_ (.A0(net494),
    .A1(_1843_),
    .S(net94),
    .X(_1844_));
 sky130_fd_sc_hd__mux2_1 _4958_ (.A0(_1844_),
    .A1(net603),
    .S(net59),
    .X(_0228_));
 sky130_fd_sc_hd__mux4_1 _4959_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][0] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][0] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][0] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][0] ),
    .S0(net167),
    .S1(net138),
    .X(_1845_));
 sky130_fd_sc_hd__mux4_1 _4960_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][0] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][0] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][0] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][0] ),
    .S0(net167),
    .S1(net138),
    .X(_1846_));
 sky130_fd_sc_hd__mux2_2 _4961_ (.A0(_1846_),
    .A1(_1845_),
    .S(net169),
    .X(_1847_));
 sky130_fd_sc_hd__nand2_1 _4962_ (.A(net90),
    .B(_1847_),
    .Y(_1848_));
 sky130_fd_sc_hd__and2_1 _4963_ (.A(\z80.tv80s.i_tv80_core.ACC[0] ),
    .B(_1691_),
    .X(_1849_));
 sky130_fd_sc_hd__a221o_1 _4964_ (.A1(\z80.tv80s.i_tv80_core.SP[8] ),
    .A2(net62),
    .B1(_1690_),
    .B2(_1847_),
    .C1(_1849_),
    .X(_1850_));
 sky130_fd_sc_hd__mux2_1 _4965_ (.A0(\z80.tv80s.i_tv80_core.PC[8] ),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[8] ),
    .S(net140),
    .X(_1851_));
 sky130_fd_sc_hd__mux2_1 _4966_ (.A0(_1847_),
    .A1(_1851_),
    .S(net104),
    .X(_1852_));
 sky130_fd_sc_hd__nor2_1 _4967_ (.A(_2881_),
    .B(_1832_),
    .Y(_1853_));
 sky130_fd_sc_hd__and2_1 _4968_ (.A(_2881_),
    .B(_1832_),
    .X(_1854_));
 sky130_fd_sc_hd__nor2_1 _4969_ (.A(_1853_),
    .B(_1854_),
    .Y(_1855_));
 sky130_fd_sc_hd__mux2_1 _4970_ (.A0(\z80.tv80s.di_reg[0] ),
    .A1(_1855_),
    .S(_1701_),
    .X(_1856_));
 sky130_fd_sc_hd__a22o_1 _4971_ (.A1(net61),
    .A2(_1852_),
    .B1(_1856_),
    .B2(_1696_),
    .X(_1857_));
 sky130_fd_sc_hd__a211o_1 _4972_ (.A1(\z80.tv80s.i_tv80_core.PC[8] ),
    .A2(_1687_),
    .B1(_1850_),
    .C1(_1857_),
    .X(_1858_));
 sky130_fd_sc_hd__mux2_1 _4973_ (.A0(\z80.tv80s.i_tv80_core.I[0] ),
    .A1(_1858_),
    .S(net99),
    .X(_1859_));
 sky130_fd_sc_hd__a22o_1 _4974_ (.A1(net593),
    .A2(net68),
    .B1(net66),
    .B2(_1859_),
    .X(_1860_));
 sky130_fd_sc_hd__a21bo_1 _4975_ (.A1(net87),
    .A2(_1860_),
    .B1_N(_1848_),
    .X(_1861_));
 sky130_fd_sc_hd__mux2_1 _4976_ (.A0(\z80.tv80s.di_reg[0] ),
    .A1(_1861_),
    .S(net79),
    .X(_1862_));
 sky130_fd_sc_hd__mux2_1 _4977_ (.A0(net581),
    .A1(_1862_),
    .S(net95),
    .X(_1863_));
 sky130_fd_sc_hd__mux2_1 _4978_ (.A0(_1863_),
    .A1(net635),
    .S(net59),
    .X(_0229_));
 sky130_fd_sc_hd__mux4_1 _4979_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][1] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][1] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][1] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][1] ),
    .S0(net138),
    .S1(net167),
    .X(_1864_));
 sky130_fd_sc_hd__mux4_1 _4980_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][1] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][1] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][1] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][1] ),
    .S0(net138),
    .S1(net167),
    .X(_1865_));
 sky130_fd_sc_hd__mux2_2 _4981_ (.A0(_1865_),
    .A1(_1864_),
    .S(net169),
    .X(_1866_));
 sky130_fd_sc_hd__nand2_1 _4982_ (.A(net90),
    .B(_1866_),
    .Y(_1867_));
 sky130_fd_sc_hd__a22o_1 _4983_ (.A1(\z80.tv80s.i_tv80_core.ACC[1] ),
    .A2(_1691_),
    .B1(_1866_),
    .B2(_1690_),
    .X(_1868_));
 sky130_fd_sc_hd__a21o_1 _4984_ (.A1(\z80.tv80s.i_tv80_core.SP[9] ),
    .A2(net62),
    .B1(_1868_),
    .X(_1869_));
 sky130_fd_sc_hd__mux2_1 _4985_ (.A0(\z80.tv80s.i_tv80_core.PC[9] ),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[9] ),
    .S(net140),
    .X(_1870_));
 sky130_fd_sc_hd__mux2_1 _4986_ (.A0(_1866_),
    .A1(_1870_),
    .S(net104),
    .X(_1871_));
 sky130_fd_sc_hd__and2_1 _4987_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[9] ),
    .B(_1853_),
    .X(_1872_));
 sky130_fd_sc_hd__nor2_1 _4988_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[9] ),
    .B(_1853_),
    .Y(_1873_));
 sky130_fd_sc_hd__o21a_1 _4989_ (.A1(_1872_),
    .A2(_1873_),
    .B1(_1701_),
    .X(_1874_));
 sky130_fd_sc_hd__a21oi_1 _4990_ (.A1(_2871_),
    .A2(_1702_),
    .B1(_1874_),
    .Y(_1875_));
 sky130_fd_sc_hd__a22o_1 _4991_ (.A1(net61),
    .A2(_1871_),
    .B1(_1875_),
    .B2(_1696_),
    .X(_1876_));
 sky130_fd_sc_hd__a211o_1 _4992_ (.A1(\z80.tv80s.i_tv80_core.PC[9] ),
    .A2(_1687_),
    .B1(_1869_),
    .C1(_1876_),
    .X(_1877_));
 sky130_fd_sc_hd__mux2_1 _4993_ (.A0(\z80.tv80s.i_tv80_core.I[1] ),
    .A1(_1877_),
    .S(net98),
    .X(_1878_));
 sky130_fd_sc_hd__a22o_1 _4994_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[9] ),
    .A2(net67),
    .B1(net65),
    .B2(_1878_),
    .X(_1879_));
 sky130_fd_sc_hd__a21bo_1 _4995_ (.A1(net87),
    .A2(_1879_),
    .B1_N(_1867_),
    .X(_1880_));
 sky130_fd_sc_hd__mux2_1 _4996_ (.A0(\z80.tv80s.di_reg[1] ),
    .A1(_1880_),
    .S(net79),
    .X(_1881_));
 sky130_fd_sc_hd__mux2_1 _4997_ (.A0(\z80.tv80s.i_tv80_core.I[1] ),
    .A1(_1881_),
    .S(net95),
    .X(_1882_));
 sky130_fd_sc_hd__mux2_1 _4998_ (.A0(_1882_),
    .A1(net556),
    .S(net59),
    .X(_0230_));
 sky130_fd_sc_hd__mux4_1 _4999_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][2] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][2] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][2] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][2] ),
    .S0(net139),
    .S1(net167),
    .X(_1883_));
 sky130_fd_sc_hd__mux4_1 _5000_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][2] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][2] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][2] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][2] ),
    .S0(net139),
    .S1(net168),
    .X(_1884_));
 sky130_fd_sc_hd__mux2_2 _5001_ (.A0(_1884_),
    .A1(_1883_),
    .S(net169),
    .X(_1885_));
 sky130_fd_sc_hd__nand2_1 _5002_ (.A(net90),
    .B(_1885_),
    .Y(_1886_));
 sky130_fd_sc_hd__a22o_1 _5003_ (.A1(\z80.tv80s.i_tv80_core.ACC[2] ),
    .A2(_1691_),
    .B1(_1885_),
    .B2(_1690_),
    .X(_1887_));
 sky130_fd_sc_hd__a21o_1 _5004_ (.A1(\z80.tv80s.i_tv80_core.SP[10] ),
    .A2(net62),
    .B1(_1887_),
    .X(_1888_));
 sky130_fd_sc_hd__mux2_1 _5005_ (.A0(\z80.tv80s.i_tv80_core.PC[10] ),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[10] ),
    .S(net140),
    .X(_1889_));
 sky130_fd_sc_hd__mux2_1 _5006_ (.A0(_1885_),
    .A1(_1889_),
    .S(net104),
    .X(_1890_));
 sky130_fd_sc_hd__xor2_1 _5007_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[10] ),
    .B(_1872_),
    .X(_1891_));
 sky130_fd_sc_hd__mux2_1 _5008_ (.A0(\z80.tv80s.di_reg[2] ),
    .A1(_1891_),
    .S(_1701_),
    .X(_1892_));
 sky130_fd_sc_hd__a22o_1 _5009_ (.A1(net61),
    .A2(_1890_),
    .B1(_1892_),
    .B2(_1696_),
    .X(_1893_));
 sky130_fd_sc_hd__a211o_1 _5010_ (.A1(\z80.tv80s.i_tv80_core.PC[10] ),
    .A2(_1687_),
    .B1(_1888_),
    .C1(_1893_),
    .X(_1894_));
 sky130_fd_sc_hd__mux2_1 _5011_ (.A0(\z80.tv80s.i_tv80_core.I[2] ),
    .A1(_1894_),
    .S(net98),
    .X(_1895_));
 sky130_fd_sc_hd__a22oi_1 _5012_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[10] ),
    .A2(net67),
    .B1(net65),
    .B2(_1895_),
    .Y(_1896_));
 sky130_fd_sc_hd__o21a_1 _5013_ (.A1(net90),
    .A2(_1896_),
    .B1(_1886_),
    .X(_1897_));
 sky130_fd_sc_hd__nand2_1 _5014_ (.A(\z80.tv80s.di_reg[2] ),
    .B(net78),
    .Y(_1898_));
 sky130_fd_sc_hd__o21ai_1 _5015_ (.A1(net78),
    .A2(_1897_),
    .B1(_1898_),
    .Y(_1899_));
 sky130_fd_sc_hd__mux2_1 _5016_ (.A0(\z80.tv80s.i_tv80_core.I[2] ),
    .A1(_1899_),
    .S(net95),
    .X(_1900_));
 sky130_fd_sc_hd__mux2_1 _5017_ (.A0(_1900_),
    .A1(net607),
    .S(net59),
    .X(_0231_));
 sky130_fd_sc_hd__mux4_1 _5018_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][3] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][3] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][3] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][3] ),
    .S0(net138),
    .S1(net167),
    .X(_1901_));
 sky130_fd_sc_hd__mux4_1 _5019_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][3] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][3] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][3] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][3] ),
    .S0(net138),
    .S1(net167),
    .X(_1902_));
 sky130_fd_sc_hd__mux2_4 _5020_ (.A0(_1902_),
    .A1(_1901_),
    .S(net169),
    .X(_1903_));
 sky130_fd_sc_hd__nand2_1 _5021_ (.A(net90),
    .B(_1903_),
    .Y(_1904_));
 sky130_fd_sc_hd__a22o_1 _5022_ (.A1(\z80.tv80s.i_tv80_core.ACC[3] ),
    .A2(_1691_),
    .B1(_1903_),
    .B2(_1690_),
    .X(_1905_));
 sky130_fd_sc_hd__a21o_1 _5023_ (.A1(\z80.tv80s.i_tv80_core.SP[11] ),
    .A2(net62),
    .B1(_1905_),
    .X(_1906_));
 sky130_fd_sc_hd__mux2_1 _5024_ (.A0(\z80.tv80s.i_tv80_core.PC[11] ),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[11] ),
    .S(net140),
    .X(_1907_));
 sky130_fd_sc_hd__mux2_1 _5025_ (.A0(_1903_),
    .A1(_1907_),
    .S(net104),
    .X(_1908_));
 sky130_fd_sc_hd__and3_1 _5026_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[10] ),
    .B(\z80.tv80s.i_tv80_core.TmpAddr[11] ),
    .C(_1872_),
    .X(_1909_));
 sky130_fd_sc_hd__a21oi_1 _5027_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[10] ),
    .A2(_1872_),
    .B1(\z80.tv80s.i_tv80_core.TmpAddr[11] ),
    .Y(_1910_));
 sky130_fd_sc_hd__nor2_1 _5028_ (.A(_1909_),
    .B(_1910_),
    .Y(_1911_));
 sky130_fd_sc_hd__mux2_1 _5029_ (.A0(\z80.tv80s.di_reg[3] ),
    .A1(_1911_),
    .S(_1701_),
    .X(_1912_));
 sky130_fd_sc_hd__a22o_1 _5030_ (.A1(net61),
    .A2(_1908_),
    .B1(_1912_),
    .B2(_1696_),
    .X(_1913_));
 sky130_fd_sc_hd__a211o_1 _5031_ (.A1(\z80.tv80s.i_tv80_core.PC[11] ),
    .A2(_1687_),
    .B1(_1906_),
    .C1(_1913_),
    .X(_1914_));
 sky130_fd_sc_hd__mux2_1 _5032_ (.A0(\z80.tv80s.i_tv80_core.I[3] ),
    .A1(_1914_),
    .S(net98),
    .X(_1915_));
 sky130_fd_sc_hd__a22o_1 _5033_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[11] ),
    .A2(net67),
    .B1(net65),
    .B2(_1915_),
    .X(_1916_));
 sky130_fd_sc_hd__a21bo_1 _5034_ (.A1(net87),
    .A2(_1916_),
    .B1_N(_1904_),
    .X(_1917_));
 sky130_fd_sc_hd__mux2_1 _5035_ (.A0(\z80.tv80s.di_reg[3] ),
    .A1(_1917_),
    .S(net79),
    .X(_1918_));
 sky130_fd_sc_hd__mux2_1 _5036_ (.A0(\z80.tv80s.i_tv80_core.I[3] ),
    .A1(_1918_),
    .S(net93),
    .X(_1919_));
 sky130_fd_sc_hd__mux2_1 _5037_ (.A0(_1919_),
    .A1(net589),
    .S(net59),
    .X(_0232_));
 sky130_fd_sc_hd__mux4_1 _5038_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][4] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][4] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][4] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][4] ),
    .S0(net139),
    .S1(net168),
    .X(_1920_));
 sky130_fd_sc_hd__mux4_1 _5039_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][4] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][4] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][4] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][4] ),
    .S0(net138),
    .S1(net168),
    .X(_1921_));
 sky130_fd_sc_hd__mux2_2 _5040_ (.A0(_1921_),
    .A1(_1920_),
    .S(net169),
    .X(_1922_));
 sky130_fd_sc_hd__nand2_1 _5041_ (.A(net90),
    .B(_1922_),
    .Y(_1923_));
 sky130_fd_sc_hd__a22o_1 _5042_ (.A1(\z80.tv80s.i_tv80_core.ACC[4] ),
    .A2(_1691_),
    .B1(_1922_),
    .B2(_1690_),
    .X(_1924_));
 sky130_fd_sc_hd__a21o_1 _5043_ (.A1(\z80.tv80s.i_tv80_core.SP[12] ),
    .A2(net62),
    .B1(_1924_),
    .X(_1925_));
 sky130_fd_sc_hd__mux2_1 _5044_ (.A0(\z80.tv80s.i_tv80_core.PC[12] ),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[12] ),
    .S(net140),
    .X(_1926_));
 sky130_fd_sc_hd__mux2_1 _5045_ (.A0(_1922_),
    .A1(_1926_),
    .S(net104),
    .X(_1927_));
 sky130_fd_sc_hd__and2_1 _5046_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[12] ),
    .B(_1909_),
    .X(_1928_));
 sky130_fd_sc_hd__nor2_1 _5047_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[12] ),
    .B(_1909_),
    .Y(_1929_));
 sky130_fd_sc_hd__o21ai_1 _5048_ (.A1(_1928_),
    .A2(_1929_),
    .B1(_1701_),
    .Y(_1930_));
 sky130_fd_sc_hd__o21a_1 _5049_ (.A1(\z80.tv80s.di_reg[4] ),
    .A2(_1701_),
    .B1(_1930_),
    .X(_1931_));
 sky130_fd_sc_hd__a22o_1 _5050_ (.A1(net61),
    .A2(_1927_),
    .B1(_1931_),
    .B2(_1696_),
    .X(_1932_));
 sky130_fd_sc_hd__a211o_1 _5051_ (.A1(\z80.tv80s.i_tv80_core.PC[12] ),
    .A2(_1687_),
    .B1(_1925_),
    .C1(_1932_),
    .X(_1933_));
 sky130_fd_sc_hd__mux2_1 _5052_ (.A0(\z80.tv80s.i_tv80_core.I[4] ),
    .A1(_1933_),
    .S(net98),
    .X(_1934_));
 sky130_fd_sc_hd__a22o_1 _5053_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[12] ),
    .A2(net67),
    .B1(net65),
    .B2(_1934_),
    .X(_1935_));
 sky130_fd_sc_hd__a21bo_1 _5054_ (.A1(net87),
    .A2(_1935_),
    .B1_N(_1923_),
    .X(_1936_));
 sky130_fd_sc_hd__mux2_1 _5055_ (.A0(\z80.tv80s.di_reg[4] ),
    .A1(_1936_),
    .S(net79),
    .X(_1937_));
 sky130_fd_sc_hd__mux2_1 _5056_ (.A0(net579),
    .A1(_1937_),
    .S(net93),
    .X(_1938_));
 sky130_fd_sc_hd__mux2_1 _5057_ (.A0(_1938_),
    .A1(net631),
    .S(net59),
    .X(_0233_));
 sky130_fd_sc_hd__mux4_1 _5058_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][5] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][5] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][5] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][5] ),
    .S0(net138),
    .S1(net167),
    .X(_1939_));
 sky130_fd_sc_hd__nand2b_1 _5059_ (.A_N(_1939_),
    .B(net169),
    .Y(_1940_));
 sky130_fd_sc_hd__mux4_2 _5060_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][5] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][5] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][5] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][5] ),
    .S0(net138),
    .S1(net167),
    .X(_1941_));
 sky130_fd_sc_hd__o21ai_4 _5061_ (.A1(net169),
    .A2(_1941_),
    .B1(_1940_),
    .Y(_1942_));
 sky130_fd_sc_hd__inv_2 _5062_ (.A(_1942_),
    .Y(_1943_));
 sky130_fd_sc_hd__nand2_1 _5063_ (.A(net90),
    .B(_1943_),
    .Y(_1944_));
 sky130_fd_sc_hd__nor2_1 _5064_ (.A(_1689_),
    .B(_1942_),
    .Y(_1945_));
 sky130_fd_sc_hd__a221o_1 _5065_ (.A1(\z80.tv80s.i_tv80_core.SP[13] ),
    .A2(net62),
    .B1(_1691_),
    .B2(\z80.tv80s.i_tv80_core.ACC[5] ),
    .C1(_1945_),
    .X(_1946_));
 sky130_fd_sc_hd__mux2_1 _5066_ (.A0(\z80.tv80s.i_tv80_core.PC[13] ),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[13] ),
    .S(net140),
    .X(_1947_));
 sky130_fd_sc_hd__mux2_1 _5067_ (.A0(_1943_),
    .A1(_1947_),
    .S(net104),
    .X(_1948_));
 sky130_fd_sc_hd__xor2_1 _5068_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[13] ),
    .B(_1928_),
    .X(_1949_));
 sky130_fd_sc_hd__mux2_1 _5069_ (.A0(\z80.tv80s.di_reg[5] ),
    .A1(_1949_),
    .S(_1701_),
    .X(_1950_));
 sky130_fd_sc_hd__a22o_1 _5070_ (.A1(net61),
    .A2(_1948_),
    .B1(_1950_),
    .B2(_1696_),
    .X(_1951_));
 sky130_fd_sc_hd__a211o_1 _5071_ (.A1(\z80.tv80s.i_tv80_core.PC[13] ),
    .A2(_1687_),
    .B1(_1946_),
    .C1(_1951_),
    .X(_1952_));
 sky130_fd_sc_hd__mux2_1 _5072_ (.A0(\z80.tv80s.i_tv80_core.I[5] ),
    .A1(_1952_),
    .S(net98),
    .X(_1953_));
 sky130_fd_sc_hd__a22o_1 _5073_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[13] ),
    .A2(net67),
    .B1(net65),
    .B2(_1953_),
    .X(_1954_));
 sky130_fd_sc_hd__a21bo_1 _5074_ (.A1(net87),
    .A2(_1954_),
    .B1_N(_1944_),
    .X(_1955_));
 sky130_fd_sc_hd__mux2_1 _5075_ (.A0(\z80.tv80s.di_reg[5] ),
    .A1(_1955_),
    .S(net79),
    .X(_1956_));
 sky130_fd_sc_hd__mux2_1 _5076_ (.A0(\z80.tv80s.i_tv80_core.I[5] ),
    .A1(_1956_),
    .S(net93),
    .X(_1957_));
 sky130_fd_sc_hd__mux2_1 _5077_ (.A0(_1957_),
    .A1(net647),
    .S(net59),
    .X(_0234_));
 sky130_fd_sc_hd__mux4_1 _5078_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][6] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][6] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][6] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][6] ),
    .S0(net139),
    .S1(net168),
    .X(_1958_));
 sky130_fd_sc_hd__mux4_1 _5079_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][6] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][6] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][6] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][6] ),
    .S0(net138),
    .S1(net167),
    .X(_1959_));
 sky130_fd_sc_hd__mux2_2 _5080_ (.A0(_1959_),
    .A1(_1958_),
    .S(net169),
    .X(_1960_));
 sky130_fd_sc_hd__nand2_1 _5081_ (.A(net90),
    .B(_1960_),
    .Y(_1961_));
 sky130_fd_sc_hd__a22o_1 _5082_ (.A1(\z80.tv80s.i_tv80_core.ACC[6] ),
    .A2(_1691_),
    .B1(_1960_),
    .B2(_1690_),
    .X(_1962_));
 sky130_fd_sc_hd__a21o_1 _5083_ (.A1(\z80.tv80s.i_tv80_core.SP[14] ),
    .A2(net62),
    .B1(_1962_),
    .X(_1963_));
 sky130_fd_sc_hd__mux2_1 _5084_ (.A0(\z80.tv80s.i_tv80_core.PC[14] ),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[14] ),
    .S(net140),
    .X(_1964_));
 sky130_fd_sc_hd__mux2_1 _5085_ (.A0(_1960_),
    .A1(_1964_),
    .S(net104),
    .X(_1965_));
 sky130_fd_sc_hd__and3_1 _5086_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[13] ),
    .B(\z80.tv80s.i_tv80_core.TmpAddr[14] ),
    .C(_1928_),
    .X(_1966_));
 sky130_fd_sc_hd__a21oi_1 _5087_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[13] ),
    .A2(_1928_),
    .B1(\z80.tv80s.i_tv80_core.TmpAddr[14] ),
    .Y(_1967_));
 sky130_fd_sc_hd__o21a_1 _5088_ (.A1(_1966_),
    .A2(_1967_),
    .B1(_1701_),
    .X(_1968_));
 sky130_fd_sc_hd__o21ba_1 _5089_ (.A1(\z80.tv80s.di_reg[6] ),
    .A2(_1701_),
    .B1_N(_1968_),
    .X(_1969_));
 sky130_fd_sc_hd__a22o_1 _5090_ (.A1(net61),
    .A2(_1965_),
    .B1(_1969_),
    .B2(_1696_),
    .X(_1970_));
 sky130_fd_sc_hd__a211o_1 _5091_ (.A1(\z80.tv80s.i_tv80_core.PC[14] ),
    .A2(_1687_),
    .B1(_1963_),
    .C1(_1970_),
    .X(_1971_));
 sky130_fd_sc_hd__mux2_1 _5092_ (.A0(\z80.tv80s.i_tv80_core.I[6] ),
    .A1(_1971_),
    .S(net98),
    .X(_1972_));
 sky130_fd_sc_hd__a22oi_1 _5093_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[14] ),
    .A2(net67),
    .B1(net65),
    .B2(_1972_),
    .Y(_1973_));
 sky130_fd_sc_hd__o21a_1 _5094_ (.A1(net90),
    .A2(_1973_),
    .B1(_1961_),
    .X(_1974_));
 sky130_fd_sc_hd__nand2_1 _5095_ (.A(\z80.tv80s.di_reg[6] ),
    .B(net78),
    .Y(_1975_));
 sky130_fd_sc_hd__o21ai_1 _5096_ (.A1(net78),
    .A2(_1974_),
    .B1(_1975_),
    .Y(_1976_));
 sky130_fd_sc_hd__mux2_1 _5097_ (.A0(\z80.tv80s.i_tv80_core.I[6] ),
    .A1(_1976_),
    .S(net93),
    .X(_1977_));
 sky130_fd_sc_hd__mux2_1 _5098_ (.A0(_1977_),
    .A1(net724),
    .S(net59),
    .X(_0235_));
 sky130_fd_sc_hd__mux4_1 _5099_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][7] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][7] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][7] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][7] ),
    .S0(net138),
    .S1(net167),
    .X(_1978_));
 sky130_fd_sc_hd__mux4_1 _5100_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][7] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][7] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][7] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][7] ),
    .S0(net138),
    .S1(net167),
    .X(_1979_));
 sky130_fd_sc_hd__mux2_2 _5101_ (.A0(_1979_),
    .A1(_1978_),
    .S(net169),
    .X(_1980_));
 sky130_fd_sc_hd__nand2_1 _5102_ (.A(net90),
    .B(_1980_),
    .Y(_1981_));
 sky130_fd_sc_hd__a22o_1 _5103_ (.A1(\z80.tv80s.i_tv80_core.ACC[7] ),
    .A2(_1691_),
    .B1(_1980_),
    .B2(_1690_),
    .X(_1982_));
 sky130_fd_sc_hd__a21o_1 _5104_ (.A1(\z80.tv80s.i_tv80_core.SP[15] ),
    .A2(net62),
    .B1(_1982_),
    .X(_1983_));
 sky130_fd_sc_hd__mux2_1 _5105_ (.A0(\z80.tv80s.i_tv80_core.PC[15] ),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[15] ),
    .S(net140),
    .X(_1984_));
 sky130_fd_sc_hd__mux2_1 _5106_ (.A0(_1980_),
    .A1(_1984_),
    .S(net104),
    .X(_1985_));
 sky130_fd_sc_hd__xor2_1 _5107_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[15] ),
    .B(_1966_),
    .X(_1986_));
 sky130_fd_sc_hd__mux2_1 _5108_ (.A0(\z80.tv80s.di_reg[7] ),
    .A1(_1986_),
    .S(_1701_),
    .X(_1987_));
 sky130_fd_sc_hd__a22o_1 _5109_ (.A1(net61),
    .A2(_1985_),
    .B1(_1987_),
    .B2(_1696_),
    .X(_1988_));
 sky130_fd_sc_hd__a211o_1 _5110_ (.A1(\z80.tv80s.i_tv80_core.PC[15] ),
    .A2(_1687_),
    .B1(_1983_),
    .C1(_1988_),
    .X(_1989_));
 sky130_fd_sc_hd__mux2_1 _5111_ (.A0(\z80.tv80s.i_tv80_core.I[7] ),
    .A1(_1989_),
    .S(net98),
    .X(_1990_));
 sky130_fd_sc_hd__a22o_1 _5112_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[15] ),
    .A2(net67),
    .B1(net65),
    .B2(_1990_),
    .X(_1991_));
 sky130_fd_sc_hd__a21bo_1 _5113_ (.A1(net87),
    .A2(_1991_),
    .B1_N(_1981_),
    .X(_1992_));
 sky130_fd_sc_hd__mux2_1 _5114_ (.A0(\z80.tv80s.di_reg[7] ),
    .A1(_1992_),
    .S(net79),
    .X(_1993_));
 sky130_fd_sc_hd__mux2_1 _5115_ (.A0(\z80.tv80s.i_tv80_core.I[7] ),
    .A1(_1993_),
    .S(net93),
    .X(_1994_));
 sky130_fd_sc_hd__mux2_1 _5116_ (.A0(_1994_),
    .A1(net629),
    .S(_1666_),
    .X(_0236_));
 sky130_fd_sc_hd__or3b_1 _5117_ (.A(_2873_),
    .B(_2875_),
    .C_N(_0781_),
    .X(_1995_));
 sky130_fd_sc_hd__or4b_4 _5118_ (.A(net501),
    .B(_2874_),
    .C(_1995_),
    .D_N(net508),
    .X(_1996_));
 sky130_fd_sc_hd__nor2_1 _5119_ (.A(_0856_),
    .B(_1996_),
    .Y(_1997_));
 sky130_fd_sc_hd__a21oi_4 _5120_ (.A1(net837),
    .A2(_0713_),
    .B1(_0851_),
    .Y(_1998_));
 sky130_fd_sc_hd__a21o_2 _5121_ (.A1(\z80.tv80s.i_tv80_core.Save_ALU_r ),
    .A2(_0713_),
    .B1(_0851_),
    .X(_1999_));
 sky130_fd_sc_hd__or2_1 _5122_ (.A(net60),
    .B(net92),
    .X(_2000_));
 sky130_fd_sc_hd__inv_2 _5123_ (.A(_2000_),
    .Y(_2001_));
 sky130_fd_sc_hd__or3_4 _5124_ (.A(_2846_),
    .B(net118),
    .C(_2930_),
    .X(_2002_));
 sky130_fd_sc_hd__inv_2 _5125_ (.A(_2002_),
    .Y(_2003_));
 sky130_fd_sc_hd__a21oi_1 _5126_ (.A1(net154),
    .A2(\z80.tv80s.i_tv80_core.F[0] ),
    .B1(_2002_),
    .Y(_2004_));
 sky130_fd_sc_hd__a211o_1 _5127_ (.A1(\z80.tv80s.i_tv80_core.F[0] ),
    .A2(_2002_),
    .B1(_2004_),
    .C1(_2000_),
    .X(_2005_));
 sky130_fd_sc_hd__o21ai_1 _5128_ (.A1(net734),
    .A2(_1498_),
    .B1(_2005_),
    .Y(_2006_));
 sky130_fd_sc_hd__nor2_1 _5129_ (.A(net60),
    .B(net102),
    .Y(_2007_));
 sky130_fd_sc_hd__or2_2 _5130_ (.A(net60),
    .B(net102),
    .X(_2008_));
 sky130_fd_sc_hd__nor2_1 _5131_ (.A(_1502_),
    .B(_2007_),
    .Y(_2009_));
 sky130_fd_sc_hd__or2_1 _5132_ (.A(_1502_),
    .B(_2007_),
    .X(_2010_));
 sky130_fd_sc_hd__a2bb2o_1 _5133_ (.A1_N(\z80.tv80s.i_tv80_core.F[0] ),
    .A2_N(_2010_),
    .B1(_2006_),
    .B2(net94),
    .X(_2011_));
 sky130_fd_sc_hd__o21ai_1 _5134_ (.A1(net526),
    .A2(_1998_),
    .B1(_2011_),
    .Y(_2012_));
 sky130_fd_sc_hd__a21bo_1 _5135_ (.A1(net162),
    .A2(_1260_),
    .B1_N(_1264_),
    .X(_2013_));
 sky130_fd_sc_hd__nor2_1 _5136_ (.A(net111),
    .B(_0815_),
    .Y(_2014_));
 sky130_fd_sc_hd__nor2_1 _5137_ (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[2] ),
    .B(\z80.tv80s.i_tv80_core.ALU_Op_r[1] ),
    .Y(_2015_));
 sky130_fd_sc_hd__mux2_1 _5138_ (.A0(_2014_),
    .A1(_2015_),
    .S(_2013_),
    .X(_2016_));
 sky130_fd_sc_hd__o211a_1 _5139_ (.A1(\z80.tv80s.i_tv80_core.ALU_Op_r[0] ),
    .A2(net143),
    .B1(\z80.tv80s.i_tv80_core.F[0] ),
    .C1(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ),
    .X(_2017_));
 sky130_fd_sc_hd__a21o_1 _5140_ (.A1(net120),
    .A2(net162),
    .B1(_1285_),
    .X(_2018_));
 sky130_fd_sc_hd__a2111o_1 _5141_ (.A1(_0839_),
    .A2(_2018_),
    .B1(_1998_),
    .C1(net526),
    .D1(_2017_),
    .X(_2019_));
 sky130_fd_sc_hd__a221o_1 _5142_ (.A1(_0848_),
    .A2(_1174_),
    .B1(_2016_),
    .B2(_2862_),
    .C1(_2019_),
    .X(_2020_));
 sky130_fd_sc_hd__a31o_1 _5143_ (.A1(_1996_),
    .A2(_2012_),
    .A3(_2020_),
    .B1(_1997_),
    .X(_2021_));
 sky130_fd_sc_hd__mux2_1 _5144_ (.A0(net863),
    .A1(_2021_),
    .S(net115),
    .X(_0237_));
 sky130_fd_sc_hd__or4_4 _5145_ (.A(_2848_),
    .B(net105),
    .C(net60),
    .D(_1327_),
    .X(_2022_));
 sky130_fd_sc_hd__or4_4 _5146_ (.A(_2855_),
    .B(_3049_),
    .C(net105),
    .D(_0653_),
    .X(_2023_));
 sky130_fd_sc_hd__and3_1 _5147_ (.A(_1996_),
    .B(_2022_),
    .C(_2023_),
    .X(_2024_));
 sky130_fd_sc_hd__o221a_1 _5148_ (.A1(_2862_),
    .A2(\z80.tv80s.i_tv80_core.F[1] ),
    .B1(_0848_),
    .B2(_2014_),
    .C1(_1999_),
    .X(_2025_));
 sky130_fd_sc_hd__o21a_1 _5149_ (.A1(\z80.tv80s.i_tv80_core.F[1] ),
    .A2(_1618_),
    .B1(_2002_),
    .X(_2026_));
 sky130_fd_sc_hd__o22a_1 _5150_ (.A1(\z80.tv80s.i_tv80_core.Fp[1] ),
    .A2(_1498_),
    .B1(_2000_),
    .B2(_2026_),
    .X(_2027_));
 sky130_fd_sc_hd__nor2_1 _5151_ (.A(_1626_),
    .B(_1999_),
    .Y(_2028_));
 sky130_fd_sc_hd__o22a_1 _5152_ (.A1(\z80.tv80s.i_tv80_core.F[1] ),
    .A2(_2010_),
    .B1(_2027_),
    .B2(net102),
    .X(_2029_));
 sky130_fd_sc_hd__a21o_1 _5153_ (.A1(_2028_),
    .A2(_2029_),
    .B1(_2025_),
    .X(_2030_));
 sky130_fd_sc_hd__a2bb2o_1 _5154_ (.A1_N(_1014_),
    .A2_N(_1996_),
    .B1(_2024_),
    .B2(_2030_),
    .X(_2031_));
 sky130_fd_sc_hd__mux2_1 _5155_ (.A0(net865),
    .A1(_2031_),
    .S(net115),
    .X(_0238_));
 sky130_fd_sc_hd__mux2_1 _5156_ (.A0(\z80.tv80s.i_tv80_core.F[2] ),
    .A1(\z80.tv80s.i_tv80_core.Fp[2] ),
    .S(_1502_),
    .X(_2032_));
 sky130_fd_sc_hd__mux2_1 _5157_ (.A0(_2032_),
    .A1(\z80.tv80s.i_tv80_core.IntE_FF2 ),
    .S(_1626_),
    .X(_2033_));
 sky130_fd_sc_hd__or3b_1 _5158_ (.A(net162),
    .B(_1262_),
    .C_N(_1260_),
    .X(_2034_));
 sky130_fd_sc_hd__o21ai_1 _5159_ (.A1(_1260_),
    .A2(_1264_),
    .B1(_2034_),
    .Y(_2035_));
 sky130_fd_sc_hd__xor2_1 _5160_ (.A(_1228_),
    .B(_1270_),
    .X(_2036_));
 sky130_fd_sc_hd__xnor2_1 _5161_ (.A(_1141_),
    .B(_1169_),
    .Y(_2037_));
 sky130_fd_sc_hd__xor2_1 _5162_ (.A(_0831_),
    .B(_0998_),
    .X(_2038_));
 sky130_fd_sc_hd__xnor2_1 _5163_ (.A(_1051_),
    .B(_1083_),
    .Y(_2039_));
 sky130_fd_sc_hd__xnor2_1 _5164_ (.A(_2038_),
    .B(_2039_),
    .Y(_2040_));
 sky130_fd_sc_hd__xnor2_1 _5165_ (.A(_2037_),
    .B(_2040_),
    .Y(_2041_));
 sky130_fd_sc_hd__nor2_1 _5166_ (.A(_2036_),
    .B(_2041_),
    .Y(_2042_));
 sky130_fd_sc_hd__a21o_1 _5167_ (.A1(_2036_),
    .A2(_2041_),
    .B1(_0827_),
    .X(_2043_));
 sky130_fd_sc_hd__o22a_1 _5168_ (.A1(_0826_),
    .A2(_2035_),
    .B1(_2042_),
    .B2(_2043_),
    .X(_2044_));
 sky130_fd_sc_hd__mux2_1 _5169_ (.A0(\z80.tv80s.i_tv80_core.F[2] ),
    .A1(_2044_),
    .S(_2870_),
    .X(_2045_));
 sky130_fd_sc_hd__xor2_1 _5170_ (.A(\z80.tv80s.i_tv80_core.BusA[0] ),
    .B(_1010_),
    .X(_2046_));
 sky130_fd_sc_hd__xor2_1 _5171_ (.A(_1236_),
    .B(_1282_),
    .X(_2047_));
 sky130_fd_sc_hd__xnor2_1 _5172_ (.A(_2046_),
    .B(_2047_),
    .Y(_2048_));
 sky130_fd_sc_hd__nand2_1 _5173_ (.A(_1127_),
    .B(_1182_),
    .Y(_2049_));
 sky130_fd_sc_hd__xnor2_1 _5174_ (.A(_1127_),
    .B(_1181_),
    .Y(_2050_));
 sky130_fd_sc_hd__xnor2_1 _5175_ (.A(_1055_),
    .B(_1089_),
    .Y(_2051_));
 sky130_fd_sc_hd__xnor2_1 _5176_ (.A(_2050_),
    .B(_2051_),
    .Y(_2052_));
 sky130_fd_sc_hd__xnor2_1 _5177_ (.A(_2048_),
    .B(_2052_),
    .Y(_2053_));
 sky130_fd_sc_hd__nand2_1 _5178_ (.A(\z80.tv80s.i_tv80_core.F[1] ),
    .B(_1279_),
    .Y(_2054_));
 sky130_fd_sc_hd__o211a_1 _5179_ (.A1(\z80.tv80s.i_tv80_core.F[1] ),
    .A2(_1172_),
    .B1(_1174_),
    .C1(_2054_),
    .X(_2055_));
 sky130_fd_sc_hd__xnor2_1 _5180_ (.A(_2053_),
    .B(_2055_),
    .Y(_2056_));
 sky130_fd_sc_hd__xor2_1 _5181_ (.A(_1238_),
    .B(_1287_),
    .X(_2057_));
 sky130_fd_sc_hd__xnor2_1 _5182_ (.A(_0842_),
    .B(_1000_),
    .Y(_2058_));
 sky130_fd_sc_hd__xor2_1 _5183_ (.A(_1057_),
    .B(_1091_),
    .X(_2059_));
 sky130_fd_sc_hd__xor2_1 _5184_ (.A(_1129_),
    .B(_1184_),
    .X(_2060_));
 sky130_fd_sc_hd__xnor2_1 _5185_ (.A(_2059_),
    .B(_2060_),
    .Y(_2061_));
 sky130_fd_sc_hd__xnor2_1 _5186_ (.A(_2058_),
    .B(_2061_),
    .Y(_2062_));
 sky130_fd_sc_hd__nor2_1 _5187_ (.A(_2057_),
    .B(_2062_),
    .Y(_2063_));
 sky130_fd_sc_hd__a21o_1 _5188_ (.A1(_2057_),
    .A2(_2062_),
    .B1(net166),
    .X(_2064_));
 sky130_fd_sc_hd__o22a_1 _5189_ (.A1(net119),
    .A2(\z80.tv80s.i_tv80_core.F[2] ),
    .B1(_2063_),
    .B2(_2064_),
    .X(_2065_));
 sky130_fd_sc_hd__xor2_1 _5190_ (.A(_1056_),
    .B(_1090_),
    .X(_2066_));
 sky130_fd_sc_hd__xor2_1 _5191_ (.A(_0846_),
    .B(_0999_),
    .X(_2067_));
 sky130_fd_sc_hd__xnor2_1 _5192_ (.A(_2066_),
    .B(_2067_),
    .Y(_2068_));
 sky130_fd_sc_hd__xor2_1 _5193_ (.A(\z80.tv80s.i_tv80_core.BusA[4] ),
    .B(\z80.tv80s.i_tv80_core.BusA[5] ),
    .X(_2069_));
 sky130_fd_sc_hd__xnor2_1 _5194_ (.A(_1272_),
    .B(_2069_),
    .Y(_2070_));
 sky130_fd_sc_hd__xnor2_1 _5195_ (.A(_2068_),
    .B(_2070_),
    .Y(_2071_));
 sky130_fd_sc_hd__a22o_1 _5196_ (.A1(\z80.tv80s.i_tv80_core.BusB[1] ),
    .A2(_1001_),
    .B1(_1059_),
    .B2(\z80.tv80s.i_tv80_core.BusB[2] ),
    .X(_2072_));
 sky130_fd_sc_hd__a22o_1 _5197_ (.A1(\z80.tv80s.i_tv80_core.BusB[5] ),
    .A2(_0470_),
    .B1(_0835_),
    .B2(\z80.tv80s.i_tv80_core.BusB[0] ),
    .X(_2073_));
 sky130_fd_sc_hd__a22o_1 _5198_ (.A1(\z80.tv80s.i_tv80_core.BusB[6] ),
    .A2(_0405_),
    .B1(_0468_),
    .B2(\z80.tv80s.i_tv80_core.BusB[3] ),
    .X(_2074_));
 sky130_fd_sc_hd__or4b_1 _5199_ (.A(_1290_),
    .B(_2073_),
    .C(_2074_),
    .D_N(_0851_),
    .X(_2075_));
 sky130_fd_sc_hd__a211o_1 _5200_ (.A1(\z80.tv80s.i_tv80_core.BusB[4] ),
    .A2(_0471_),
    .B1(_2072_),
    .C1(_2075_),
    .X(_2076_));
 sky130_fd_sc_hd__and2_2 _5201_ (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ),
    .B(_2014_),
    .X(_2077_));
 sky130_fd_sc_hd__inv_2 _5202_ (.A(_2077_),
    .Y(_2078_));
 sky130_fd_sc_hd__a22o_1 _5203_ (.A1(_0839_),
    .A2(_2065_),
    .B1(_2071_),
    .B2(_0844_),
    .X(_2079_));
 sky130_fd_sc_hd__a221o_1 _5204_ (.A1(_0848_),
    .A2(_2056_),
    .B1(_2077_),
    .B2(\z80.tv80s.i_tv80_core.F[2] ),
    .C1(_1998_),
    .X(_2080_));
 sky130_fd_sc_hd__a21o_1 _5205_ (.A1(_2862_),
    .A2(_2045_),
    .B1(_2080_),
    .X(_2081_));
 sky130_fd_sc_hd__or3b_1 _5206_ (.A(_2079_),
    .B(_2081_),
    .C_N(_2076_),
    .X(_2082_));
 sky130_fd_sc_hd__or2_1 _5207_ (.A(\z80.tv80s.di_reg[5] ),
    .B(\z80.tv80s.di_reg[4] ),
    .X(_2083_));
 sky130_fd_sc_hd__nand2_1 _5208_ (.A(\z80.tv80s.di_reg[5] ),
    .B(\z80.tv80s.di_reg[4] ),
    .Y(_2084_));
 sky130_fd_sc_hd__nand2_1 _5209_ (.A(_2083_),
    .B(_2084_),
    .Y(_2085_));
 sky130_fd_sc_hd__xor2_1 _5210_ (.A(\z80.tv80s.di_reg[1] ),
    .B(\z80.tv80s.di_reg[0] ),
    .X(_2086_));
 sky130_fd_sc_hd__xor2_1 _5211_ (.A(\z80.tv80s.di_reg[7] ),
    .B(\z80.tv80s.di_reg[6] ),
    .X(_2087_));
 sky130_fd_sc_hd__xor2_1 _5212_ (.A(\z80.tv80s.di_reg[3] ),
    .B(\z80.tv80s.di_reg[2] ),
    .X(_2088_));
 sky130_fd_sc_hd__xnor2_1 _5213_ (.A(_2087_),
    .B(_2088_),
    .Y(_2089_));
 sky130_fd_sc_hd__xnor2_1 _5214_ (.A(_2086_),
    .B(_2089_),
    .Y(_2090_));
 sky130_fd_sc_hd__xnor2_1 _5215_ (.A(_2085_),
    .B(_2090_),
    .Y(_2091_));
 sky130_fd_sc_hd__o21a_1 _5216_ (.A1(_1999_),
    .A2(_2033_),
    .B1(_2022_),
    .X(_2092_));
 sky130_fd_sc_hd__a2bb2o_1 _5217_ (.A1_N(_2022_),
    .A2_N(_2091_),
    .B1(_2092_),
    .B2(_2082_),
    .X(_2093_));
 sky130_fd_sc_hd__mux2_1 _5218_ (.A0(net429),
    .A1(_2093_),
    .S(_0672_),
    .X(_2094_));
 sky130_fd_sc_hd__mux2_1 _5219_ (.A0(_1067_),
    .A1(_2094_),
    .S(_1996_),
    .X(_2095_));
 sky130_fd_sc_hd__mux2_1 _5220_ (.A0(net856),
    .A1(_2095_),
    .S(net116),
    .X(_0239_));
 sky130_fd_sc_hd__and2b_1 _5221_ (.A_N(_2023_),
    .B(_1097_),
    .X(_2096_));
 sky130_fd_sc_hd__mux2_1 _5222_ (.A0(\z80.tv80s.i_tv80_core.F[3] ),
    .A1(_2878_),
    .S(_1618_),
    .X(_2097_));
 sky130_fd_sc_hd__mux2_1 _5223_ (.A0(\z80.tv80s.i_tv80_core.ACC[3] ),
    .A1(_2097_),
    .S(_2002_),
    .X(_2098_));
 sky130_fd_sc_hd__a22o_1 _5224_ (.A1(\z80.tv80s.i_tv80_core.Fp[3] ),
    .A2(net91),
    .B1(_2001_),
    .B2(_2098_),
    .X(_2099_));
 sky130_fd_sc_hd__a221o_1 _5225_ (.A1(\z80.tv80s.i_tv80_core.F[3] ),
    .A2(_2009_),
    .B1(_2099_),
    .B2(net95),
    .C1(_1999_),
    .X(_2100_));
 sky130_fd_sc_hd__mux2_1 _5226_ (.A0(\z80.tv80s.i_tv80_core.BusB[3] ),
    .A1(_1083_),
    .S(_0778_),
    .X(_2101_));
 sky130_fd_sc_hd__a31o_1 _5227_ (.A1(\z80.tv80s.i_tv80_core.BusB[3] ),
    .A2(net97),
    .A3(_0851_),
    .B1(_1092_),
    .X(_2102_));
 sky130_fd_sc_hd__a211o_1 _5228_ (.A1(\z80.tv80s.i_tv80_core.F[3] ),
    .A2(_2077_),
    .B1(_2102_),
    .C1(_1998_),
    .X(_2103_));
 sky130_fd_sc_hd__a211o_1 _5229_ (.A1(_2862_),
    .A2(_2101_),
    .B1(_2103_),
    .C1(_1095_),
    .X(_2104_));
 sky130_fd_sc_hd__a31o_1 _5230_ (.A1(_2023_),
    .A2(_2100_),
    .A3(_2104_),
    .B1(_2096_),
    .X(_2105_));
 sky130_fd_sc_hd__mux2_1 _5231_ (.A0(_1101_),
    .A1(_2105_),
    .S(_1996_),
    .X(_2106_));
 sky130_fd_sc_hd__mux2_1 _5232_ (.A0(net823),
    .A1(_2106_),
    .S(net115),
    .X(_0240_));
 sky130_fd_sc_hd__and2b_1 _5233_ (.A_N(_1136_),
    .B(_2014_),
    .X(_2107_));
 sky130_fd_sc_hd__a221o_1 _5234_ (.A1(\z80.tv80s.i_tv80_core.ALU_Op_r[2] ),
    .A2(_0821_),
    .B1(_1136_),
    .B2(_2015_),
    .C1(_2107_),
    .X(_2108_));
 sky130_fd_sc_hd__a2bb2o_1 _5235_ (.A1_N(_0849_),
    .A2_N(_1126_),
    .B1(_2108_),
    .B2(_2862_),
    .X(_2109_));
 sky130_fd_sc_hd__a211o_1 _5236_ (.A1(\z80.tv80s.i_tv80_core.F[4] ),
    .A2(_2077_),
    .B1(_2109_),
    .C1(_0851_),
    .X(_2110_));
 sky130_fd_sc_hd__a311o_1 _5237_ (.A1(net154),
    .A2(_2003_),
    .A3(_2007_),
    .B1(\z80.tv80s.i_tv80_core.F[4] ),
    .C1(_1621_),
    .X(_2111_));
 sky130_fd_sc_hd__o2bb2a_1 _5238_ (.A1_N(_2001_),
    .A2_N(_2004_),
    .B1(\z80.tv80s.i_tv80_core.Fp[4] ),
    .B2(_1498_),
    .X(_2112_));
 sky130_fd_sc_hd__or2_1 _5239_ (.A(net102),
    .B(_2112_),
    .X(_2113_));
 sky130_fd_sc_hd__a32o_1 _5240_ (.A1(_2028_),
    .A2(_2111_),
    .A3(_2113_),
    .B1(_2110_),
    .B2(_1999_),
    .X(_2114_));
 sky130_fd_sc_hd__a2bb2o_1 _5241_ (.A1_N(_1150_),
    .A2_N(_1996_),
    .B1(_2024_),
    .B2(_2114_),
    .X(_2115_));
 sky130_fd_sc_hd__mux2_1 _5242_ (.A0(net830),
    .A1(_2115_),
    .S(net116),
    .X(_0241_));
 sky130_fd_sc_hd__mux2_1 _5243_ (.A0(\z80.tv80s.i_tv80_core.F[5] ),
    .A1(_2879_),
    .S(_1618_),
    .X(_2116_));
 sky130_fd_sc_hd__mux2_1 _5244_ (.A0(\z80.tv80s.i_tv80_core.ACC[5] ),
    .A1(_2116_),
    .S(_2002_),
    .X(_2117_));
 sky130_fd_sc_hd__a22o_1 _5245_ (.A1(\z80.tv80s.i_tv80_core.Fp[5] ),
    .A2(net92),
    .B1(_2001_),
    .B2(_2117_),
    .X(_2118_));
 sky130_fd_sc_hd__a221o_1 _5246_ (.A1(\z80.tv80s.i_tv80_core.F[5] ),
    .A2(_2009_),
    .B1(_2118_),
    .B2(net94),
    .C1(_1999_),
    .X(_2119_));
 sky130_fd_sc_hd__mux2_1 _5247_ (.A0(\z80.tv80s.i_tv80_core.BusB[5] ),
    .A1(_1169_),
    .S(_0778_),
    .X(_2120_));
 sky130_fd_sc_hd__a311o_1 _5248_ (.A1(\z80.tv80s.i_tv80_core.BusB[5] ),
    .A2(net97),
    .A3(_0851_),
    .B1(_1183_),
    .C1(_1185_),
    .X(_2121_));
 sky130_fd_sc_hd__a221o_1 _5249_ (.A1(\z80.tv80s.i_tv80_core.F[5] ),
    .A2(_2077_),
    .B1(_2120_),
    .B2(_2862_),
    .C1(_2121_),
    .X(_2122_));
 sky130_fd_sc_hd__o21a_1 _5250_ (.A1(_1998_),
    .A2(_2122_),
    .B1(_2023_),
    .X(_2123_));
 sky130_fd_sc_hd__o2bb2a_1 _5251_ (.A1_N(_2123_),
    .A2_N(_2119_),
    .B1(_2023_),
    .B2(_1012_),
    .X(_2124_));
 sky130_fd_sc_hd__mux2_1 _5252_ (.A0(_1191_),
    .A1(_2124_),
    .S(_1996_),
    .X(_2125_));
 sky130_fd_sc_hd__inv_2 _5253_ (.A(_2125_),
    .Y(_2126_));
 sky130_fd_sc_hd__mux2_1 _5254_ (.A0(net818),
    .A1(_2126_),
    .S(net116),
    .X(_0242_));
 sky130_fd_sc_hd__a211o_1 _5255_ (.A1(_2852_),
    .A2(\z80.tv80s.i_tv80_core.Z16_r ),
    .B1(_0831_),
    .C1(_0998_),
    .X(_2127_));
 sky130_fd_sc_hd__or3b_1 _5256_ (.A(_2127_),
    .B(_1083_),
    .C_N(_1051_),
    .X(_2128_));
 sky130_fd_sc_hd__or3_1 _5257_ (.A(_1142_),
    .B(_1169_),
    .C(_2128_),
    .X(_2129_));
 sky130_fd_sc_hd__o31a_1 _5258_ (.A1(_1228_),
    .A2(_1270_),
    .A3(_2129_),
    .B1(_2870_),
    .X(_2130_));
 sky130_fd_sc_hd__a211o_1 _5259_ (.A1(_2852_),
    .A2(\z80.tv80s.i_tv80_core.Arith16_r ),
    .B1(_2130_),
    .C1(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ),
    .X(_2131_));
 sky130_fd_sc_hd__or3b_1 _5260_ (.A(_0849_),
    .B(_1055_),
    .C_N(_1089_),
    .X(_2132_));
 sky130_fd_sc_hd__or4b_1 _5261_ (.A(\z80.tv80s.i_tv80_core.BusA[0] ),
    .B(_2049_),
    .C(_2132_),
    .D_N(_1010_),
    .X(_2133_));
 sky130_fd_sc_hd__or4_1 _5262_ (.A(_1057_),
    .B(_1091_),
    .C(_1129_),
    .D(_1184_),
    .X(_2134_));
 sky130_fd_sc_hd__or3_1 _5263_ (.A(_1238_),
    .B(_1287_),
    .C(_2134_),
    .X(_2135_));
 sky130_fd_sc_hd__or3_1 _5264_ (.A(_0843_),
    .B(_1000_),
    .C(_2135_),
    .X(_2136_));
 sky130_fd_sc_hd__o21ai_1 _5265_ (.A1(net118),
    .A2(\z80.tv80s.i_tv80_core.F[6] ),
    .B1(_0839_),
    .Y(_2137_));
 sky130_fd_sc_hd__a21o_1 _5266_ (.A1(net118),
    .A2(_2136_),
    .B1(_2137_),
    .X(_2138_));
 sky130_fd_sc_hd__or4_1 _5267_ (.A(_0846_),
    .B(_0999_),
    .C(_1056_),
    .D(_1090_),
    .X(_2139_));
 sky130_fd_sc_hd__or4_1 _5268_ (.A(net162),
    .B(\z80.tv80s.i_tv80_core.BusA[4] ),
    .C(\z80.tv80s.i_tv80_core.BusA[5] ),
    .D(\z80.tv80s.i_tv80_core.BusA[6] ),
    .X(_2140_));
 sky130_fd_sc_hd__o311a_1 _5269_ (.A1(_0845_),
    .A2(_2139_),
    .A3(_2140_),
    .B1(_2076_),
    .C1(_2078_),
    .X(_2141_));
 sky130_fd_sc_hd__o31a_1 _5270_ (.A1(_1236_),
    .A2(_1282_),
    .A3(_2133_),
    .B1(_2141_),
    .X(_2142_));
 sky130_fd_sc_hd__a32o_1 _5271_ (.A1(_2131_),
    .A2(_2138_),
    .A3(_2142_),
    .B1(_2077_),
    .B2(_2852_),
    .X(_2143_));
 sky130_fd_sc_hd__o31a_1 _5272_ (.A1(\z80.tv80s.i_tv80_core.Fp[6] ),
    .A2(net102),
    .A3(_1498_),
    .B1(_1625_),
    .X(_2144_));
 sky130_fd_sc_hd__o21ai_1 _5273_ (.A1(\z80.tv80s.i_tv80_core.F[6] ),
    .A2(_1502_),
    .B1(_2144_),
    .Y(_2145_));
 sky130_fd_sc_hd__or4_1 _5274_ (.A(\z80.tv80s.i_tv80_core.I[1] ),
    .B(\z80.tv80s.i_tv80_core.I[0] ),
    .C(\z80.tv80s.i_tv80_core.I[3] ),
    .D(\z80.tv80s.i_tv80_core.I[2] ),
    .X(_2146_));
 sky130_fd_sc_hd__or4_1 _5275_ (.A(\z80.tv80s.i_tv80_core.I[5] ),
    .B(\z80.tv80s.i_tv80_core.I[4] ),
    .C(\z80.tv80s.i_tv80_core.I[6] ),
    .D(_2146_),
    .X(_2147_));
 sky130_fd_sc_hd__o31a_1 _5276_ (.A1(\z80.tv80s.i_tv80_core.I[7] ),
    .A2(_1625_),
    .A3(_2147_),
    .B1(_2145_),
    .X(_2148_));
 sky130_fd_sc_hd__mux2_1 _5277_ (.A0(_2143_),
    .A1(_2148_),
    .S(_1998_),
    .X(_2149_));
 sky130_fd_sc_hd__or4_1 _5278_ (.A(\z80.tv80s.di_reg[3] ),
    .B(\z80.tv80s.di_reg[2] ),
    .C(\z80.tv80s.di_reg[7] ),
    .D(\z80.tv80s.di_reg[6] ),
    .X(_2150_));
 sky130_fd_sc_hd__or4_1 _5279_ (.A(\z80.tv80s.di_reg[1] ),
    .B(\z80.tv80s.di_reg[0] ),
    .C(_2083_),
    .D(_2150_),
    .X(_2151_));
 sky130_fd_sc_hd__mux2_1 _5280_ (.A0(_2151_),
    .A1(_2149_),
    .S(_2022_),
    .X(_2152_));
 sky130_fd_sc_hd__mux2_1 _5281_ (.A0(_1245_),
    .A1(_2152_),
    .S(_1996_),
    .X(_2153_));
 sky130_fd_sc_hd__inv_2 _5282_ (.A(_2153_),
    .Y(_2154_));
 sky130_fd_sc_hd__mux2_1 _5283_ (.A0(net854),
    .A1(_2154_),
    .S(net116),
    .X(_0243_));
 sky130_fd_sc_hd__mux2_1 _5284_ (.A0(\z80.tv80s.i_tv80_core.F[7] ),
    .A1(_1270_),
    .S(_2870_),
    .X(_2155_));
 sky130_fd_sc_hd__mux2_1 _5285_ (.A0(\z80.tv80s.i_tv80_core.F[7] ),
    .A1(_1287_),
    .S(net119),
    .X(_2156_));
 sky130_fd_sc_hd__a22o_1 _5286_ (.A1(_2862_),
    .A2(_2155_),
    .B1(_2156_),
    .B2(_0839_),
    .X(_2157_));
 sky130_fd_sc_hd__a2111o_1 _5287_ (.A1(\z80.tv80s.i_tv80_core.F[7] ),
    .A2(_2077_),
    .B1(_2157_),
    .C1(_1284_),
    .D1(_1291_),
    .X(_2158_));
 sky130_fd_sc_hd__mux2_1 _5288_ (.A0(\z80.tv80s.i_tv80_core.F[7] ),
    .A1(\z80.tv80s.i_tv80_core.Fp[7] ),
    .S(_1502_),
    .X(_2159_));
 sky130_fd_sc_hd__mux2_1 _5289_ (.A0(_2159_),
    .A1(net792),
    .S(_1626_),
    .X(_2160_));
 sky130_fd_sc_hd__mux2_1 _5290_ (.A0(_2158_),
    .A1(_2160_),
    .S(_1998_),
    .X(_2161_));
 sky130_fd_sc_hd__mux2_1 _5291_ (.A0(\z80.tv80s.di_reg[7] ),
    .A1(_2161_),
    .S(_2022_),
    .X(_2162_));
 sky130_fd_sc_hd__mux2_1 _5292_ (.A0(_1295_),
    .A1(_2162_),
    .S(_1996_),
    .X(_2163_));
 sky130_fd_sc_hd__mux2_1 _5293_ (.A0(net833),
    .A1(_2163_),
    .S(net116),
    .X(_0244_));
 sky130_fd_sc_hd__or2_1 _5294_ (.A(_2861_),
    .B(_0713_),
    .X(_2164_));
 sky130_fd_sc_hd__and2_1 _5295_ (.A(_2856_),
    .B(_0741_),
    .X(_2165_));
 sky130_fd_sc_hd__or4b_4 _5296_ (.A(_0754_),
    .B(_0761_),
    .C(_2165_),
    .D_N(_0769_),
    .X(_2166_));
 sky130_fd_sc_hd__a21o_1 _5297_ (.A1(_2164_),
    .A2(_2166_),
    .B1(net125),
    .X(_2167_));
 sky130_fd_sc_hd__a21oi_1 _5298_ (.A1(_2143_),
    .A2(_2166_),
    .B1(_2167_),
    .Y(_2168_));
 sky130_fd_sc_hd__or3_1 _5299_ (.A(_0955_),
    .B(_0964_),
    .C(_2166_),
    .X(_2169_));
 sky130_fd_sc_hd__and4bb_1 _5300_ (.A_N(_2169_),
    .B_N(_0966_),
    .C(_0943_),
    .D(_1459_),
    .X(_2170_));
 sky130_fd_sc_hd__or4b_1 _5301_ (.A(_1464_),
    .B(_1470_),
    .C(_1477_),
    .D_N(_2170_),
    .X(_2171_));
 sky130_fd_sc_hd__or4_1 _5302_ (.A(_0978_),
    .B(_1024_),
    .C(_1484_),
    .D(_2171_),
    .X(_2172_));
 sky130_fd_sc_hd__or4b_1 _5303_ (.A(_1040_),
    .B(_1110_),
    .C(_2172_),
    .D_N(_1124_),
    .X(_2173_));
 sky130_fd_sc_hd__or4_2 _5304_ (.A(_1204_),
    .B(_1218_),
    .C(_1259_),
    .D(_2173_),
    .X(_2174_));
 sky130_fd_sc_hd__a22o_1 _5305_ (.A1(net429),
    .A2(_2167_),
    .B1(_2168_),
    .B2(_2174_),
    .X(_0245_));
 sky130_fd_sc_hd__a211o_1 _5306_ (.A1(net150),
    .A2(_2912_),
    .B1(_2917_),
    .C1(_2925_),
    .X(_2175_));
 sky130_fd_sc_hd__or4_1 _5307_ (.A(_2947_),
    .B(_0697_),
    .C(_0700_),
    .D(_2175_),
    .X(_2176_));
 sky130_fd_sc_hd__a211o_1 _5308_ (.A1(_2929_),
    .A2(_0477_),
    .B1(_0415_),
    .C1(_2962_),
    .X(_2177_));
 sky130_fd_sc_hd__or4_1 _5309_ (.A(_2909_),
    .B(_2914_),
    .C(_2942_),
    .D(_2177_),
    .X(_2178_));
 sky130_fd_sc_hd__or4_1 _5310_ (.A(_2926_),
    .B(_0412_),
    .C(_0425_),
    .D(_0701_),
    .X(_2179_));
 sky130_fd_sc_hd__or4_1 _5311_ (.A(_0509_),
    .B(_2176_),
    .C(_2178_),
    .D(_2179_),
    .X(_2180_));
 sky130_fd_sc_hd__a21o_1 _5312_ (.A1(_0397_),
    .A2(_0524_),
    .B1(_2180_),
    .X(_2181_));
 sky130_fd_sc_hd__a211o_1 _5313_ (.A1(net144),
    .A2(_2181_),
    .B1(_1318_),
    .C1(_1313_),
    .X(_2182_));
 sky130_fd_sc_hd__mux2_1 _5314_ (.A0(_0537_),
    .A1(_2849_),
    .S(net97),
    .X(_2183_));
 sky130_fd_sc_hd__nor2_1 _5315_ (.A(_2847_),
    .B(_2851_),
    .Y(_2184_));
 sky130_fd_sc_hd__nor2_1 _5316_ (.A(_2999_),
    .B(_0530_),
    .Y(_2185_));
 sky130_fd_sc_hd__nor2_1 _5317_ (.A(_2992_),
    .B(_0398_),
    .Y(_2186_));
 sky130_fd_sc_hd__o31a_1 _5318_ (.A1(_0671_),
    .A2(_2185_),
    .A3(_2186_),
    .B1(net146),
    .X(_2187_));
 sky130_fd_sc_hd__o41a_1 _5319_ (.A1(_3050_),
    .A2(_0392_),
    .A3(_0465_),
    .A4(_2187_),
    .B1(net106),
    .X(_2188_));
 sky130_fd_sc_hd__a221o_1 _5320_ (.A1(net166),
    .A2(_2182_),
    .B1(_2183_),
    .B2(_2184_),
    .C1(_2188_),
    .X(_2189_));
 sky130_fd_sc_hd__o2bb2a_1 _5321_ (.A1_N(net150),
    .A2_N(_2180_),
    .B1(_0525_),
    .B2(net131),
    .X(_2190_));
 sky130_fd_sc_hd__nor2_1 _5322_ (.A(net118),
    .B(_2190_),
    .Y(_2191_));
 sky130_fd_sc_hd__or4_1 _5323_ (.A(_2993_),
    .B(_3050_),
    .C(_0465_),
    .D(_0671_),
    .X(_2192_));
 sky130_fd_sc_hd__o32a_1 _5324_ (.A1(net152),
    .A2(_0678_),
    .A3(_1426_),
    .B1(_2185_),
    .B2(_2192_),
    .X(_2193_));
 sky130_fd_sc_hd__a211o_1 _5325_ (.A1(net152),
    .A2(_2991_),
    .B1(_0676_),
    .C1(_2193_),
    .X(_2194_));
 sky130_fd_sc_hd__a31o_1 _5326_ (.A1(_2916_),
    .A2(_2975_),
    .A3(_2987_),
    .B1(_3002_),
    .X(_2195_));
 sky130_fd_sc_hd__and4_1 _5327_ (.A(_3017_),
    .B(_3044_),
    .C(_3053_),
    .D(_2195_),
    .X(_2196_));
 sky130_fd_sc_hd__o2bb2a_1 _5328_ (.A1_N(_3000_),
    .A2_N(_2196_),
    .B1(net153),
    .B2(net137),
    .X(_2197_));
 sky130_fd_sc_hd__o21a_1 _5329_ (.A1(_2971_),
    .A2(_2980_),
    .B1(_0538_),
    .X(_2198_));
 sky130_fd_sc_hd__a211o_1 _5330_ (.A1(net153),
    .A2(_2183_),
    .B1(_2197_),
    .C1(_2198_),
    .X(_2199_));
 sky130_fd_sc_hd__a221o_1 _5331_ (.A1(net107),
    .A2(_2194_),
    .B1(_2199_),
    .B2(net824),
    .C1(_2191_),
    .X(_2200_));
 sky130_fd_sc_hd__and4bb_1 _5332_ (.A_N(net125),
    .B_N(_2189_),
    .C(\z80.tv80s.i_tv80_core.i_mcode.MCycle[2] ),
    .D(\z80.tv80s.i_tv80_core.ISet[1] ),
    .X(_2201_));
 sky130_fd_sc_hd__a22o_1 _5333_ (.A1(net125),
    .A2(net450),
    .B1(_2200_),
    .B2(_2201_),
    .X(_0246_));
 sky130_fd_sc_hd__nor2_2 _5334_ (.A(net125),
    .B(_2008_),
    .Y(_2202_));
 sky130_fd_sc_hd__a22o_1 _5335_ (.A1(net125),
    .A2(net839),
    .B1(_2200_),
    .B2(_2202_),
    .X(_0247_));
 sky130_fd_sc_hd__or2_1 _5336_ (.A(_1318_),
    .B(_2181_),
    .X(_2203_));
 sky130_fd_sc_hd__a221o_1 _5337_ (.A1(net161),
    .A2(_0433_),
    .B1(_2203_),
    .B2(net148),
    .C1(_3021_),
    .X(_2204_));
 sky130_fd_sc_hd__a31o_1 _5338_ (.A1(net152),
    .A2(_2991_),
    .A3(_0397_),
    .B1(_0465_),
    .X(_2205_));
 sky130_fd_sc_hd__o32a_1 _5339_ (.A1(_3050_),
    .A2(_0531_),
    .A3(_2205_),
    .B1(_1426_),
    .B2(net147),
    .X(_2206_));
 sky130_fd_sc_hd__o21a_1 _5340_ (.A1(\z80.tv80s.i_tv80_core.IR[4] ),
    .A2(_0398_),
    .B1(_2993_),
    .X(_2207_));
 sky130_fd_sc_hd__or2_1 _5341_ (.A(net147),
    .B(\z80.tv80s.i_tv80_core.i_mcode.MCycle[0] ),
    .X(_2208_));
 sky130_fd_sc_hd__a221o_1 _5342_ (.A1(net120),
    .A2(_0558_),
    .B1(_2208_),
    .B2(_3041_),
    .C1(_2207_),
    .X(_2209_));
 sky130_fd_sc_hd__o31a_1 _5343_ (.A1(_2999_),
    .A2(_2206_),
    .A3(_2209_),
    .B1(net107),
    .X(_2210_));
 sky130_fd_sc_hd__or3b_1 _5344_ (.A(_2926_),
    .B(_2950_),
    .C_N(_3032_),
    .X(_2211_));
 sky130_fd_sc_hd__or4_1 _5345_ (.A(_2914_),
    .B(_2942_),
    .C(_2947_),
    .D(_2211_),
    .X(_2212_));
 sky130_fd_sc_hd__or4_1 _5346_ (.A(_2948_),
    .B(_0425_),
    .C(_2175_),
    .D(_2212_),
    .X(_2213_));
 sky130_fd_sc_hd__o211a_1 _5347_ (.A1(net145),
    .A2(_2989_),
    .B1(_2987_),
    .C1(_2976_),
    .X(_2214_));
 sky130_fd_sc_hd__o311a_1 _5348_ (.A1(_2845_),
    .A2(_2937_),
    .A3(_2960_),
    .B1(_3006_),
    .C1(_3045_),
    .X(_2215_));
 sky130_fd_sc_hd__o31a_1 _5349_ (.A1(_2897_),
    .A2(_2995_),
    .A3(_2214_),
    .B1(_2215_),
    .X(_2216_));
 sky130_fd_sc_hd__nand2_1 _5350_ (.A(_2196_),
    .B(_2216_),
    .Y(_2217_));
 sky130_fd_sc_hd__o21a_1 _5351_ (.A1(_2213_),
    .A2(_2217_),
    .B1(_2208_),
    .X(_2218_));
 sky130_fd_sc_hd__a221o_1 _5352_ (.A1(\z80.tv80s.i_tv80_core.IR[7] ),
    .A2(_0538_),
    .B1(_2183_),
    .B2(net148),
    .C1(_2218_),
    .X(_2219_));
 sky130_fd_sc_hd__a221o_1 _5353_ (.A1(net166),
    .A2(_2204_),
    .B1(_2219_),
    .B2(net824),
    .C1(_2210_),
    .X(_2220_));
 sky130_fd_sc_hd__a22o_1 _5354_ (.A1(net125),
    .A2(net143),
    .B1(_2202_),
    .B2(net825),
    .X(_0248_));
 sky130_fd_sc_hd__a22o_1 _5355_ (.A1(net126),
    .A2(net832),
    .B1(_2189_),
    .B2(_2202_),
    .X(_0249_));
 sky130_fd_sc_hd__a21oi_1 _5356_ (.A1(_2982_),
    .A2(_0537_),
    .B1(_0568_),
    .Y(_2221_));
 sky130_fd_sc_hd__a211o_1 _5357_ (.A1(net166),
    .A2(_1314_),
    .B1(_2221_),
    .C1(net107),
    .X(_2222_));
 sky130_fd_sc_hd__a32o_1 _5358_ (.A1(_1330_),
    .A2(_2202_),
    .A3(_2222_),
    .B1(net805),
    .B2(net125),
    .X(_0250_));
 sky130_fd_sc_hd__o31a_1 _5359_ (.A1(_2970_),
    .A2(_3037_),
    .A3(_2217_),
    .B1(net137),
    .X(_2223_));
 sky130_fd_sc_hd__nor3_1 _5360_ (.A(_2980_),
    .B(_2983_),
    .C(_0537_),
    .Y(_2224_));
 sky130_fd_sc_hd__o21a_1 _5361_ (.A1(_2223_),
    .A2(_2224_),
    .B1(net824),
    .X(_2225_));
 sky130_fd_sc_hd__or4_1 _5362_ (.A(_0684_),
    .B(_1312_),
    .C(_1316_),
    .D(_1393_),
    .X(_2226_));
 sky130_fd_sc_hd__a211o_1 _5363_ (.A1(net875),
    .A2(_3041_),
    .B1(_0558_),
    .C1(_0678_),
    .X(_2227_));
 sky130_fd_sc_hd__or3_1 _5364_ (.A(_2999_),
    .B(_1426_),
    .C(_2227_),
    .X(_2228_));
 sky130_fd_sc_hd__a221o_1 _5365_ (.A1(net166),
    .A2(_2226_),
    .B1(_2228_),
    .B2(net107),
    .C1(_2225_),
    .X(_2229_));
 sky130_fd_sc_hd__a22o_1 _5366_ (.A1(net126),
    .A2(net837),
    .B1(_2202_),
    .B2(_2229_),
    .X(_0251_));
 sky130_fd_sc_hd__nor2_1 _5367_ (.A(\z80.tv80s.i_tv80_core.No_BTR ),
    .B(_0673_),
    .Y(_2230_));
 sky130_fd_sc_hd__mux2_1 _5368_ (.A0(net263),
    .A1(_2230_),
    .S(_2202_),
    .X(_0252_));
 sky130_fd_sc_hd__or4_1 _5369_ (.A(_2926_),
    .B(_2929_),
    .C(_2943_),
    .D(_0412_),
    .X(_2231_));
 sky130_fd_sc_hd__or4_1 _5370_ (.A(_2965_),
    .B(_0422_),
    .C(_0443_),
    .D(_1390_),
    .X(_2232_));
 sky130_fd_sc_hd__or4_1 _5371_ (.A(_2925_),
    .B(_2944_),
    .C(_0507_),
    .D(_2232_),
    .X(_2233_));
 sky130_fd_sc_hd__or4_1 _5372_ (.A(_0505_),
    .B(_0706_),
    .C(_2231_),
    .D(_2233_),
    .X(_2234_));
 sky130_fd_sc_hd__nor2_1 _5373_ (.A(_0704_),
    .B(_2234_),
    .Y(_2235_));
 sky130_fd_sc_hd__and3_1 _5374_ (.A(\z80.tv80s.i_tv80_core.i_mcode.MCycle[3] ),
    .B(_3026_),
    .C(_0474_),
    .X(_2236_));
 sky130_fd_sc_hd__a31o_1 _5375_ (.A1(net152),
    .A2(_2912_),
    .A3(_0512_),
    .B1(_2236_),
    .X(_2237_));
 sky130_fd_sc_hd__mux2_1 _5376_ (.A0(_2237_),
    .A1(net131),
    .S(_2235_),
    .X(_2238_));
 sky130_fd_sc_hd__a22oi_4 _5377_ (.A1(_2999_),
    .A2(net106),
    .B1(_2238_),
    .B2(net164),
    .Y(_2239_));
 sky130_fd_sc_hd__a21oi_1 _5378_ (.A1(_1525_),
    .A2(_2239_),
    .B1(net60),
    .Y(_2240_));
 sky130_fd_sc_hd__mux2_1 _5379_ (.A0(net633),
    .A1(_2240_),
    .S(net113),
    .X(_0253_));
 sky130_fd_sc_hd__a21oi_1 _5380_ (.A1(_1333_),
    .A2(_2239_),
    .B1(net60),
    .Y(_2241_));
 sky130_fd_sc_hd__mux2_1 _5381_ (.A0(net508),
    .A1(_2241_),
    .S(net113),
    .X(_0254_));
 sky130_fd_sc_hd__a21oi_1 _5382_ (.A1(_1349_),
    .A2(_2239_),
    .B1(net60),
    .Y(_2242_));
 sky130_fd_sc_hd__mux2_1 _5383_ (.A0(net501),
    .A1(_2242_),
    .S(net114),
    .X(_0255_));
 sky130_fd_sc_hd__nor2_1 _5384_ (.A(net124),
    .B(_1506_),
    .Y(_2243_));
 sky130_fd_sc_hd__a32o_1 _5385_ (.A1(_0577_),
    .A2(_2239_),
    .A3(_2243_),
    .B1(net464),
    .B2(\z80.tv80s.i_tv80_core.BusAck ),
    .X(_0256_));
 sky130_fd_sc_hd__nor2_1 _5386_ (.A(net114),
    .B(_2875_),
    .Y(_2244_));
 sky130_fd_sc_hd__or3_1 _5387_ (.A(net110),
    .B(_2918_),
    .C(_0397_),
    .X(_2245_));
 sky130_fd_sc_hd__or4b_1 _5388_ (.A(net109),
    .B(_1312_),
    .C(_1322_),
    .D_N(_2245_),
    .X(_2246_));
 sky130_fd_sc_hd__o41a_1 _5389_ (.A1(_1316_),
    .A2(_1339_),
    .A3(_1393_),
    .A4(_2246_),
    .B1(_1311_),
    .X(_2247_));
 sky130_fd_sc_hd__o31a_1 _5390_ (.A1(_1328_),
    .A2(_1331_),
    .A3(_2227_),
    .B1(net106),
    .X(_2248_));
 sky130_fd_sc_hd__or4b_1 _5391_ (.A(_2225_),
    .B(_2247_),
    .C(_2248_),
    .D_N(_2239_),
    .X(_2249_));
 sky130_fd_sc_hd__a31o_1 _5392_ (.A1(net114),
    .A2(_0577_),
    .A3(_2249_),
    .B1(_2244_),
    .X(_0257_));
 sky130_fd_sc_hd__a22o_1 _5393_ (.A1(net126),
    .A2(net625),
    .B1(_0624_),
    .B2(_0684_),
    .X(_0258_));
 sky130_fd_sc_hd__a31o_1 _5394_ (.A1(_2859_),
    .A2(net103),
    .A3(_1412_),
    .B1(_1401_),
    .X(_2250_));
 sky130_fd_sc_hd__mux2_1 _5395_ (.A0(net142),
    .A1(_2250_),
    .S(net113),
    .X(_0259_));
 sky130_fd_sc_hd__mux2_1 _5396_ (.A0(net542),
    .A1(_1412_),
    .S(net114),
    .X(_0260_));
 sky130_fd_sc_hd__a21oi_1 _5397_ (.A1(\z80.tv80s.i_tv80_core.i_mcode.MCycle[5] ),
    .A2(_0602_),
    .B1(net534),
    .Y(_2251_));
 sky130_fd_sc_hd__or2_1 _5398_ (.A(_2934_),
    .B(_0611_),
    .X(_2252_));
 sky130_fd_sc_hd__a21oi_1 _5399_ (.A1(_0608_),
    .A2(_2252_),
    .B1(net535),
    .Y(_0261_));
 sky130_fd_sc_hd__or2_1 _5400_ (.A(_0600_),
    .B(_0609_),
    .X(_2253_));
 sky130_fd_sc_hd__a22o_1 _5401_ (.A1(_2847_),
    .A2(_0627_),
    .B1(_2253_),
    .B2(net467),
    .X(_0262_));
 sky130_fd_sc_hd__a22o_1 _5402_ (.A1(net96),
    .A2(_0627_),
    .B1(_2253_),
    .B2(net566),
    .X(_0263_));
 sky130_fd_sc_hd__o21ai_1 _5403_ (.A1(_0459_),
    .A2(_1419_),
    .B1(_1420_),
    .Y(_2254_));
 sky130_fd_sc_hd__mux2_1 _5404_ (.A0(net139),
    .A1(_2254_),
    .S(net114),
    .X(_0264_));
 sky130_fd_sc_hd__nand2_1 _5405_ (.A(_0391_),
    .B(_0463_),
    .Y(_2255_));
 sky130_fd_sc_hd__nor2_1 _5406_ (.A(net134),
    .B(_0424_),
    .Y(_2256_));
 sky130_fd_sc_hd__or4b_1 _5407_ (.A(_0416_),
    .B(_2256_),
    .C(_0439_),
    .D_N(_0442_),
    .X(_2257_));
 sky130_fd_sc_hd__a22o_1 _5408_ (.A1(_0555_),
    .A2(_0623_),
    .B1(_2257_),
    .B2(net131),
    .X(_2258_));
 sky130_fd_sc_hd__a32o_1 _5409_ (.A1(\z80.tv80s.i_tv80_core.i_mcode.MCycle[1] ),
    .A2(net107),
    .A3(_2255_),
    .B1(_2258_),
    .B2(net166),
    .X(_2259_));
 sky130_fd_sc_hd__nand2_4 _5410_ (.A(net736),
    .B(_2259_),
    .Y(_2260_));
 sky130_fd_sc_hd__nor2_1 _5411_ (.A(_2854_),
    .B(_2872_),
    .Y(_2261_));
 sky130_fd_sc_hd__a22o_1 _5412_ (.A1(_2854_),
    .A2(\z80.tv80s.i_tv80_core.SP[0] ),
    .B1(_1673_),
    .B2(_2261_),
    .X(_2262_));
 sky130_fd_sc_hd__nor2_1 _5413_ (.A(\z80.tv80s.di_reg[0] ),
    .B(_1673_),
    .Y(_2263_));
 sky130_fd_sc_hd__a21oi_1 _5414_ (.A1(net122),
    .A2(_2263_),
    .B1(_2262_),
    .Y(_2264_));
 sky130_fd_sc_hd__and2_2 _5415_ (.A(\z80.tv80s.i_tv80_core.i_mcode.MCycle[5] ),
    .B(\z80.tv80s.i_tv80_core.ts[3] ),
    .X(_2265_));
 sky130_fd_sc_hd__nand2_4 _5416_ (.A(\z80.tv80s.i_tv80_core.i_mcode.MCycle[5] ),
    .B(net122),
    .Y(_2266_));
 sky130_fd_sc_hd__nor2_1 _5417_ (.A(net100),
    .B(_2266_),
    .Y(_2267_));
 sky130_fd_sc_hd__and3_4 _5418_ (.A(_0603_),
    .B(_1566_),
    .C(_1571_),
    .X(_2268_));
 sky130_fd_sc_hd__mux2_1 _5419_ (.A0(net801),
    .A1(net13),
    .S(_2268_),
    .X(_2269_));
 sky130_fd_sc_hd__a22o_1 _5420_ (.A1(_2264_),
    .A2(_2267_),
    .B1(_2269_),
    .B2(net101),
    .X(_2270_));
 sky130_fd_sc_hd__mux2_1 _5421_ (.A0(\z80.tv80s.di_reg[0] ),
    .A1(_2270_),
    .S(_2260_),
    .X(_2271_));
 sky130_fd_sc_hd__or2_2 _5422_ (.A(_0604_),
    .B(_1677_),
    .X(_2272_));
 sky130_fd_sc_hd__and2_4 _5423_ (.A(_2266_),
    .B(_2272_),
    .X(_2273_));
 sky130_fd_sc_hd__a31o_1 _5424_ (.A1(net94),
    .A2(_2260_),
    .A3(_2273_),
    .B1(net128),
    .X(_2274_));
 sky130_fd_sc_hd__a22o_1 _5425_ (.A1(net116),
    .A2(_2271_),
    .B1(_2274_),
    .B2(net801),
    .X(_0265_));
 sky130_fd_sc_hd__a311o_4 _5426_ (.A1(net106),
    .A2(_0864_),
    .A3(_0865_),
    .B1(_0863_),
    .C1(net122),
    .X(_2275_));
 sky130_fd_sc_hd__nand2_1 _5427_ (.A(\z80.tv80s.i_tv80_core.ts[3] ),
    .B(_2871_),
    .Y(_2276_));
 sky130_fd_sc_hd__mux2_1 _5428_ (.A0(\z80.tv80s.i_tv80_core.SP[1] ),
    .A1(_1715_),
    .S(net122),
    .X(_2277_));
 sky130_fd_sc_hd__and3_1 _5429_ (.A(_2275_),
    .B(_2276_),
    .C(_2277_),
    .X(_2278_));
 sky130_fd_sc_hd__a21o_1 _5430_ (.A1(_2275_),
    .A2(_2276_),
    .B1(_2277_),
    .X(_2279_));
 sky130_fd_sc_hd__and2b_1 _5431_ (.A_N(_2278_),
    .B(_2279_),
    .X(_2280_));
 sky130_fd_sc_hd__xnor2_1 _5432_ (.A(_2262_),
    .B(_2280_),
    .Y(_2281_));
 sky130_fd_sc_hd__inv_2 _5433_ (.A(_2281_),
    .Y(_2282_));
 sky130_fd_sc_hd__a22o_1 _5434_ (.A1(net790),
    .A2(_2273_),
    .B1(_2282_),
    .B2(_2265_),
    .X(_2283_));
 sky130_fd_sc_hd__mux2_1 _5435_ (.A0(net790),
    .A1(net12),
    .S(_2268_),
    .X(_2284_));
 sky130_fd_sc_hd__mux2_1 _5436_ (.A0(_2283_),
    .A1(_2284_),
    .S(_0598_),
    .X(_2285_));
 sky130_fd_sc_hd__mux2_1 _5437_ (.A0(\z80.tv80s.di_reg[1] ),
    .A1(_2285_),
    .S(_2260_),
    .X(_2286_));
 sky130_fd_sc_hd__mux2_1 _5438_ (.A0(net790),
    .A1(_2286_),
    .S(net116),
    .X(_0266_));
 sky130_fd_sc_hd__or2_1 _5439_ (.A(_2854_),
    .B(\z80.tv80s.di_reg[2] ),
    .X(_2287_));
 sky130_fd_sc_hd__mux2_1 _5440_ (.A0(\z80.tv80s.i_tv80_core.SP[2] ),
    .A1(_1736_),
    .S(net121),
    .X(_2288_));
 sky130_fd_sc_hd__and3_1 _5441_ (.A(_2275_),
    .B(_2287_),
    .C(_2288_),
    .X(_2289_));
 sky130_fd_sc_hd__a21oi_1 _5442_ (.A1(_2275_),
    .A2(_2287_),
    .B1(_2288_),
    .Y(_2290_));
 sky130_fd_sc_hd__nor2_1 _5443_ (.A(_2289_),
    .B(_2290_),
    .Y(_2291_));
 sky130_fd_sc_hd__a21o_1 _5444_ (.A1(_2262_),
    .A2(_2279_),
    .B1(_2278_),
    .X(_2292_));
 sky130_fd_sc_hd__xor2_1 _5445_ (.A(_2291_),
    .B(_2292_),
    .X(_2293_));
 sky130_fd_sc_hd__a22o_1 _5446_ (.A1(net803),
    .A2(_2273_),
    .B1(_2293_),
    .B2(_2265_),
    .X(_2294_));
 sky130_fd_sc_hd__mux2_1 _5447_ (.A0(net803),
    .A1(net10),
    .S(_2268_),
    .X(_2295_));
 sky130_fd_sc_hd__mux2_1 _5448_ (.A0(_2294_),
    .A1(_2295_),
    .S(_0598_),
    .X(_2296_));
 sky130_fd_sc_hd__mux2_1 _5449_ (.A0(\z80.tv80s.di_reg[2] ),
    .A1(_2296_),
    .S(_2260_),
    .X(_2297_));
 sky130_fd_sc_hd__mux2_1 _5450_ (.A0(net803),
    .A1(_2297_),
    .S(net116),
    .X(_0267_));
 sky130_fd_sc_hd__or2_1 _5451_ (.A(_2854_),
    .B(\z80.tv80s.di_reg[3] ),
    .X(_2298_));
 sky130_fd_sc_hd__mux2_1 _5452_ (.A0(\z80.tv80s.i_tv80_core.SP[3] ),
    .A1(_1754_),
    .S(net121),
    .X(_2299_));
 sky130_fd_sc_hd__nand3_1 _5453_ (.A(_2275_),
    .B(_2298_),
    .C(_2299_),
    .Y(_2300_));
 sky130_fd_sc_hd__a21o_1 _5454_ (.A1(_2275_),
    .A2(_2298_),
    .B1(_2299_),
    .X(_2301_));
 sky130_fd_sc_hd__and2_1 _5455_ (.A(_2300_),
    .B(_2301_),
    .X(_2302_));
 sky130_fd_sc_hd__a21o_1 _5456_ (.A1(_2291_),
    .A2(_2292_),
    .B1(_2289_),
    .X(_2303_));
 sky130_fd_sc_hd__xor2_1 _5457_ (.A(_2302_),
    .B(_2303_),
    .X(_2304_));
 sky130_fd_sc_hd__mux2_1 _5458_ (.A0(net154),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[3] ),
    .S(_2272_),
    .X(_2305_));
 sky130_fd_sc_hd__mux2_1 _5459_ (.A0(_2304_),
    .A1(_2305_),
    .S(_2266_),
    .X(_2306_));
 sky130_fd_sc_hd__mux2_1 _5460_ (.A0(net827),
    .A1(net7),
    .S(_2268_),
    .X(_2307_));
 sky130_fd_sc_hd__mux2_1 _5461_ (.A0(_2306_),
    .A1(_2307_),
    .S(net101),
    .X(_2308_));
 sky130_fd_sc_hd__mux2_1 _5462_ (.A0(\z80.tv80s.di_reg[3] ),
    .A1(_2308_),
    .S(_2260_),
    .X(_2309_));
 sky130_fd_sc_hd__mux2_1 _5463_ (.A0(net827),
    .A1(_2309_),
    .S(net114),
    .X(_0268_));
 sky130_fd_sc_hd__or2_1 _5464_ (.A(_2854_),
    .B(\z80.tv80s.di_reg[4] ),
    .X(_2310_));
 sky130_fd_sc_hd__mux2_1 _5465_ (.A0(\z80.tv80s.i_tv80_core.SP[4] ),
    .A1(_1771_),
    .S(net121),
    .X(_2311_));
 sky130_fd_sc_hd__nand3_1 _5466_ (.A(_2275_),
    .B(_2310_),
    .C(_2311_),
    .Y(_2312_));
 sky130_fd_sc_hd__a21o_1 _5467_ (.A1(_2275_),
    .A2(_2310_),
    .B1(_2311_),
    .X(_2313_));
 sky130_fd_sc_hd__and2_1 _5468_ (.A(_2312_),
    .B(_2313_),
    .X(_2314_));
 sky130_fd_sc_hd__a21bo_1 _5469_ (.A1(_2301_),
    .A2(_2303_),
    .B1_N(_2300_),
    .X(_2315_));
 sky130_fd_sc_hd__xor2_2 _5470_ (.A(_2314_),
    .B(_2315_),
    .X(_2316_));
 sky130_fd_sc_hd__mux2_1 _5471_ (.A0(net147),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[4] ),
    .S(_2272_),
    .X(_2317_));
 sky130_fd_sc_hd__mux2_1 _5472_ (.A0(_2316_),
    .A1(_2317_),
    .S(_2266_),
    .X(_2318_));
 sky130_fd_sc_hd__mux2_1 _5473_ (.A0(net815),
    .A1(net6),
    .S(_2268_),
    .X(_2319_));
 sky130_fd_sc_hd__mux2_1 _5474_ (.A0(_2318_),
    .A1(_2319_),
    .S(net101),
    .X(_2320_));
 sky130_fd_sc_hd__mux2_1 _5475_ (.A0(\z80.tv80s.di_reg[4] ),
    .A1(_2320_),
    .S(_2260_),
    .X(_2321_));
 sky130_fd_sc_hd__mux2_1 _5476_ (.A0(net815),
    .A1(_2321_),
    .S(net114),
    .X(_0269_));
 sky130_fd_sc_hd__or2_1 _5477_ (.A(_2854_),
    .B(\z80.tv80s.di_reg[5] ),
    .X(_2322_));
 sky130_fd_sc_hd__mux2_1 _5478_ (.A0(\z80.tv80s.i_tv80_core.SP[5] ),
    .A1(_1789_),
    .S(net122),
    .X(_2323_));
 sky130_fd_sc_hd__and3_1 _5479_ (.A(_2275_),
    .B(_2322_),
    .C(_2323_),
    .X(_2324_));
 sky130_fd_sc_hd__a21oi_1 _5480_ (.A1(_2275_),
    .A2(_2322_),
    .B1(_2323_),
    .Y(_2325_));
 sky130_fd_sc_hd__nor2_1 _5481_ (.A(_2324_),
    .B(_2325_),
    .Y(_2326_));
 sky130_fd_sc_hd__a21bo_1 _5482_ (.A1(_2313_),
    .A2(_2315_),
    .B1_N(_2312_),
    .X(_2327_));
 sky130_fd_sc_hd__xor2_2 _5483_ (.A(_2326_),
    .B(_2327_),
    .X(_2328_));
 sky130_fd_sc_hd__mux2_1 _5484_ (.A0(net146),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[5] ),
    .S(_2272_),
    .X(_2329_));
 sky130_fd_sc_hd__mux2_1 _5485_ (.A0(_2328_),
    .A1(_2329_),
    .S(_2266_),
    .X(_2330_));
 sky130_fd_sc_hd__mux2_1 _5486_ (.A0(net821),
    .A1(net8),
    .S(_2268_),
    .X(_2331_));
 sky130_fd_sc_hd__mux2_1 _5487_ (.A0(_2330_),
    .A1(_2331_),
    .S(net101),
    .X(_2332_));
 sky130_fd_sc_hd__mux2_1 _5488_ (.A0(\z80.tv80s.di_reg[5] ),
    .A1(_2332_),
    .S(_2260_),
    .X(_2333_));
 sky130_fd_sc_hd__mux2_1 _5489_ (.A0(net821),
    .A1(_2333_),
    .S(net116),
    .X(_0270_));
 sky130_fd_sc_hd__or2_1 _5490_ (.A(_2854_),
    .B(\z80.tv80s.di_reg[6] ),
    .X(_2334_));
 sky130_fd_sc_hd__mux2_1 _5491_ (.A0(\z80.tv80s.i_tv80_core.SP[6] ),
    .A1(_1807_),
    .S(net121),
    .X(_2335_));
 sky130_fd_sc_hd__and3_1 _5492_ (.A(_2275_),
    .B(_2334_),
    .C(_2335_),
    .X(_2336_));
 sky130_fd_sc_hd__a21oi_1 _5493_ (.A1(_2275_),
    .A2(_2334_),
    .B1(_2335_),
    .Y(_2337_));
 sky130_fd_sc_hd__nor2_1 _5494_ (.A(_2336_),
    .B(_2337_),
    .Y(_2338_));
 sky130_fd_sc_hd__a21oi_1 _5495_ (.A1(_2326_),
    .A2(_2327_),
    .B1(_2324_),
    .Y(_2339_));
 sky130_fd_sc_hd__xnor2_1 _5496_ (.A(_2338_),
    .B(_2339_),
    .Y(_2340_));
 sky130_fd_sc_hd__a22o_1 _5497_ (.A1(net810),
    .A2(_2273_),
    .B1(_2340_),
    .B2(_2265_),
    .X(_2341_));
 sky130_fd_sc_hd__mux2_1 _5498_ (.A0(net810),
    .A1(net9),
    .S(_2268_),
    .X(_2342_));
 sky130_fd_sc_hd__mux2_1 _5499_ (.A0(_2341_),
    .A1(_2342_),
    .S(_0598_),
    .X(_2343_));
 sky130_fd_sc_hd__mux2_1 _5500_ (.A0(\z80.tv80s.di_reg[6] ),
    .A1(_2343_),
    .S(_2260_),
    .X(_2344_));
 sky130_fd_sc_hd__mux2_1 _5501_ (.A0(net810),
    .A1(_2344_),
    .S(net114),
    .X(_0271_));
 sky130_fd_sc_hd__o21ba_1 _5502_ (.A1(_2337_),
    .A2(_2339_),
    .B1_N(_2336_),
    .X(_2345_));
 sky130_fd_sc_hd__o21a_1 _5503_ (.A1(_2854_),
    .A2(\z80.tv80s.di_reg[7] ),
    .B1(_2275_),
    .X(_2346_));
 sky130_fd_sc_hd__mux2_1 _5504_ (.A0(\z80.tv80s.i_tv80_core.SP[7] ),
    .A1(_1828_),
    .S(net121),
    .X(_2347_));
 sky130_fd_sc_hd__nor2_1 _5505_ (.A(net72),
    .B(_2347_),
    .Y(_2348_));
 sky130_fd_sc_hd__nand2_1 _5506_ (.A(net72),
    .B(_2347_),
    .Y(_2349_));
 sky130_fd_sc_hd__nand2b_1 _5507_ (.A_N(_2348_),
    .B(_2349_),
    .Y(_2350_));
 sky130_fd_sc_hd__xnor2_2 _5508_ (.A(_2345_),
    .B(_2350_),
    .Y(_2351_));
 sky130_fd_sc_hd__o2bb2ai_1 _5509_ (.A1_N(net812),
    .A2_N(_2273_),
    .B1(_2351_),
    .B2(_2266_),
    .Y(_2352_));
 sky130_fd_sc_hd__mux2_1 _5510_ (.A0(net812),
    .A1(net11),
    .S(_2268_),
    .X(_2353_));
 sky130_fd_sc_hd__mux2_1 _5511_ (.A0(_2352_),
    .A1(_2353_),
    .S(net101),
    .X(_2354_));
 sky130_fd_sc_hd__mux2_1 _5512_ (.A0(\z80.tv80s.di_reg[7] ),
    .A1(_2354_),
    .S(_2260_),
    .X(_2355_));
 sky130_fd_sc_hd__mux2_1 _5513_ (.A0(net812),
    .A1(_2355_),
    .S(net114),
    .X(_0272_));
 sky130_fd_sc_hd__o21a_1 _5514_ (.A1(_2345_),
    .A2(_2348_),
    .B1(_2349_),
    .X(_2356_));
 sky130_fd_sc_hd__mux2_1 _5515_ (.A0(\z80.tv80s.i_tv80_core.SP[8] ),
    .A1(_1847_),
    .S(net121),
    .X(_2357_));
 sky130_fd_sc_hd__nand2_1 _5516_ (.A(net72),
    .B(_2357_),
    .Y(_2358_));
 sky130_fd_sc_hd__or2_1 _5517_ (.A(net72),
    .B(_2357_),
    .X(_2359_));
 sky130_fd_sc_hd__nand2_1 _5518_ (.A(_2358_),
    .B(_2359_),
    .Y(_2360_));
 sky130_fd_sc_hd__xnor2_1 _5519_ (.A(_2356_),
    .B(_2360_),
    .Y(_2361_));
 sky130_fd_sc_hd__or2_1 _5520_ (.A(net100),
    .B(_2273_),
    .X(_2362_));
 sky130_fd_sc_hd__nand2_1 _5521_ (.A(net593),
    .B(_2362_),
    .Y(_2363_));
 sky130_fd_sc_hd__and4_1 _5522_ (.A(net165),
    .B(_2924_),
    .C(_0508_),
    .D(_0512_),
    .X(_2364_));
 sky130_fd_sc_hd__or4b_4 _5523_ (.A(_0697_),
    .B(_1679_),
    .C(_2231_),
    .D_N(_2364_),
    .X(_2365_));
 sky130_fd_sc_hd__o21ai_4 _5524_ (.A1(_0391_),
    .A2(_0670_),
    .B1(_2365_),
    .Y(_2366_));
 sky130_fd_sc_hd__nand2_4 _5525_ (.A(net121),
    .B(_2366_),
    .Y(_2367_));
 sky130_fd_sc_hd__o311a_1 _5526_ (.A1(net100),
    .A2(_2266_),
    .A3(_2361_),
    .B1(_2363_),
    .C1(_2367_),
    .X(_2368_));
 sky130_fd_sc_hd__a31o_1 _5527_ (.A1(net121),
    .A2(_2872_),
    .A3(_2366_),
    .B1(net128),
    .X(_2369_));
 sky130_fd_sc_hd__a2bb2o_1 _5528_ (.A1_N(_2368_),
    .A2_N(_2369_),
    .B1(net128),
    .B2(net593),
    .X(_0273_));
 sky130_fd_sc_hd__mux2_1 _5529_ (.A0(\z80.tv80s.i_tv80_core.SP[9] ),
    .A1(_1866_),
    .S(net121),
    .X(_2370_));
 sky130_fd_sc_hd__nor2_1 _5530_ (.A(net72),
    .B(_2370_),
    .Y(_2371_));
 sky130_fd_sc_hd__and2_1 _5531_ (.A(_2346_),
    .B(_2370_),
    .X(_2372_));
 sky130_fd_sc_hd__nor2_1 _5532_ (.A(_2371_),
    .B(_2372_),
    .Y(_2373_));
 sky130_fd_sc_hd__o21a_1 _5533_ (.A1(_2356_),
    .A2(_2360_),
    .B1(_2358_),
    .X(_2374_));
 sky130_fd_sc_hd__xnor2_1 _5534_ (.A(_2373_),
    .B(_2374_),
    .Y(_2375_));
 sky130_fd_sc_hd__a22o_1 _5535_ (.A1(net611),
    .A2(_2362_),
    .B1(_2375_),
    .B2(_2267_),
    .X(_2376_));
 sky130_fd_sc_hd__mux2_1 _5536_ (.A0(\z80.tv80s.di_reg[1] ),
    .A1(_2376_),
    .S(_2367_),
    .X(_2377_));
 sky130_fd_sc_hd__mux2_1 _5537_ (.A0(net611),
    .A1(_2377_),
    .S(net117),
    .X(_0274_));
 sky130_fd_sc_hd__o21ai_1 _5538_ (.A1(_2357_),
    .A2(_2370_),
    .B1(_2346_),
    .Y(_2378_));
 sky130_fd_sc_hd__o41a_1 _5539_ (.A1(_2356_),
    .A2(_2360_),
    .A3(_2371_),
    .A4(_2372_),
    .B1(_2378_),
    .X(_2379_));
 sky130_fd_sc_hd__mux2_1 _5540_ (.A0(\z80.tv80s.i_tv80_core.SP[10] ),
    .A1(_1885_),
    .S(net121),
    .X(_2380_));
 sky130_fd_sc_hd__nand2_1 _5541_ (.A(net72),
    .B(_2380_),
    .Y(_2381_));
 sky130_fd_sc_hd__or2_1 _5542_ (.A(net72),
    .B(_2380_),
    .X(_2382_));
 sky130_fd_sc_hd__and2_1 _5543_ (.A(_2381_),
    .B(_2382_),
    .X(_2383_));
 sky130_fd_sc_hd__inv_2 _5544_ (.A(_2383_),
    .Y(_2384_));
 sky130_fd_sc_hd__xnor2_1 _5545_ (.A(_2379_),
    .B(_2383_),
    .Y(_2385_));
 sky130_fd_sc_hd__a22o_1 _5546_ (.A1(net761),
    .A2(_2273_),
    .B1(_2385_),
    .B2(_2265_),
    .X(_2386_));
 sky130_fd_sc_hd__mux2_1 _5547_ (.A0(net761),
    .A1(_2386_),
    .S(net93),
    .X(_2387_));
 sky130_fd_sc_hd__mux2_1 _5548_ (.A0(\z80.tv80s.di_reg[2] ),
    .A1(_2387_),
    .S(_2367_),
    .X(_2388_));
 sky130_fd_sc_hd__mux2_1 _5549_ (.A0(net761),
    .A1(_2388_),
    .S(net117),
    .X(_0275_));
 sky130_fd_sc_hd__mux2_1 _5550_ (.A0(\z80.tv80s.i_tv80_core.SP[11] ),
    .A1(_1903_),
    .S(net121),
    .X(_2389_));
 sky130_fd_sc_hd__xnor2_1 _5551_ (.A(net72),
    .B(_2389_),
    .Y(_2390_));
 sky130_fd_sc_hd__o21a_1 _5552_ (.A1(_2379_),
    .A2(_2384_),
    .B1(_2381_),
    .X(_2391_));
 sky130_fd_sc_hd__xnor2_1 _5553_ (.A(_2390_),
    .B(_2391_),
    .Y(_2392_));
 sky130_fd_sc_hd__inv_2 _5554_ (.A(_2392_),
    .Y(_2393_));
 sky130_fd_sc_hd__a22o_1 _5555_ (.A1(net776),
    .A2(_2273_),
    .B1(_2393_),
    .B2(_2265_),
    .X(_2394_));
 sky130_fd_sc_hd__mux2_1 _5556_ (.A0(net776),
    .A1(_2394_),
    .S(net93),
    .X(_2395_));
 sky130_fd_sc_hd__mux2_1 _5557_ (.A0(\z80.tv80s.di_reg[3] ),
    .A1(_2395_),
    .S(_2367_),
    .X(_2396_));
 sky130_fd_sc_hd__mux2_1 _5558_ (.A0(net776),
    .A1(_2396_),
    .S(net112),
    .X(_0276_));
 sky130_fd_sc_hd__mux2_1 _5559_ (.A0(\z80.tv80s.i_tv80_core.SP[12] ),
    .A1(_1922_),
    .S(net121),
    .X(_2397_));
 sky130_fd_sc_hd__and2_1 _5560_ (.A(net72),
    .B(_2397_),
    .X(_2398_));
 sky130_fd_sc_hd__nor2_1 _5561_ (.A(net72),
    .B(_2397_),
    .Y(_2399_));
 sky130_fd_sc_hd__or2_1 _5562_ (.A(_2398_),
    .B(_2399_),
    .X(_2400_));
 sky130_fd_sc_hd__o21ai_1 _5563_ (.A1(_2380_),
    .A2(_2389_),
    .B1(net72),
    .Y(_2401_));
 sky130_fd_sc_hd__o31a_1 _5564_ (.A1(_2379_),
    .A2(_2384_),
    .A3(_2390_),
    .B1(_2401_),
    .X(_2402_));
 sky130_fd_sc_hd__xnor2_1 _5565_ (.A(_2400_),
    .B(_2402_),
    .Y(_2403_));
 sky130_fd_sc_hd__o2bb2a_1 _5566_ (.A1_N(\z80.tv80s.i_tv80_core.TmpAddr[12] ),
    .A2_N(_2273_),
    .B1(_2403_),
    .B2(_2266_),
    .X(_2404_));
 sky130_fd_sc_hd__nand2_1 _5567_ (.A(net753),
    .B(net101),
    .Y(_2405_));
 sky130_fd_sc_hd__o211a_1 _5568_ (.A1(net101),
    .A2(_2404_),
    .B1(_2405_),
    .C1(_2367_),
    .X(_2406_));
 sky130_fd_sc_hd__o21ba_1 _5569_ (.A1(\z80.tv80s.di_reg[4] ),
    .A2(_2367_),
    .B1_N(_2406_),
    .X(_2407_));
 sky130_fd_sc_hd__mux2_1 _5570_ (.A0(net753),
    .A1(_2407_),
    .S(net117),
    .X(_0277_));
 sky130_fd_sc_hd__mux2_1 _5571_ (.A0(\z80.tv80s.i_tv80_core.SP[13] ),
    .A1(_1943_),
    .S(net121),
    .X(_2408_));
 sky130_fd_sc_hd__nand2_1 _5572_ (.A(net72),
    .B(_2408_),
    .Y(_2409_));
 sky130_fd_sc_hd__or2_1 _5573_ (.A(net72),
    .B(_2408_),
    .X(_2410_));
 sky130_fd_sc_hd__nand2_1 _5574_ (.A(_2409_),
    .B(_2410_),
    .Y(_2411_));
 sky130_fd_sc_hd__o21ba_1 _5575_ (.A1(_2399_),
    .A2(_2402_),
    .B1_N(_2398_),
    .X(_2412_));
 sky130_fd_sc_hd__xnor2_1 _5576_ (.A(_2411_),
    .B(_2412_),
    .Y(_2413_));
 sky130_fd_sc_hd__inv_2 _5577_ (.A(_2413_),
    .Y(_2414_));
 sky130_fd_sc_hd__a22o_1 _5578_ (.A1(net782),
    .A2(_2273_),
    .B1(_2414_),
    .B2(_2265_),
    .X(_2415_));
 sky130_fd_sc_hd__mux2_1 _5579_ (.A0(net782),
    .A1(_2415_),
    .S(net93),
    .X(_2416_));
 sky130_fd_sc_hd__mux2_1 _5580_ (.A0(\z80.tv80s.di_reg[5] ),
    .A1(_2416_),
    .S(_2367_),
    .X(_2417_));
 sky130_fd_sc_hd__mux2_1 _5581_ (.A0(net782),
    .A1(_2417_),
    .S(net117),
    .X(_0278_));
 sky130_fd_sc_hd__mux2_1 _5582_ (.A0(\z80.tv80s.i_tv80_core.SP[14] ),
    .A1(_1960_),
    .S(net121),
    .X(_2418_));
 sky130_fd_sc_hd__and2_1 _5583_ (.A(net72),
    .B(_2418_),
    .X(_2419_));
 sky130_fd_sc_hd__nor2_1 _5584_ (.A(net72),
    .B(_2418_),
    .Y(_2420_));
 sky130_fd_sc_hd__nor2_1 _5585_ (.A(_2419_),
    .B(_2420_),
    .Y(_2421_));
 sky130_fd_sc_hd__o21ai_1 _5586_ (.A1(_2411_),
    .A2(_2412_),
    .B1(_2409_),
    .Y(_2422_));
 sky130_fd_sc_hd__xor2_1 _5587_ (.A(_2421_),
    .B(_2422_),
    .X(_2423_));
 sky130_fd_sc_hd__a22o_1 _5588_ (.A1(net751),
    .A2(_2273_),
    .B1(_2423_),
    .B2(_2265_),
    .X(_2424_));
 sky130_fd_sc_hd__mux2_1 _5589_ (.A0(net751),
    .A1(_2424_),
    .S(net93),
    .X(_2425_));
 sky130_fd_sc_hd__mux2_1 _5590_ (.A0(\z80.tv80s.di_reg[6] ),
    .A1(_2425_),
    .S(_2367_),
    .X(_2426_));
 sky130_fd_sc_hd__mux2_1 _5591_ (.A0(net751),
    .A1(_2426_),
    .S(net112),
    .X(_0279_));
 sky130_fd_sc_hd__a21oi_1 _5592_ (.A1(_2421_),
    .A2(_2422_),
    .B1(_2419_),
    .Y(_2427_));
 sky130_fd_sc_hd__mux2_1 _5593_ (.A0(\z80.tv80s.i_tv80_core.SP[15] ),
    .A1(_1980_),
    .S(net121),
    .X(_2428_));
 sky130_fd_sc_hd__xor2_1 _5594_ (.A(net72),
    .B(_2428_),
    .X(_2429_));
 sky130_fd_sc_hd__xnor2_1 _5595_ (.A(_2427_),
    .B(_2429_),
    .Y(_2430_));
 sky130_fd_sc_hd__a22o_1 _5596_ (.A1(net759),
    .A2(_2273_),
    .B1(_2430_),
    .B2(_2265_),
    .X(_2431_));
 sky130_fd_sc_hd__mux2_1 _5597_ (.A0(net759),
    .A1(_2431_),
    .S(net93),
    .X(_2432_));
 sky130_fd_sc_hd__mux2_1 _5598_ (.A0(\z80.tv80s.di_reg[7] ),
    .A1(_2432_),
    .S(_2367_),
    .X(_2433_));
 sky130_fd_sc_hd__mux2_1 _5599_ (.A0(net759),
    .A1(_2433_),
    .S(net112),
    .X(_0280_));
 sky130_fd_sc_hd__and3_1 _5600_ (.A(net166),
    .B(_2946_),
    .C(_0602_),
    .X(_2434_));
 sky130_fd_sc_hd__xor2_1 _5601_ (.A(net473),
    .B(_2434_),
    .X(_0281_));
 sky130_fd_sc_hd__a221o_1 _5602_ (.A1(_2948_),
    .A2(_0401_),
    .B1(_0684_),
    .B2(net96),
    .C1(_1393_),
    .X(_2435_));
 sky130_fd_sc_hd__or4_1 _5603_ (.A(_0746_),
    .B(_0748_),
    .C(_0749_),
    .D(_2435_),
    .X(_2436_));
 sky130_fd_sc_hd__a31o_1 _5604_ (.A1(net96),
    .A2(_0422_),
    .A3(_0461_),
    .B1(_2436_),
    .X(_2437_));
 sky130_fd_sc_hd__and4_1 _5605_ (.A(net120),
    .B(net147),
    .C(net146),
    .D(_1384_),
    .X(_2438_));
 sky130_fd_sc_hd__a221o_1 _5606_ (.A1(net134),
    .A2(_3041_),
    .B1(_1385_),
    .B2(net96),
    .C1(_2438_),
    .X(_2439_));
 sky130_fd_sc_hd__a22o_1 _5607_ (.A1(net164),
    .A2(_2437_),
    .B1(_2439_),
    .B2(net106),
    .X(_2440_));
 sky130_fd_sc_hd__and2_2 _5608_ (.A(_2842_),
    .B(_2440_),
    .X(_2441_));
 sky130_fd_sc_hd__inv_2 _5609_ (.A(_2441_),
    .Y(_2442_));
 sky130_fd_sc_hd__and2_1 _5610_ (.A(_1412_),
    .B(_2441_),
    .X(_2443_));
 sky130_fd_sc_hd__a21oi_4 _5611_ (.A1(_1401_),
    .A2(_2443_),
    .B1(net128),
    .Y(_2444_));
 sky130_fd_sc_hd__nor2_1 _5612_ (.A(_1412_),
    .B(_2442_),
    .Y(_2445_));
 sky130_fd_sc_hd__a31o_1 _5613_ (.A1(net166),
    .A2(net109),
    .A3(_1397_),
    .B1(_1383_),
    .X(_2446_));
 sky130_fd_sc_hd__a21oi_1 _5614_ (.A1(\z80.tv80s.i_tv80_core.i_mcode.MCycle[3] ),
    .A2(net96),
    .B1(net130),
    .Y(_2447_));
 sky130_fd_sc_hd__a221oi_1 _5615_ (.A1(net152),
    .A2(_1384_),
    .B1(_1512_),
    .B2(_2991_),
    .C1(_2999_),
    .Y(_2448_));
 sky130_fd_sc_hd__o31a_1 _5616_ (.A1(_0666_),
    .A2(_1510_),
    .A3(_2447_),
    .B1(_2448_),
    .X(_2449_));
 sky130_fd_sc_hd__nor2_1 _5617_ (.A(_0437_),
    .B(_0481_),
    .Y(_2450_));
 sky130_fd_sc_hd__a211o_1 _5618_ (.A1(_3026_),
    .A2(_0405_),
    .B1(_1403_),
    .C1(_2450_),
    .X(_2451_));
 sky130_fd_sc_hd__nor2_1 _5619_ (.A(_0525_),
    .B(_1511_),
    .Y(_2452_));
 sky130_fd_sc_hd__a221o_1 _5620_ (.A1(net160),
    .A2(_2971_),
    .B1(_0461_),
    .B2(_2944_),
    .C1(_2452_),
    .X(_2453_));
 sky130_fd_sc_hd__o211a_1 _5621_ (.A1(_2849_),
    .A2(net96),
    .B1(_0401_),
    .C1(_0422_),
    .X(_2454_));
 sky130_fd_sc_hd__a211o_1 _5622_ (.A1(_2909_),
    .A2(_0484_),
    .B1(_1390_),
    .C1(_2948_),
    .X(_2455_));
 sky130_fd_sc_hd__a22o_1 _5623_ (.A1(_0512_),
    .A2(_2451_),
    .B1(_2455_),
    .B2(net134),
    .X(_2456_));
 sky130_fd_sc_hd__or4_1 _5624_ (.A(_1394_),
    .B(_2453_),
    .C(_2454_),
    .D(_2456_),
    .X(_2457_));
 sky130_fd_sc_hd__o2bb2a_1 _5625_ (.A1_N(net164),
    .A2_N(_2457_),
    .B1(net105),
    .B2(_2449_),
    .X(_2458_));
 sky130_fd_sc_hd__o2bb2a_4 _5626_ (.A1_N(net161),
    .A2_N(_2446_),
    .B1(_2458_),
    .B2(\z80.tv80s.i_tv80_core.i_mcode.MCycle[6] ),
    .X(_2459_));
 sky130_fd_sc_hd__inv_2 _5627_ (.A(_2459_),
    .Y(_2460_));
 sky130_fd_sc_hd__and3_2 _5628_ (.A(_1401_),
    .B(_2445_),
    .C(_2460_),
    .X(_2461_));
 sky130_fd_sc_hd__and3b_2 _5629_ (.A_N(_1401_),
    .B(_2445_),
    .C(_2459_),
    .X(_2462_));
 sky130_fd_sc_hd__and4_2 _5630_ (.A(_1401_),
    .B(_1412_),
    .C(_2442_),
    .D(_2460_),
    .X(_2463_));
 sky130_fd_sc_hd__a21o_1 _5631_ (.A1(_1401_),
    .A2(_1412_),
    .B1(_2441_),
    .X(_2464_));
 sky130_fd_sc_hd__inv_2 _5632_ (.A(_2464_),
    .Y(_2465_));
 sky130_fd_sc_hd__a221o_1 _5633_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][0] ),
    .A2(net142),
    .B1(net84),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][0] ),
    .C1(net75),
    .X(_2466_));
 sky130_fd_sc_hd__a221o_1 _5634_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][0] ),
    .A2(net142),
    .B1(net84),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][0] ),
    .C1(_0984_),
    .X(_2467_));
 sky130_fd_sc_hd__a221o_1 _5635_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][0] ),
    .A2(net141),
    .B1(net83),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][0] ),
    .C1(net75),
    .X(_2468_));
 sky130_fd_sc_hd__a221o_1 _5636_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][0] ),
    .A2(net141),
    .B1(net83),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][0] ),
    .C1(net73),
    .X(_2469_));
 sky130_fd_sc_hd__and2_1 _5637_ (.A(_1300_),
    .B(_1434_),
    .X(_2470_));
 sky130_fd_sc_hd__a31o_1 _5638_ (.A1(_1299_),
    .A2(_2466_),
    .A3(_2467_),
    .B1(_2470_),
    .X(_2471_));
 sky130_fd_sc_hd__and3_1 _5639_ (.A(_1299_),
    .B(_2468_),
    .C(_2469_),
    .X(_2472_));
 sky130_fd_sc_hd__a211o_1 _5640_ (.A1(_0985_),
    .A2(_1300_),
    .B1(_2460_),
    .C1(_2472_),
    .X(_2473_));
 sky130_fd_sc_hd__o211a_1 _5641_ (.A1(_2459_),
    .A2(_2471_),
    .B1(_2473_),
    .C1(_2465_),
    .X(_2474_));
 sky130_fd_sc_hd__nor2_1 _5642_ (.A(_1401_),
    .B(_2459_),
    .Y(_2475_));
 sky130_fd_sc_hd__and2_2 _5643_ (.A(_2443_),
    .B(_2475_),
    .X(_2476_));
 sky130_fd_sc_hd__and2_1 _5644_ (.A(_1401_),
    .B(_2459_),
    .X(_2477_));
 sky130_fd_sc_hd__and3_2 _5645_ (.A(_1412_),
    .B(_2442_),
    .C(_2477_),
    .X(_2478_));
 sky130_fd_sc_hd__and3b_2 _5646_ (.A_N(_1401_),
    .B(_2443_),
    .C(_2459_),
    .X(_2479_));
 sky130_fd_sc_hd__a21o_1 _5647_ (.A1(\z80.tv80s.i_tv80_core.SP[8] ),
    .A2(_2475_),
    .B1(_2477_),
    .X(_2480_));
 sky130_fd_sc_hd__a22o_1 _5648_ (.A1(\z80.tv80s.i_tv80_core.F[0] ),
    .A2(_2461_),
    .B1(_2463_),
    .B2(\z80.tv80s.i_tv80_core.ACC[0] ),
    .X(_2481_));
 sky130_fd_sc_hd__a211o_1 _5649_ (.A1(net637),
    .A2(_2462_),
    .B1(_2474_),
    .C1(_2481_),
    .X(_2482_));
 sky130_fd_sc_hd__a221o_1 _5650_ (.A1(\z80.tv80s.di_reg[0] ),
    .A2(_2478_),
    .B1(_2480_),
    .B2(_2445_),
    .C1(_2482_),
    .X(_2483_));
 sky130_fd_sc_hd__a221o_1 _5651_ (.A1(\z80.tv80s.i_tv80_core.PC[8] ),
    .A2(_2476_),
    .B1(_2479_),
    .B2(net641),
    .C1(_2483_),
    .X(_2484_));
 sky130_fd_sc_hd__a22o_1 _5652_ (.A1(net125),
    .A2(net709),
    .B1(_2444_),
    .B2(_2484_),
    .X(_0282_));
 sky130_fd_sc_hd__and2_2 _5653_ (.A(_2445_),
    .B(_2475_),
    .X(_2485_));
 sky130_fd_sc_hd__a22o_1 _5654_ (.A1(\z80.tv80s.i_tv80_core.PC[9] ),
    .A2(_2476_),
    .B1(_2478_),
    .B2(\z80.tv80s.di_reg[1] ),
    .X(_2486_));
 sky130_fd_sc_hd__or2_1 _5655_ (.A(_1027_),
    .B(_1299_),
    .X(_2487_));
 sky130_fd_sc_hd__o221a_1 _5656_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][1] ),
    .A2(net142),
    .B1(net83),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][1] ),
    .C1(net73),
    .X(_2488_));
 sky130_fd_sc_hd__o221a_1 _5657_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][1] ),
    .A2(net142),
    .B1(net83),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][1] ),
    .C1(net75),
    .X(_2489_));
 sky130_fd_sc_hd__o31a_1 _5658_ (.A1(_1300_),
    .A2(_2488_),
    .A3(_2489_),
    .B1(_2487_),
    .X(_2490_));
 sky130_fd_sc_hd__mux2_1 _5659_ (.A0(_1442_),
    .A1(_2490_),
    .S(_2459_),
    .X(_2491_));
 sky130_fd_sc_hd__a221o_1 _5660_ (.A1(\z80.tv80s.i_tv80_core.F[1] ),
    .A2(_2461_),
    .B1(_2485_),
    .B2(\z80.tv80s.i_tv80_core.SP[9] ),
    .C1(_2486_),
    .X(_2492_));
 sky130_fd_sc_hd__a22o_1 _5661_ (.A1(\z80.tv80s.i_tv80_core.SP[1] ),
    .A2(_2462_),
    .B1(_2465_),
    .B2(_2491_),
    .X(_2493_));
 sky130_fd_sc_hd__a22o_1 _5662_ (.A1(\z80.tv80s.i_tv80_core.ACC[1] ),
    .A2(_2463_),
    .B1(_2479_),
    .B2(\z80.tv80s.i_tv80_core.PC[1] ),
    .X(_2494_));
 sky130_fd_sc_hd__or3_1 _5663_ (.A(_2492_),
    .B(_2493_),
    .C(_2494_),
    .X(_2495_));
 sky130_fd_sc_hd__a22o_1 _5664_ (.A1(net125),
    .A2(net645),
    .B1(_2444_),
    .B2(_2495_),
    .X(_0283_));
 sky130_fd_sc_hd__a22o_1 _5665_ (.A1(\z80.tv80s.di_reg[2] ),
    .A2(_2478_),
    .B1(_2479_),
    .B2(net617),
    .X(_2496_));
 sky130_fd_sc_hd__a22o_1 _5666_ (.A1(\z80.tv80s.i_tv80_core.F[2] ),
    .A2(_2461_),
    .B1(_2476_),
    .B2(\z80.tv80s.i_tv80_core.PC[10] ),
    .X(_2497_));
 sky130_fd_sc_hd__o221a_1 _5667_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][2] ),
    .A2(net141),
    .B1(net83),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][2] ),
    .C1(net73),
    .X(_2498_));
 sky130_fd_sc_hd__o221a_1 _5668_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][2] ),
    .A2(net141),
    .B1(net83),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][2] ),
    .C1(net75),
    .X(_2499_));
 sky130_fd_sc_hd__or2_1 _5669_ (.A(_1300_),
    .B(_2499_),
    .X(_2500_));
 sky130_fd_sc_hd__o22a_1 _5670_ (.A1(_1029_),
    .A2(_1299_),
    .B1(_2498_),
    .B2(_2500_),
    .X(_2501_));
 sky130_fd_sc_hd__mux2_1 _5671_ (.A0(_1453_),
    .A1(_2501_),
    .S(_2459_),
    .X(_2502_));
 sky130_fd_sc_hd__a22o_1 _5672_ (.A1(\z80.tv80s.i_tv80_core.ACC[2] ),
    .A2(_2463_),
    .B1(_2465_),
    .B2(_2502_),
    .X(_2503_));
 sky130_fd_sc_hd__a221o_1 _5673_ (.A1(net713),
    .A2(_2462_),
    .B1(_2485_),
    .B2(net583),
    .C1(_2503_),
    .X(_2504_));
 sky130_fd_sc_hd__or3_1 _5674_ (.A(_2496_),
    .B(_2497_),
    .C(_2504_),
    .X(_2505_));
 sky130_fd_sc_hd__a22o_1 _5675_ (.A1(net125),
    .A2(net774),
    .B1(_2444_),
    .B2(_2505_),
    .X(_0284_));
 sky130_fd_sc_hd__a22o_1 _5676_ (.A1(\z80.tv80s.i_tv80_core.SP[3] ),
    .A2(_2462_),
    .B1(_2479_),
    .B2(net595),
    .X(_2506_));
 sky130_fd_sc_hd__a22o_1 _5677_ (.A1(\z80.tv80s.i_tv80_core.F[3] ),
    .A2(_2461_),
    .B1(_2476_),
    .B2(\z80.tv80s.i_tv80_core.PC[11] ),
    .X(_2507_));
 sky130_fd_sc_hd__o221a_1 _5678_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][3] ),
    .A2(net142),
    .B1(net84),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][3] ),
    .C1(_0984_),
    .X(_2508_));
 sky130_fd_sc_hd__o221a_1 _5679_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][3] ),
    .A2(net142),
    .B1(net84),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][3] ),
    .C1(net75),
    .X(_2509_));
 sky130_fd_sc_hd__or2_1 _5680_ (.A(_2508_),
    .B(_2509_),
    .X(_2510_));
 sky130_fd_sc_hd__o221a_1 _5681_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][3] ),
    .A2(net141),
    .B1(net82),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][3] ),
    .C1(net73),
    .X(_2511_));
 sky130_fd_sc_hd__o221a_1 _5682_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][3] ),
    .A2(net141),
    .B1(net82),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][3] ),
    .C1(net74),
    .X(_2512_));
 sky130_fd_sc_hd__or2_1 _5683_ (.A(_2511_),
    .B(_2512_),
    .X(_2513_));
 sky130_fd_sc_hd__mux4_2 _5684_ (.A0(_1462_),
    .A1(_2510_),
    .A2(_1113_),
    .A3(_2513_),
    .S0(_1299_),
    .S1(_2459_),
    .X(_2514_));
 sky130_fd_sc_hd__a22o_1 _5685_ (.A1(\z80.tv80s.di_reg[3] ),
    .A2(_2478_),
    .B1(_2514_),
    .B2(_2465_),
    .X(_2515_));
 sky130_fd_sc_hd__a221o_1 _5686_ (.A1(\z80.tv80s.i_tv80_core.ACC[3] ),
    .A2(_2463_),
    .B1(_2485_),
    .B2(\z80.tv80s.i_tv80_core.SP[11] ),
    .C1(_2515_),
    .X(_2516_));
 sky130_fd_sc_hd__or3_1 _5687_ (.A(_2506_),
    .B(_2507_),
    .C(_2516_),
    .X(_2517_));
 sky130_fd_sc_hd__a22o_1 _5688_ (.A1(net125),
    .A2(net649),
    .B1(_2444_),
    .B2(_2517_),
    .X(_0285_));
 sky130_fd_sc_hd__a22o_1 _5689_ (.A1(net662),
    .A2(_2462_),
    .B1(_2479_),
    .B2(net599),
    .X(_2518_));
 sky130_fd_sc_hd__a22o_1 _5690_ (.A1(\z80.tv80s.i_tv80_core.F[4] ),
    .A2(_2461_),
    .B1(_2476_),
    .B2(\z80.tv80s.i_tv80_core.PC[12] ),
    .X(_2519_));
 sky130_fd_sc_hd__o221a_1 _5691_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][4] ),
    .A2(net141),
    .B1(net82),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][4] ),
    .C1(net73),
    .X(_2520_));
 sky130_fd_sc_hd__o221a_1 _5692_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][4] ),
    .A2(net141),
    .B1(net82),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][4] ),
    .C1(net74),
    .X(_2521_));
 sky130_fd_sc_hd__or2_1 _5693_ (.A(_2520_),
    .B(_2521_),
    .X(_2522_));
 sky130_fd_sc_hd__o221a_1 _5694_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][4] ),
    .A2(net141),
    .B1(net83),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][4] ),
    .C1(net73),
    .X(_2523_));
 sky130_fd_sc_hd__o221a_1 _5695_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][4] ),
    .A2(net141),
    .B1(net83),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][4] ),
    .C1(net74),
    .X(_2524_));
 sky130_fd_sc_hd__or2_1 _5696_ (.A(_2523_),
    .B(_2524_),
    .X(_2525_));
 sky130_fd_sc_hd__mux4_2 _5697_ (.A0(_1467_),
    .A1(_2522_),
    .A2(_1155_),
    .A3(_2525_),
    .S0(_1299_),
    .S1(_2459_),
    .X(_2526_));
 sky130_fd_sc_hd__a22o_1 _5698_ (.A1(\z80.tv80s.di_reg[4] ),
    .A2(_2478_),
    .B1(_2526_),
    .B2(_2465_),
    .X(_2527_));
 sky130_fd_sc_hd__a221o_1 _5699_ (.A1(\z80.tv80s.i_tv80_core.ACC[4] ),
    .A2(_2463_),
    .B1(_2485_),
    .B2(\z80.tv80s.i_tv80_core.SP[12] ),
    .C1(_2527_),
    .X(_2528_));
 sky130_fd_sc_hd__or3_1 _5700_ (.A(_2518_),
    .B(_2519_),
    .C(_2528_),
    .X(_2529_));
 sky130_fd_sc_hd__a22o_1 _5701_ (.A1(net128),
    .A2(net728),
    .B1(_2444_),
    .B2(_2529_),
    .X(_0286_));
 sky130_fd_sc_hd__a22o_1 _5702_ (.A1(\z80.tv80s.i_tv80_core.SP[5] ),
    .A2(_2462_),
    .B1(_2479_),
    .B2(net577),
    .X(_2530_));
 sky130_fd_sc_hd__a22o_1 _5703_ (.A1(\z80.tv80s.i_tv80_core.F[5] ),
    .A2(_2461_),
    .B1(_2476_),
    .B2(\z80.tv80s.i_tv80_core.PC[13] ),
    .X(_2531_));
 sky130_fd_sc_hd__o221a_1 _5704_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][5] ),
    .A2(net141),
    .B1(net82),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][5] ),
    .C1(net73),
    .X(_2532_));
 sky130_fd_sc_hd__o221a_1 _5705_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][5] ),
    .A2(net141),
    .B1(net82),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][5] ),
    .C1(net74),
    .X(_2533_));
 sky130_fd_sc_hd__or2_1 _5706_ (.A(_2532_),
    .B(_2533_),
    .X(_2534_));
 sky130_fd_sc_hd__o221a_1 _5707_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][5] ),
    .A2(net141),
    .B1(net82),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][5] ),
    .C1(net73),
    .X(_2535_));
 sky130_fd_sc_hd__o221a_1 _5708_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][5] ),
    .A2(net141),
    .B1(net82),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][5] ),
    .C1(net74),
    .X(_2536_));
 sky130_fd_sc_hd__or2_1 _5709_ (.A(_2535_),
    .B(_2536_),
    .X(_2537_));
 sky130_fd_sc_hd__mux4_2 _5710_ (.A0(_1473_),
    .A1(_2534_),
    .A2(_1207_),
    .A3(_2537_),
    .S0(_1299_),
    .S1(_2459_),
    .X(_2538_));
 sky130_fd_sc_hd__a22o_1 _5711_ (.A1(\z80.tv80s.di_reg[5] ),
    .A2(_2478_),
    .B1(_2538_),
    .B2(_2465_),
    .X(_2539_));
 sky130_fd_sc_hd__a221o_1 _5712_ (.A1(\z80.tv80s.i_tv80_core.ACC[5] ),
    .A2(_2463_),
    .B1(_2485_),
    .B2(\z80.tv80s.i_tv80_core.SP[13] ),
    .C1(_2539_),
    .X(_2540_));
 sky130_fd_sc_hd__or3_1 _5713_ (.A(_2530_),
    .B(_2531_),
    .C(_2540_),
    .X(_2541_));
 sky130_fd_sc_hd__a22o_1 _5714_ (.A1(net128),
    .A2(net643),
    .B1(_2444_),
    .B2(_2541_),
    .X(_0287_));
 sky130_fd_sc_hd__a22o_1 _5715_ (.A1(\z80.tv80s.i_tv80_core.SP[6] ),
    .A2(_2462_),
    .B1(_2479_),
    .B2(\z80.tv80s.i_tv80_core.PC[6] ),
    .X(_2542_));
 sky130_fd_sc_hd__a22o_1 _5716_ (.A1(\z80.tv80s.i_tv80_core.F[6] ),
    .A2(_2461_),
    .B1(_2476_),
    .B2(\z80.tv80s.i_tv80_core.PC[14] ),
    .X(_2543_));
 sky130_fd_sc_hd__o221a_1 _5717_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][6] ),
    .A2(\z80.tv80s.i_tv80_core.RegAddrB_r[0] ),
    .B1(net84),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][6] ),
    .C1(_0984_),
    .X(_2544_));
 sky130_fd_sc_hd__o221a_1 _5718_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][6] ),
    .A2(\z80.tv80s.i_tv80_core.RegAddrB_r[0] ),
    .B1(net84),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][6] ),
    .C1(_0983_),
    .X(_2545_));
 sky130_fd_sc_hd__or2_1 _5719_ (.A(_2544_),
    .B(_2545_),
    .X(_2546_));
 sky130_fd_sc_hd__o221a_1 _5720_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][6] ),
    .A2(net141),
    .B1(net82),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][6] ),
    .C1(net73),
    .X(_2547_));
 sky130_fd_sc_hd__o221a_1 _5721_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][6] ),
    .A2(net141),
    .B1(net82),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][6] ),
    .C1(net74),
    .X(_2548_));
 sky130_fd_sc_hd__or2_1 _5722_ (.A(_2547_),
    .B(_2548_),
    .X(_2549_));
 sky130_fd_sc_hd__mux4_2 _5723_ (.A0(_1480_),
    .A1(_2546_),
    .A2(_1250_),
    .A3(_2549_),
    .S0(_1299_),
    .S1(_2459_),
    .X(_2550_));
 sky130_fd_sc_hd__a22o_1 _5724_ (.A1(\z80.tv80s.di_reg[6] ),
    .A2(_2478_),
    .B1(_2550_),
    .B2(_2465_),
    .X(_2551_));
 sky130_fd_sc_hd__a221o_1 _5725_ (.A1(\z80.tv80s.i_tv80_core.ACC[6] ),
    .A2(_2463_),
    .B1(_2485_),
    .B2(\z80.tv80s.i_tv80_core.SP[14] ),
    .C1(_2551_),
    .X(_2552_));
 sky130_fd_sc_hd__or3_1 _5726_ (.A(_2542_),
    .B(_2543_),
    .C(_2552_),
    .X(_2553_));
 sky130_fd_sc_hd__a22o_1 _5727_ (.A1(net128),
    .A2(net619),
    .B1(_2444_),
    .B2(_2553_),
    .X(_0288_));
 sky130_fd_sc_hd__a22o_1 _5728_ (.A1(\z80.tv80s.i_tv80_core.F[7] ),
    .A2(_2461_),
    .B1(_2462_),
    .B2(\z80.tv80s.i_tv80_core.SP[7] ),
    .X(_2554_));
 sky130_fd_sc_hd__a22o_1 _5729_ (.A1(\z80.tv80s.i_tv80_core.ACC[7] ),
    .A2(_2463_),
    .B1(_2485_),
    .B2(\z80.tv80s.i_tv80_core.SP[15] ),
    .X(_2555_));
 sky130_fd_sc_hd__o221a_1 _5730_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][7] ),
    .A2(net142),
    .B1(net84),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][7] ),
    .C1(net73),
    .X(_2556_));
 sky130_fd_sc_hd__o221a_1 _5731_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][7] ),
    .A2(net142),
    .B1(net84),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][7] ),
    .C1(net75),
    .X(_2557_));
 sky130_fd_sc_hd__or2_1 _5732_ (.A(_1300_),
    .B(_2557_),
    .X(_2558_));
 sky130_fd_sc_hd__o22a_1 _5733_ (.A1(_1299_),
    .A2(_1482_),
    .B1(_2556_),
    .B2(_2558_),
    .X(_2559_));
 sky130_fd_sc_hd__mux2_1 _5734_ (.A0(_2559_),
    .A1(_1307_),
    .S(_2459_),
    .X(_2560_));
 sky130_fd_sc_hd__a22o_1 _5735_ (.A1(\z80.tv80s.i_tv80_core.PC[7] ),
    .A2(_2479_),
    .B1(_2560_),
    .B2(_2465_),
    .X(_2561_));
 sky130_fd_sc_hd__a221o_1 _5736_ (.A1(\z80.tv80s.i_tv80_core.PC[15] ),
    .A2(_2476_),
    .B1(_2478_),
    .B2(\z80.tv80s.di_reg[7] ),
    .C1(_2561_),
    .X(_2562_));
 sky130_fd_sc_hd__or3_1 _5737_ (.A(_2554_),
    .B(_2555_),
    .C(_2562_),
    .X(_2563_));
 sky130_fd_sc_hd__a22o_1 _5738_ (.A1(net125),
    .A2(net639),
    .B1(_2444_),
    .B2(_2563_),
    .X(_0289_));
 sky130_fd_sc_hd__mux2_1 _5739_ (.A0(_2882_),
    .A1(_0964_),
    .S(net113),
    .X(_2564_));
 sky130_fd_sc_hd__inv_2 _5740_ (.A(_2564_),
    .Y(_0290_));
 sky130_fd_sc_hd__mux2_1 _5741_ (.A0(_2883_),
    .A1(_0952_),
    .S(net113),
    .X(_2565_));
 sky130_fd_sc_hd__inv_2 _5742_ (.A(_2565_),
    .Y(_0291_));
 sky130_fd_sc_hd__mux2_1 _5743_ (.A0(net249),
    .A1(_0942_),
    .S(net113),
    .X(_0292_));
 sky130_fd_sc_hd__mux2_1 _5744_ (.A0(net253),
    .A1(_0931_),
    .S(net113),
    .X(_0293_));
 sky130_fd_sc_hd__mux2_1 _5745_ (.A0(net223),
    .A1(_0921_),
    .S(net112),
    .X(_0294_));
 sky130_fd_sc_hd__mux2_1 _5746_ (.A0(net247),
    .A1(_0913_),
    .S(net112),
    .X(_0295_));
 sky130_fd_sc_hd__mux2_1 _5747_ (.A0(net251),
    .A1(_0905_),
    .S(net112),
    .X(_0296_));
 sky130_fd_sc_hd__mux2_1 _5748_ (.A0(net233),
    .A1(_0897_),
    .S(net112),
    .X(_0297_));
 sky130_fd_sc_hd__mux2_1 _5749_ (.A0(net229),
    .A1(_0889_),
    .S(net112),
    .X(_0298_));
 sky130_fd_sc_hd__mux2_1 _5750_ (.A0(net243),
    .A1(_1021_),
    .S(net112),
    .X(_0299_));
 sky130_fd_sc_hd__mux2_1 _5751_ (.A0(net237),
    .A1(_1034_),
    .S(net112),
    .X(_0300_));
 sky130_fd_sc_hd__mux2_1 _5752_ (.A0(net235),
    .A1(_1107_),
    .S(net112),
    .X(_0301_));
 sky130_fd_sc_hd__mux2_1 _5753_ (.A0(net245),
    .A1(_1122_),
    .S(net112),
    .X(_0302_));
 sky130_fd_sc_hd__mux2_1 _5754_ (.A0(net241),
    .A1(_1198_),
    .S(net112),
    .X(_0303_));
 sky130_fd_sc_hd__mux2_1 _5755_ (.A0(net227),
    .A1(_1213_),
    .S(net112),
    .X(_0304_));
 sky130_fd_sc_hd__mux2_1 _5756_ (.A0(net231),
    .A1(_1257_),
    .S(net112),
    .X(_0305_));
 sky130_fd_sc_hd__or4b_4 _5757_ (.A(_2854_),
    .B(net125),
    .C(_0477_),
    .D_N(_1354_),
    .X(_2566_));
 sky130_fd_sc_hd__mux2_1 _5758_ (.A0(\z80.tv80s.i_tv80_core.ACC[0] ),
    .A1(net581),
    .S(_2566_),
    .X(_0306_));
 sky130_fd_sc_hd__mux2_1 _5759_ (.A0(\z80.tv80s.i_tv80_core.ACC[1] ),
    .A1(net676),
    .S(_2566_),
    .X(_0307_));
 sky130_fd_sc_hd__mux2_1 _5760_ (.A0(\z80.tv80s.i_tv80_core.ACC[2] ),
    .A1(net623),
    .S(_2566_),
    .X(_0308_));
 sky130_fd_sc_hd__mux2_1 _5761_ (.A0(\z80.tv80s.i_tv80_core.ACC[3] ),
    .A1(net627),
    .S(_2566_),
    .X(_0309_));
 sky130_fd_sc_hd__mux2_1 _5762_ (.A0(\z80.tv80s.i_tv80_core.ACC[4] ),
    .A1(net579),
    .S(_2566_),
    .X(_0310_));
 sky130_fd_sc_hd__mux2_1 _5763_ (.A0(\z80.tv80s.i_tv80_core.ACC[5] ),
    .A1(net722),
    .S(_2566_),
    .X(_0311_));
 sky130_fd_sc_hd__mux2_1 _5764_ (.A0(\z80.tv80s.i_tv80_core.ACC[6] ),
    .A1(net732),
    .S(_2566_),
    .X(_0312_));
 sky130_fd_sc_hd__mux2_1 _5765_ (.A0(\z80.tv80s.i_tv80_core.ACC[7] ),
    .A1(net792),
    .S(_2566_),
    .X(_0313_));
 sky130_fd_sc_hd__mux2_1 _5766_ (.A0(\z80.tv80s.i_tv80_core.ACC[7] ),
    .A1(net494),
    .S(_1382_),
    .X(_0314_));
 sky130_fd_sc_hd__nand2_1 _5767_ (.A(_1333_),
    .B(_1351_),
    .Y(_2567_));
 sky130_fd_sc_hd__mux2_1 _5768_ (.A0(net261),
    .A1(_2567_),
    .S(net113),
    .X(_0315_));
 sky130_fd_sc_hd__mux2_1 _5769_ (.A0(net239),
    .A1(_1350_),
    .S(net113),
    .X(_0316_));
 sky130_fd_sc_hd__or4b_2 _5770_ (.A(\z80.tv80s.i_tv80_core.Halt_FF ),
    .B(_0484_),
    .C(_0735_),
    .D_N(_1680_),
    .X(_2568_));
 sky130_fd_sc_hd__nor2_1 _5771_ (.A(net78),
    .B(_2568_),
    .Y(_2569_));
 sky130_fd_sc_hd__o21a_2 _5772_ (.A1(net94),
    .A2(_2569_),
    .B1(_0605_),
    .X(_2570_));
 sky130_fd_sc_hd__a2111o_1 _5773_ (.A1(_2896_),
    .A2(_2982_),
    .B1(_0418_),
    .C1(_0429_),
    .D1(_2912_),
    .X(_2571_));
 sky130_fd_sc_hd__or4b_1 _5774_ (.A(_2965_),
    .B(_0416_),
    .C(_0439_),
    .D_N(_0442_),
    .X(_2572_));
 sky130_fd_sc_hd__a21oi_1 _5775_ (.A1(\z80.tv80s.i_tv80_core.i_mcode.MCycle[1] ),
    .A2(_2571_),
    .B1(_2572_),
    .Y(_2573_));
 sky130_fd_sc_hd__o32a_1 _5776_ (.A1(_2908_),
    .A2(_3020_),
    .A3(_0462_),
    .B1(_2573_),
    .B2(_0397_),
    .X(_2574_));
 sky130_fd_sc_hd__or3b_1 _5777_ (.A(net134),
    .B(_0554_),
    .C_N(_0623_),
    .X(_2575_));
 sky130_fd_sc_hd__a21oi_1 _5778_ (.A1(_2574_),
    .A2(_2575_),
    .B1(net118),
    .Y(_2576_));
 sky130_fd_sc_hd__o21bai_4 _5779_ (.A1(net119),
    .A2(_0685_),
    .B1_N(\z80.tv80s.i_tv80_core.BTR_r ),
    .Y(_2577_));
 sky130_fd_sc_hd__o21a_1 _5780_ (.A1(net163),
    .A2(_2893_),
    .B1(net129),
    .X(_2578_));
 sky130_fd_sc_hd__a311o_1 _5781_ (.A1(net107),
    .A2(_0390_),
    .A3(_0398_),
    .B1(_2578_),
    .C1(\z80.tv80s.i_tv80_core.i_mcode.MCycle[5] ),
    .X(_2579_));
 sky130_fd_sc_hd__o31a_1 _5782_ (.A1(_2576_),
    .A2(_2577_),
    .A3(_2579_),
    .B1(_0603_),
    .X(_2580_));
 sky130_fd_sc_hd__or2_2 _5783_ (.A(net102),
    .B(_2580_),
    .X(_2581_));
 sky130_fd_sc_hd__o21a_2 _5784_ (.A1(_0577_),
    .A2(net64),
    .B1(net63),
    .X(_2582_));
 sky130_fd_sc_hd__o21ai_4 _5785_ (.A1(_0577_),
    .A2(net64),
    .B1(net63),
    .Y(_2583_));
 sky130_fd_sc_hd__nor2_4 _5786_ (.A(_2008_),
    .B(_2580_),
    .Y(_2584_));
 sky130_fd_sc_hd__mux2_1 _5787_ (.A0(\z80.tv80s.i_tv80_core.TmpAddr[0] ),
    .A1(\z80.tv80s.i_tv80_core.PC[0] ),
    .S(net99),
    .X(_2585_));
 sky130_fd_sc_hd__a221o_1 _5788_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[0] ),
    .A2(net68),
    .B1(net66),
    .B2(_2585_),
    .C1(net90),
    .X(_2586_));
 sky130_fd_sc_hd__a22oi_1 _5789_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[0] ),
    .A2(net78),
    .B1(_1674_),
    .B2(_2586_),
    .Y(_2587_));
 sky130_fd_sc_hd__o31ai_1 _5790_ (.A1(net119),
    .A2(_2872_),
    .A3(_0685_),
    .B1(_2577_),
    .Y(_2588_));
 sky130_fd_sc_hd__nand2_1 _5791_ (.A(net641),
    .B(_2588_),
    .Y(_2589_));
 sky130_fd_sc_hd__or2_1 _5792_ (.A(net641),
    .B(_2588_),
    .X(_2590_));
 sky130_fd_sc_hd__nand2_1 _5793_ (.A(_2589_),
    .B(_2590_),
    .Y(_2591_));
 sky130_fd_sc_hd__a22o_1 _5794_ (.A1(_2584_),
    .A2(_2587_),
    .B1(_2591_),
    .B2(net64),
    .X(_2592_));
 sky130_fd_sc_hd__o2bb2a_1 _5795_ (.A1_N(net63),
    .A2_N(_2592_),
    .B1(_2582_),
    .B2(net641),
    .X(_0317_));
 sky130_fd_sc_hd__a21o_1 _5796_ (.A1(net694),
    .A2(net99),
    .B1(_1711_),
    .X(_2593_));
 sky130_fd_sc_hd__mux2_1 _5797_ (.A0(_2593_),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[1] ),
    .S(net68),
    .X(_2594_));
 sky130_fd_sc_hd__a211o_1 _5798_ (.A1(net88),
    .A2(_2594_),
    .B1(_1728_),
    .C1(net78),
    .X(_2595_));
 sky130_fd_sc_hd__or3_1 _5799_ (.A(net119),
    .B(\z80.tv80s.di_reg[1] ),
    .C(_0685_),
    .X(_2596_));
 sky130_fd_sc_hd__and3_1 _5800_ (.A(\z80.tv80s.i_tv80_core.PC[1] ),
    .B(_2577_),
    .C(_2596_),
    .X(_2597_));
 sky130_fd_sc_hd__a21oi_1 _5801_ (.A1(_2577_),
    .A2(_2596_),
    .B1(\z80.tv80s.i_tv80_core.PC[1] ),
    .Y(_2598_));
 sky130_fd_sc_hd__or2_1 _5802_ (.A(_2597_),
    .B(_2598_),
    .X(_2599_));
 sky130_fd_sc_hd__and2_1 _5803_ (.A(_2589_),
    .B(_2599_),
    .X(_2600_));
 sky130_fd_sc_hd__nor2_1 _5804_ (.A(_2589_),
    .B(_2599_),
    .Y(_2601_));
 sky130_fd_sc_hd__nor2_1 _5805_ (.A(_2600_),
    .B(_2601_),
    .Y(_2602_));
 sky130_fd_sc_hd__a32o_1 _5806_ (.A1(_1730_),
    .A2(_2584_),
    .A3(_2595_),
    .B1(_2602_),
    .B2(net64),
    .X(_2603_));
 sky130_fd_sc_hd__a22o_1 _5807_ (.A1(net694),
    .A2(_2583_),
    .B1(_2603_),
    .B2(net63),
    .X(_0318_));
 sky130_fd_sc_hd__or3_1 _5808_ (.A(net119),
    .B(\z80.tv80s.di_reg[2] ),
    .C(_0685_),
    .X(_2604_));
 sky130_fd_sc_hd__and3_1 _5809_ (.A(\z80.tv80s.i_tv80_core.PC[2] ),
    .B(_2577_),
    .C(_2604_),
    .X(_2605_));
 sky130_fd_sc_hd__a21oi_1 _5810_ (.A1(_2577_),
    .A2(_2604_),
    .B1(\z80.tv80s.i_tv80_core.PC[2] ),
    .Y(_2606_));
 sky130_fd_sc_hd__or2_1 _5811_ (.A(_2605_),
    .B(_2606_),
    .X(_2607_));
 sky130_fd_sc_hd__o21ba_1 _5812_ (.A1(_2597_),
    .A2(_2601_),
    .B1_N(_2607_),
    .X(_2608_));
 sky130_fd_sc_hd__or3b_1 _5813_ (.A(_2597_),
    .B(_2601_),
    .C_N(_2607_),
    .X(_2609_));
 sky130_fd_sc_hd__nand2b_1 _5814_ (.A_N(_2608_),
    .B(_2609_),
    .Y(_2610_));
 sky130_fd_sc_hd__a21o_1 _5815_ (.A1(\z80.tv80s.i_tv80_core.PC[2] ),
    .A2(net99),
    .B1(_1733_),
    .X(_2611_));
 sky130_fd_sc_hd__mux2_1 _5816_ (.A0(_2611_),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[2] ),
    .S(_1681_),
    .X(_2612_));
 sky130_fd_sc_hd__nand2_1 _5817_ (.A(net88),
    .B(_2612_),
    .Y(_2613_));
 sky130_fd_sc_hd__a22o_1 _5818_ (.A1(_2880_),
    .A2(net78),
    .B1(_1749_),
    .B2(_2613_),
    .X(_2614_));
 sky130_fd_sc_hd__a22o_1 _5819_ (.A1(net64),
    .A2(_2610_),
    .B1(_2614_),
    .B2(_2584_),
    .X(_2615_));
 sky130_fd_sc_hd__o2bb2a_1 _5820_ (.A1_N(net63),
    .A2_N(_2615_),
    .B1(_2582_),
    .B2(net617),
    .X(_0319_));
 sky130_fd_sc_hd__or3_1 _5821_ (.A(net119),
    .B(\z80.tv80s.di_reg[3] ),
    .C(_0685_),
    .X(_2616_));
 sky130_fd_sc_hd__and3_1 _5822_ (.A(\z80.tv80s.i_tv80_core.PC[3] ),
    .B(_2577_),
    .C(_2616_),
    .X(_2617_));
 sky130_fd_sc_hd__a21oi_1 _5823_ (.A1(_2577_),
    .A2(_2616_),
    .B1(\z80.tv80s.i_tv80_core.PC[3] ),
    .Y(_2618_));
 sky130_fd_sc_hd__or2_1 _5824_ (.A(_2617_),
    .B(_2618_),
    .X(_2619_));
 sky130_fd_sc_hd__o21ba_1 _5825_ (.A1(_2605_),
    .A2(_2608_),
    .B1_N(_2619_),
    .X(_2620_));
 sky130_fd_sc_hd__or3b_1 _5826_ (.A(_2605_),
    .B(_2608_),
    .C_N(_2619_),
    .X(_2621_));
 sky130_fd_sc_hd__nand2b_1 _5827_ (.A_N(_2620_),
    .B(_2621_),
    .Y(_2622_));
 sky130_fd_sc_hd__mux2_1 _5828_ (.A0(\z80.tv80s.i_tv80_core.TmpAddr[3] ),
    .A1(\z80.tv80s.i_tv80_core.PC[3] ),
    .S(net99),
    .X(_2623_));
 sky130_fd_sc_hd__a22o_1 _5829_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[3] ),
    .A2(net68),
    .B1(net66),
    .B2(_2623_),
    .X(_2624_));
 sky130_fd_sc_hd__a21o_1 _5830_ (.A1(net88),
    .A2(_2624_),
    .B1(_1755_),
    .X(_2625_));
 sky130_fd_sc_hd__o21ai_1 _5831_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[3] ),
    .A2(net79),
    .B1(_2625_),
    .Y(_2626_));
 sky130_fd_sc_hd__a22o_1 _5832_ (.A1(net64),
    .A2(_2622_),
    .B1(_2626_),
    .B2(_2584_),
    .X(_2627_));
 sky130_fd_sc_hd__o2bb2a_1 _5833_ (.A1_N(net63),
    .A2_N(_2627_),
    .B1(_2582_),
    .B2(net595),
    .X(_0320_));
 sky130_fd_sc_hd__or3_1 _5834_ (.A(net119),
    .B(\z80.tv80s.di_reg[4] ),
    .C(_0685_),
    .X(_2628_));
 sky130_fd_sc_hd__and3_1 _5835_ (.A(\z80.tv80s.i_tv80_core.PC[4] ),
    .B(_2577_),
    .C(_2628_),
    .X(_2629_));
 sky130_fd_sc_hd__a21oi_1 _5836_ (.A1(_2577_),
    .A2(_2628_),
    .B1(\z80.tv80s.i_tv80_core.PC[4] ),
    .Y(_2630_));
 sky130_fd_sc_hd__or2_1 _5837_ (.A(_2629_),
    .B(_2630_),
    .X(_2631_));
 sky130_fd_sc_hd__o21ba_1 _5838_ (.A1(_2617_),
    .A2(_2620_),
    .B1_N(_2631_),
    .X(_2632_));
 sky130_fd_sc_hd__or3b_1 _5839_ (.A(_2617_),
    .B(_2620_),
    .C_N(_2631_),
    .X(_2633_));
 sky130_fd_sc_hd__nand2b_1 _5840_ (.A_N(_2632_),
    .B(_2633_),
    .Y(_2634_));
 sky130_fd_sc_hd__mux2_1 _5841_ (.A0(\z80.tv80s.i_tv80_core.TmpAddr[4] ),
    .A1(\z80.tv80s.i_tv80_core.PC[4] ),
    .S(net99),
    .X(_2635_));
 sky130_fd_sc_hd__a22o_1 _5842_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[4] ),
    .A2(net68),
    .B1(net66),
    .B2(_2635_),
    .X(_2636_));
 sky130_fd_sc_hd__a21o_1 _5843_ (.A1(net88),
    .A2(_2636_),
    .B1(_1772_),
    .X(_2637_));
 sky130_fd_sc_hd__o21ai_1 _5844_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[4] ),
    .A2(_1669_),
    .B1(_2637_),
    .Y(_2638_));
 sky130_fd_sc_hd__a22o_1 _5845_ (.A1(_2581_),
    .A2(_2634_),
    .B1(_2638_),
    .B2(_2584_),
    .X(_2639_));
 sky130_fd_sc_hd__o2bb2a_1 _5846_ (.A1_N(net63),
    .A2_N(_2639_),
    .B1(_2582_),
    .B2(net599),
    .X(_0321_));
 sky130_fd_sc_hd__a21o_1 _5847_ (.A1(\z80.tv80s.i_tv80_core.PC[5] ),
    .A2(net98),
    .B1(_1791_),
    .X(_2640_));
 sky130_fd_sc_hd__mux2_1 _5848_ (.A0(_2640_),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[5] ),
    .S(net67),
    .X(_2641_));
 sky130_fd_sc_hd__a21bo_1 _5849_ (.A1(net88),
    .A2(_2641_),
    .B1_N(_1790_),
    .X(_2642_));
 sky130_fd_sc_hd__mux2_1 _5850_ (.A0(\z80.tv80s.i_tv80_core.TmpAddr[5] ),
    .A1(_2642_),
    .S(net79),
    .X(_2643_));
 sky130_fd_sc_hd__or3_1 _5851_ (.A(net119),
    .B(\z80.tv80s.di_reg[5] ),
    .C(_0685_),
    .X(_2644_));
 sky130_fd_sc_hd__and3_1 _5852_ (.A(net577),
    .B(_2577_),
    .C(_2644_),
    .X(_2645_));
 sky130_fd_sc_hd__a21oi_1 _5853_ (.A1(_2577_),
    .A2(_2644_),
    .B1(\z80.tv80s.i_tv80_core.PC[5] ),
    .Y(_2646_));
 sky130_fd_sc_hd__or2_1 _5854_ (.A(_2645_),
    .B(_2646_),
    .X(_2647_));
 sky130_fd_sc_hd__nor3b_1 _5855_ (.A(_2629_),
    .B(_2632_),
    .C_N(_2647_),
    .Y(_2648_));
 sky130_fd_sc_hd__o21ba_1 _5856_ (.A1(_2629_),
    .A2(_2632_),
    .B1_N(_2647_),
    .X(_2649_));
 sky130_fd_sc_hd__nor2_1 _5857_ (.A(_2648_),
    .B(_2649_),
    .Y(_2650_));
 sky130_fd_sc_hd__a22o_1 _5858_ (.A1(_2584_),
    .A2(_2643_),
    .B1(_2650_),
    .B2(_2581_),
    .X(_2651_));
 sky130_fd_sc_hd__a22o_1 _5859_ (.A1(net577),
    .A2(_2583_),
    .B1(_2651_),
    .B2(_2570_),
    .X(_0322_));
 sky130_fd_sc_hd__a21o_1 _5860_ (.A1(\z80.tv80s.i_tv80_core.PC[6] ),
    .A2(_1685_),
    .B1(_1809_),
    .X(_2652_));
 sky130_fd_sc_hd__mux2_1 _5861_ (.A0(_2652_),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[6] ),
    .S(net68),
    .X(_2653_));
 sky130_fd_sc_hd__a21o_1 _5862_ (.A1(net88),
    .A2(_2653_),
    .B1(_1808_),
    .X(_2654_));
 sky130_fd_sc_hd__mux2_1 _5863_ (.A0(\z80.tv80s.i_tv80_core.TmpAddr[6] ),
    .A1(_2654_),
    .S(_1669_),
    .X(_2655_));
 sky130_fd_sc_hd__o21ba_1 _5864_ (.A1(net60),
    .A2(_2655_),
    .B1_N(_2581_),
    .X(_2656_));
 sky130_fd_sc_hd__o21a_1 _5865_ (.A1(net744),
    .A2(_0577_),
    .B1(_2656_),
    .X(_2657_));
 sky130_fd_sc_hd__or3_1 _5866_ (.A(net119),
    .B(\z80.tv80s.di_reg[6] ),
    .C(_0685_),
    .X(_2658_));
 sky130_fd_sc_hd__and3_1 _5867_ (.A(\z80.tv80s.i_tv80_core.PC[6] ),
    .B(_2577_),
    .C(_2658_),
    .X(_2659_));
 sky130_fd_sc_hd__inv_2 _5868_ (.A(_2659_),
    .Y(_2660_));
 sky130_fd_sc_hd__a21oi_1 _5869_ (.A1(_2577_),
    .A2(_2658_),
    .B1(\z80.tv80s.i_tv80_core.PC[6] ),
    .Y(_2661_));
 sky130_fd_sc_hd__or2_1 _5870_ (.A(_2659_),
    .B(_2661_),
    .X(_2662_));
 sky130_fd_sc_hd__o21bai_1 _5871_ (.A1(_2645_),
    .A2(_2649_),
    .B1_N(_2662_),
    .Y(_2663_));
 sky130_fd_sc_hd__or3b_1 _5872_ (.A(_2645_),
    .B(_2649_),
    .C_N(_2662_),
    .X(_2664_));
 sky130_fd_sc_hd__a31o_1 _5873_ (.A1(net64),
    .A2(_2663_),
    .A3(_2664_),
    .B1(_2657_),
    .X(_2665_));
 sky130_fd_sc_hd__mux2_1 _5874_ (.A0(net744),
    .A1(_2665_),
    .S(_2570_),
    .X(_0323_));
 sky130_fd_sc_hd__mux2_1 _5875_ (.A0(\z80.tv80s.i_tv80_core.TmpAddr[7] ),
    .A1(\z80.tv80s.i_tv80_core.PC[7] ),
    .S(net99),
    .X(_2666_));
 sky130_fd_sc_hd__a22o_1 _5876_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[7] ),
    .A2(net68),
    .B1(net65),
    .B2(_2666_),
    .X(_2667_));
 sky130_fd_sc_hd__a21bo_1 _5877_ (.A1(net87),
    .A2(_2667_),
    .B1_N(_1829_),
    .X(_2668_));
 sky130_fd_sc_hd__mux2_1 _5878_ (.A0(\z80.tv80s.i_tv80_core.TmpAddr[7] ),
    .A1(_2668_),
    .S(net79),
    .X(_2669_));
 sky130_fd_sc_hd__mux2_1 _5879_ (.A0(_2669_),
    .A1(net738),
    .S(net60),
    .X(_2670_));
 sky130_fd_sc_hd__o31a_2 _5880_ (.A1(net119),
    .A2(\z80.tv80s.di_reg[7] ),
    .A3(_0685_),
    .B1(_2577_),
    .X(_2671_));
 sky130_fd_sc_hd__and2_1 _5881_ (.A(\z80.tv80s.i_tv80_core.PC[7] ),
    .B(net77),
    .X(_2672_));
 sky130_fd_sc_hd__nor2_1 _5882_ (.A(\z80.tv80s.i_tv80_core.PC[7] ),
    .B(net77),
    .Y(_2673_));
 sky130_fd_sc_hd__or2_1 _5883_ (.A(_2672_),
    .B(_2673_),
    .X(_2674_));
 sky130_fd_sc_hd__and3_1 _5884_ (.A(_2660_),
    .B(_2663_),
    .C(_2674_),
    .X(_2675_));
 sky130_fd_sc_hd__a21oi_1 _5885_ (.A1(_2660_),
    .A2(_2663_),
    .B1(_2674_),
    .Y(_2676_));
 sky130_fd_sc_hd__nor2_1 _5886_ (.A(_2675_),
    .B(_2676_),
    .Y(_2677_));
 sky130_fd_sc_hd__mux2_1 _5887_ (.A0(_2670_),
    .A1(_2677_),
    .S(_2581_),
    .X(_2678_));
 sky130_fd_sc_hd__mux2_1 _5888_ (.A0(net738),
    .A1(_2678_),
    .S(net63),
    .X(_0324_));
 sky130_fd_sc_hd__xnor2_1 _5889_ (.A(\z80.tv80s.i_tv80_core.PC[8] ),
    .B(net77),
    .Y(_2679_));
 sky130_fd_sc_hd__or3b_1 _5890_ (.A(_2672_),
    .B(_2676_),
    .C_N(_2679_),
    .X(_2680_));
 sky130_fd_sc_hd__o21ba_1 _5891_ (.A1(_2672_),
    .A2(_2676_),
    .B1_N(_2679_),
    .X(_2681_));
 sky130_fd_sc_hd__mux2_1 _5892_ (.A0(\z80.tv80s.i_tv80_core.I[0] ),
    .A1(\z80.tv80s.i_tv80_core.PC[8] ),
    .S(net99),
    .X(_2682_));
 sky130_fd_sc_hd__a22o_1 _5893_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[8] ),
    .A2(net68),
    .B1(net65),
    .B2(_2682_),
    .X(_2683_));
 sky130_fd_sc_hd__nand2_1 _5894_ (.A(net87),
    .B(_2683_),
    .Y(_2684_));
 sky130_fd_sc_hd__a21oi_1 _5895_ (.A1(_1848_),
    .A2(_2684_),
    .B1(net78),
    .Y(_2685_));
 sky130_fd_sc_hd__a211o_1 _5896_ (.A1(\z80.tv80s.di_reg[0] ),
    .A2(net78),
    .B1(_2685_),
    .C1(net60),
    .X(_2686_));
 sky130_fd_sc_hd__o21ba_1 _5897_ (.A1(net808),
    .A2(_0577_),
    .B1_N(net64),
    .X(_2687_));
 sky130_fd_sc_hd__nand2_1 _5898_ (.A(net64),
    .B(_2680_),
    .Y(_2688_));
 sky130_fd_sc_hd__a2bb2o_1 _5899_ (.A1_N(_2681_),
    .A2_N(_2688_),
    .B1(_2686_),
    .B2(_2687_),
    .X(_2689_));
 sky130_fd_sc_hd__mux2_1 _5900_ (.A0(net808),
    .A1(_2689_),
    .S(net63),
    .X(_0325_));
 sky130_fd_sc_hd__xor2_1 _5901_ (.A(net788),
    .B(_2671_),
    .X(_2690_));
 sky130_fd_sc_hd__a21oi_1 _5902_ (.A1(\z80.tv80s.i_tv80_core.PC[8] ),
    .A2(net77),
    .B1(_2681_),
    .Y(_2691_));
 sky130_fd_sc_hd__xnor2_1 _5903_ (.A(_2690_),
    .B(_2691_),
    .Y(_2692_));
 sky130_fd_sc_hd__mux2_1 _5904_ (.A0(\z80.tv80s.i_tv80_core.I[1] ),
    .A1(\z80.tv80s.i_tv80_core.PC[9] ),
    .S(net98),
    .X(_2693_));
 sky130_fd_sc_hd__a22o_1 _5905_ (.A1(net611),
    .A2(net67),
    .B1(net65),
    .B2(_2693_),
    .X(_2694_));
 sky130_fd_sc_hd__a21bo_1 _5906_ (.A1(net87),
    .A2(_2694_),
    .B1_N(_1867_),
    .X(_2695_));
 sky130_fd_sc_hd__mux2_1 _5907_ (.A0(\z80.tv80s.di_reg[1] ),
    .A1(_2695_),
    .S(net79),
    .X(_2696_));
 sky130_fd_sc_hd__a22o_1 _5908_ (.A1(net64),
    .A2(_2692_),
    .B1(_2696_),
    .B2(_2584_),
    .X(_2697_));
 sky130_fd_sc_hd__a22o_1 _5909_ (.A1(net788),
    .A2(_2583_),
    .B1(_2697_),
    .B2(net63),
    .X(_0326_));
 sky130_fd_sc_hd__xnor2_1 _5910_ (.A(\z80.tv80s.i_tv80_core.PC[10] ),
    .B(net77),
    .Y(_2698_));
 sky130_fd_sc_hd__o21ai_1 _5911_ (.A1(\z80.tv80s.i_tv80_core.PC[8] ),
    .A2(\z80.tv80s.i_tv80_core.PC[9] ),
    .B1(_2671_),
    .Y(_2699_));
 sky130_fd_sc_hd__nand2_1 _5912_ (.A(_2681_),
    .B(_2690_),
    .Y(_2700_));
 sky130_fd_sc_hd__a21oi_1 _5913_ (.A1(_2699_),
    .A2(_2700_),
    .B1(_2698_),
    .Y(_2701_));
 sky130_fd_sc_hd__and3_1 _5914_ (.A(_2698_),
    .B(_2699_),
    .C(_2700_),
    .X(_2702_));
 sky130_fd_sc_hd__or2_1 _5915_ (.A(_2701_),
    .B(_2702_),
    .X(_2703_));
 sky130_fd_sc_hd__mux2_1 _5916_ (.A0(\z80.tv80s.i_tv80_core.I[2] ),
    .A1(\z80.tv80s.i_tv80_core.PC[10] ),
    .S(net98),
    .X(_2704_));
 sky130_fd_sc_hd__a22o_1 _5917_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[10] ),
    .A2(net67),
    .B1(net65),
    .B2(_2704_),
    .X(_2705_));
 sky130_fd_sc_hd__nand2_1 _5918_ (.A(net87),
    .B(_2705_),
    .Y(_2706_));
 sky130_fd_sc_hd__a21o_1 _5919_ (.A1(_1886_),
    .A2(_2706_),
    .B1(net78),
    .X(_2707_));
 sky130_fd_sc_hd__a32o_1 _5920_ (.A1(_1898_),
    .A2(_2584_),
    .A3(_2707_),
    .B1(_2703_),
    .B2(net64),
    .X(_2708_));
 sky130_fd_sc_hd__o2bb2a_1 _5921_ (.A1_N(net63),
    .A2_N(_2708_),
    .B1(_2582_),
    .B2(net806),
    .X(_0327_));
 sky130_fd_sc_hd__xnor2_1 _5922_ (.A(net799),
    .B(net77),
    .Y(_2709_));
 sky130_fd_sc_hd__a21o_1 _5923_ (.A1(\z80.tv80s.i_tv80_core.PC[10] ),
    .A2(net77),
    .B1(_2701_),
    .X(_2710_));
 sky130_fd_sc_hd__xnor2_1 _5924_ (.A(_2709_),
    .B(_2710_),
    .Y(_2711_));
 sky130_fd_sc_hd__mux2_1 _5925_ (.A0(\z80.tv80s.i_tv80_core.I[3] ),
    .A1(\z80.tv80s.i_tv80_core.PC[11] ),
    .S(net98),
    .X(_2712_));
 sky130_fd_sc_hd__a22o_1 _5926_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[11] ),
    .A2(net67),
    .B1(net65),
    .B2(_2712_),
    .X(_2713_));
 sky130_fd_sc_hd__a21bo_1 _5927_ (.A1(net87),
    .A2(_2713_),
    .B1_N(_1904_),
    .X(_2714_));
 sky130_fd_sc_hd__mux2_1 _5928_ (.A0(\z80.tv80s.di_reg[3] ),
    .A1(_2714_),
    .S(net79),
    .X(_2715_));
 sky130_fd_sc_hd__mux2_1 _5929_ (.A0(_2715_),
    .A1(net799),
    .S(net60),
    .X(_2716_));
 sky130_fd_sc_hd__mux2_1 _5930_ (.A0(_2716_),
    .A1(_2711_),
    .S(net64),
    .X(_2717_));
 sky130_fd_sc_hd__mux2_1 _5931_ (.A0(net799),
    .A1(_2717_),
    .S(net63),
    .X(_0328_));
 sky130_fd_sc_hd__nand2_1 _5932_ (.A(net772),
    .B(net77),
    .Y(_2718_));
 sky130_fd_sc_hd__or2_1 _5933_ (.A(net772),
    .B(net77),
    .X(_2719_));
 sky130_fd_sc_hd__nand2_1 _5934_ (.A(_2718_),
    .B(_2719_),
    .Y(_2720_));
 sky130_fd_sc_hd__o41ai_1 _5935_ (.A1(\z80.tv80s.i_tv80_core.PC[8] ),
    .A2(\z80.tv80s.i_tv80_core.PC[9] ),
    .A3(\z80.tv80s.i_tv80_core.PC[10] ),
    .A4(\z80.tv80s.i_tv80_core.PC[11] ),
    .B1(net77),
    .Y(_2721_));
 sky130_fd_sc_hd__o31a_1 _5936_ (.A1(_2698_),
    .A2(_2700_),
    .A3(_2709_),
    .B1(_2721_),
    .X(_2722_));
 sky130_fd_sc_hd__xor2_1 _5937_ (.A(_2720_),
    .B(_2722_),
    .X(_2723_));
 sky130_fd_sc_hd__mux2_1 _5938_ (.A0(\z80.tv80s.i_tv80_core.I[4] ),
    .A1(\z80.tv80s.i_tv80_core.PC[12] ),
    .S(net98),
    .X(_2724_));
 sky130_fd_sc_hd__a22o_1 _5939_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[12] ),
    .A2(net67),
    .B1(net65),
    .B2(_2724_),
    .X(_2725_));
 sky130_fd_sc_hd__a21bo_1 _5940_ (.A1(net87),
    .A2(_2725_),
    .B1_N(_1923_),
    .X(_2726_));
 sky130_fd_sc_hd__mux2_1 _5941_ (.A0(\z80.tv80s.di_reg[4] ),
    .A1(_2726_),
    .S(net79),
    .X(_2727_));
 sky130_fd_sc_hd__mux2_1 _5942_ (.A0(_2727_),
    .A1(net772),
    .S(_0576_),
    .X(_2728_));
 sky130_fd_sc_hd__mux2_1 _5943_ (.A0(_2728_),
    .A1(_2723_),
    .S(net64),
    .X(_2729_));
 sky130_fd_sc_hd__mux2_1 _5944_ (.A0(net772),
    .A1(_2729_),
    .S(net63),
    .X(_0329_));
 sky130_fd_sc_hd__mux2_1 _5945_ (.A0(\z80.tv80s.i_tv80_core.I[5] ),
    .A1(\z80.tv80s.i_tv80_core.PC[13] ),
    .S(net98),
    .X(_2730_));
 sky130_fd_sc_hd__a22o_1 _5946_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[13] ),
    .A2(net67),
    .B1(net65),
    .B2(_2730_),
    .X(_2731_));
 sky130_fd_sc_hd__a21bo_1 _5947_ (.A1(net87),
    .A2(_2731_),
    .B1_N(_1944_),
    .X(_2732_));
 sky130_fd_sc_hd__mux2_1 _5948_ (.A0(\z80.tv80s.di_reg[5] ),
    .A1(_2732_),
    .S(net79),
    .X(_2733_));
 sky130_fd_sc_hd__nand2_1 _5949_ (.A(net780),
    .B(net77),
    .Y(_2734_));
 sky130_fd_sc_hd__nor2_1 _5950_ (.A(\z80.tv80s.i_tv80_core.PC[13] ),
    .B(net77),
    .Y(_2735_));
 sky130_fd_sc_hd__or2_1 _5951_ (.A(net780),
    .B(net77),
    .X(_2736_));
 sky130_fd_sc_hd__nand2_1 _5952_ (.A(_2734_),
    .B(_2736_),
    .Y(_2737_));
 sky130_fd_sc_hd__o21a_1 _5953_ (.A1(_2720_),
    .A2(_2722_),
    .B1(_2718_),
    .X(_2738_));
 sky130_fd_sc_hd__xor2_1 _5954_ (.A(_2737_),
    .B(_2738_),
    .X(_2739_));
 sky130_fd_sc_hd__a22o_1 _5955_ (.A1(_2584_),
    .A2(_2733_),
    .B1(_2739_),
    .B2(net64),
    .X(_2740_));
 sky130_fd_sc_hd__a22o_1 _5956_ (.A1(net780),
    .A2(_2583_),
    .B1(_2740_),
    .B2(net63),
    .X(_0330_));
 sky130_fd_sc_hd__and2_1 _5957_ (.A(\z80.tv80s.i_tv80_core.PC[14] ),
    .B(net77),
    .X(_2741_));
 sky130_fd_sc_hd__nor2_1 _5958_ (.A(\z80.tv80s.i_tv80_core.PC[14] ),
    .B(net77),
    .Y(_2742_));
 sky130_fd_sc_hd__or2_1 _5959_ (.A(_2741_),
    .B(_2742_),
    .X(_2743_));
 sky130_fd_sc_hd__o21a_1 _5960_ (.A1(_2735_),
    .A2(_2738_),
    .B1(_2734_),
    .X(_2744_));
 sky130_fd_sc_hd__xnor2_1 _5961_ (.A(_2743_),
    .B(_2744_),
    .Y(_2745_));
 sky130_fd_sc_hd__mux2_1 _5962_ (.A0(\z80.tv80s.i_tv80_core.I[6] ),
    .A1(\z80.tv80s.i_tv80_core.PC[14] ),
    .S(net98),
    .X(_2746_));
 sky130_fd_sc_hd__a22o_1 _5963_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[14] ),
    .A2(net67),
    .B1(net65),
    .B2(_2746_),
    .X(_2747_));
 sky130_fd_sc_hd__nand2_1 _5964_ (.A(net87),
    .B(_2747_),
    .Y(_2748_));
 sky130_fd_sc_hd__a21o_1 _5965_ (.A1(_1961_),
    .A2(_2748_),
    .B1(net78),
    .X(_2749_));
 sky130_fd_sc_hd__a32o_1 _5966_ (.A1(_1975_),
    .A2(_2584_),
    .A3(_2749_),
    .B1(_2745_),
    .B2(net64),
    .X(_2750_));
 sky130_fd_sc_hd__o2bb2a_1 _5967_ (.A1_N(net63),
    .A2_N(_2750_),
    .B1(_2582_),
    .B2(net766),
    .X(_0331_));
 sky130_fd_sc_hd__o21ba_1 _5968_ (.A1(_2742_),
    .A2(_2744_),
    .B1_N(_2741_),
    .X(_2751_));
 sky130_fd_sc_hd__xor2_1 _5969_ (.A(net757),
    .B(_2751_),
    .X(_2752_));
 sky130_fd_sc_hd__xnor2_1 _5970_ (.A(net77),
    .B(_2752_),
    .Y(_2753_));
 sky130_fd_sc_hd__mux2_1 _5971_ (.A0(\z80.tv80s.i_tv80_core.I[7] ),
    .A1(\z80.tv80s.i_tv80_core.PC[15] ),
    .S(net98),
    .X(_2754_));
 sky130_fd_sc_hd__a22o_1 _5972_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[15] ),
    .A2(net67),
    .B1(net65),
    .B2(_2754_),
    .X(_2755_));
 sky130_fd_sc_hd__a21bo_1 _5973_ (.A1(net87),
    .A2(_2755_),
    .B1_N(_1981_),
    .X(_2756_));
 sky130_fd_sc_hd__mux2_1 _5974_ (.A0(\z80.tv80s.di_reg[7] ),
    .A1(_2756_),
    .S(net79),
    .X(_2757_));
 sky130_fd_sc_hd__mux2_1 _5975_ (.A0(_2757_),
    .A1(net757),
    .S(_0576_),
    .X(_2758_));
 sky130_fd_sc_hd__mux2_1 _5976_ (.A0(_2758_),
    .A1(_2753_),
    .S(net64),
    .X(_2759_));
 sky130_fd_sc_hd__mux2_1 _5977_ (.A0(net757),
    .A1(_2759_),
    .S(net63),
    .X(_0332_));
 sky130_fd_sc_hd__nor2_1 _5978_ (.A(net129),
    .B(net716),
    .Y(_2760_));
 sky130_fd_sc_hd__nor2_1 _5979_ (.A(_0034_),
    .B(net770),
    .Y(_2761_));
 sky130_fd_sc_hd__nor2_1 _5980_ (.A(_2842_),
    .B(net698),
    .Y(_2762_));
 sky130_fd_sc_hd__or3_1 _5981_ (.A(net797),
    .B(net770),
    .C(net698),
    .X(_2763_));
 sky130_fd_sc_hd__nand3_1 _5982_ (.A(net797),
    .B(net770),
    .C(net698),
    .Y(_2764_));
 sky130_fd_sc_hd__a31oi_1 _5983_ (.A1(net129),
    .A2(_2763_),
    .A3(_2764_),
    .B1(_2760_),
    .Y(_2765_));
 sky130_fd_sc_hd__a22o_1 _5984_ (.A1(net133),
    .A2(_0580_),
    .B1(_0721_),
    .B2(_2765_),
    .X(_0333_));
 sky130_fd_sc_hd__or3b_1 _5985_ (.A(_0035_),
    .B(net698),
    .C_N(_0034_),
    .X(_2766_));
 sky130_fd_sc_hd__a21oi_1 _5986_ (.A1(net129),
    .A2(_2766_),
    .B1(_2984_),
    .Y(_2767_));
 sky130_fd_sc_hd__a32o_1 _5987_ (.A1(_0720_),
    .A2(_0721_),
    .A3(_2767_),
    .B1(_0580_),
    .B2(net131),
    .X(_0334_));
 sky130_fd_sc_hd__and2b_1 _5988_ (.A_N(_0034_),
    .B(net770),
    .X(_2768_));
 sky130_fd_sc_hd__a22o_1 _5989_ (.A1(net131),
    .A2(_2760_),
    .B1(_2762_),
    .B2(_2768_),
    .X(_2769_));
 sky130_fd_sc_hd__a22o_1 _5990_ (.A1(net130),
    .A2(_0580_),
    .B1(_0721_),
    .B2(_2769_),
    .X(_0335_));
 sky130_fd_sc_hd__a32o_1 _5991_ (.A1(_0034_),
    .A2(_0035_),
    .A3(_2762_),
    .B1(net130),
    .B2(_2842_),
    .X(_2770_));
 sky130_fd_sc_hd__a32o_1 _5992_ (.A1(_0720_),
    .A2(_0721_),
    .A3(_2770_),
    .B1(_0580_),
    .B2(net692),
    .X(_0336_));
 sky130_fd_sc_hd__a32o_1 _5993_ (.A1(net129),
    .A2(net698),
    .A3(net771),
    .B1(_2760_),
    .B2(net692),
    .X(_2771_));
 sky130_fd_sc_hd__a22o_1 _5994_ (.A1(net523),
    .A2(_0580_),
    .B1(_0721_),
    .B2(_2771_),
    .X(_0337_));
 sky130_fd_sc_hd__and4b_1 _5995_ (.A_N(net770),
    .B(net698),
    .C(net129),
    .D(net797),
    .X(_2772_));
 sky130_fd_sc_hd__a21oi_1 _5996_ (.A1(net523),
    .A2(_2760_),
    .B1(_2772_),
    .Y(_2773_));
 sky130_fd_sc_hd__o2bb2a_1 _5997_ (.A1_N(_0721_),
    .A2_N(_2773_),
    .B1(net609),
    .B2(_0581_),
    .X(_0338_));
 sky130_fd_sc_hd__a31o_1 _5998_ (.A1(net129),
    .A2(net698),
    .A3(_2768_),
    .B1(_0584_),
    .X(_2774_));
 sky130_fd_sc_hd__a32o_1 _5999_ (.A1(_0720_),
    .A2(_0721_),
    .A3(net699),
    .B1(_0580_),
    .B2(net129),
    .X(_0339_));
 sky130_fd_sc_hd__a21o_1 _6000_ (.A1(net778),
    .A2(_0722_),
    .B1(_0732_),
    .X(_0340_));
 sky130_fd_sc_hd__o21a_1 _6001_ (.A1(net124),
    .A2(_0579_),
    .B1(net221),
    .X(_0341_));
 sky130_fd_sc_hd__a22o_1 _6002_ (.A1(\z80.tv80s.i_tv80_core.NMICycle ),
    .A2(_0722_),
    .B1(_0723_),
    .B2(net518),
    .X(_0342_));
 sky130_fd_sc_hd__or2_4 _6003_ (.A(_0880_),
    .B(_1430_),
    .X(_2775_));
 sky130_fd_sc_hd__mux2_1 _6004_ (.A0(_1435_),
    .A1(net470),
    .S(_2775_),
    .X(_0343_));
 sky130_fd_sc_hd__mux2_1 _6005_ (.A0(_1446_),
    .A1(net486),
    .S(_2775_),
    .X(_0344_));
 sky130_fd_sc_hd__mux2_1 _6006_ (.A0(_1457_),
    .A1(net514),
    .S(_2775_),
    .X(_0345_));
 sky130_fd_sc_hd__mux2_1 _6007_ (.A0(_1463_),
    .A1(net375),
    .S(_2775_),
    .X(_0346_));
 sky130_fd_sc_hd__mux2_1 _6008_ (.A0(_1468_),
    .A1(net516),
    .S(_2775_),
    .X(_0347_));
 sky130_fd_sc_hd__mux2_1 _6009_ (.A0(_1474_),
    .A1(net466),
    .S(_2775_),
    .X(_0348_));
 sky130_fd_sc_hd__mux2_1 _6010_ (.A0(_1481_),
    .A1(net389),
    .S(_2775_),
    .X(_0349_));
 sky130_fd_sc_hd__mux2_1 _6011_ (.A0(_1487_),
    .A1(net520),
    .S(_2775_),
    .X(_0350_));
 sky130_fd_sc_hd__mux2_1 _6012_ (.A0(net13),
    .A1(net836),
    .S(_0604_),
    .X(_0351_));
 sky130_fd_sc_hd__mux2_1 _6013_ (.A0(net12),
    .A1(net838),
    .S(_0604_),
    .X(_0352_));
 sky130_fd_sc_hd__mux2_1 _6014_ (.A0(net10),
    .A1(net846),
    .S(_0604_),
    .X(_0353_));
 sky130_fd_sc_hd__mux2_1 _6015_ (.A0(net7),
    .A1(net844),
    .S(_0604_),
    .X(_0354_));
 sky130_fd_sc_hd__mux2_1 _6016_ (.A0(net6),
    .A1(net841),
    .S(_0604_),
    .X(_0355_));
 sky130_fd_sc_hd__mux2_1 _6017_ (.A0(net8),
    .A1(net840),
    .S(_0604_),
    .X(_0356_));
 sky130_fd_sc_hd__mux2_1 _6018_ (.A0(net9),
    .A1(net847),
    .S(_0604_),
    .X(_0357_));
 sky130_fd_sc_hd__mux2_1 _6019_ (.A0(net11),
    .A1(net848),
    .S(_0604_),
    .X(_0358_));
 sky130_fd_sc_hd__o32a_1 _6020_ (.A1(_2849_),
    .A2(net405),
    .A3(_0485_),
    .B1(_0708_),
    .B2(net340),
    .X(_2776_));
 sky130_fd_sc_hd__mux2_1 _6021_ (.A0(_2858_),
    .A1(_2776_),
    .S(net60),
    .X(_2777_));
 sky130_fd_sc_hd__nand2_4 _6022_ (.A(_0734_),
    .B(_2777_),
    .Y(_2778_));
 sky130_fd_sc_hd__nor2_2 _6023_ (.A(_0577_),
    .B(_2778_),
    .Y(_2779_));
 sky130_fd_sc_hd__a22o_1 _6024_ (.A1(\z80.tv80s.i_tv80_core.ts[0] ),
    .A2(_2778_),
    .B1(_2779_),
    .B2(net265),
    .X(_0359_));
 sky130_fd_sc_hd__or2_1 _6025_ (.A(net605),
    .B(_0574_),
    .X(_2780_));
 sky130_fd_sc_hd__mux2_1 _6026_ (.A0(_2780_),
    .A1(net573),
    .S(_2778_),
    .X(_0360_));
 sky130_fd_sc_hd__a22o_1 _6027_ (.A1(\z80.tv80s.i_tv80_core.ts[2] ),
    .A2(_2778_),
    .B1(_2779_),
    .B2(net573),
    .X(_0361_));
 sky130_fd_sc_hd__a22o_1 _6028_ (.A1(net122),
    .A2(_2778_),
    .B1(_2779_),
    .B2(net829),
    .X(_0362_));
 sky130_fd_sc_hd__a22o_1 _6029_ (.A1(net363),
    .A2(_2778_),
    .B1(_2779_),
    .B2(net122),
    .X(_0363_));
 sky130_fd_sc_hd__a22o_1 _6030_ (.A1(net297),
    .A2(_2778_),
    .B1(_2779_),
    .B2(net363),
    .X(_0364_));
 sky130_fd_sc_hd__a22o_1 _6031_ (.A1(net265),
    .A2(_2778_),
    .B1(_2779_),
    .B2(net297),
    .X(_0365_));
 sky130_fd_sc_hd__or3_1 _6032_ (.A(net508),
    .B(net501),
    .C(_2874_),
    .X(_2781_));
 sky130_fd_sc_hd__or4b_4 _6033_ (.A(net633),
    .B(_2875_),
    .C(_2781_),
    .D_N(_0781_),
    .X(_2782_));
 sky130_fd_sc_hd__a21oi_2 _6034_ (.A1(net136),
    .A2(\z80.tv80s.i_tv80_core.ts[4] ),
    .B1(_0603_),
    .Y(_2783_));
 sky130_fd_sc_hd__nor2_2 _6035_ (.A(_0763_),
    .B(_2783_),
    .Y(_2784_));
 sky130_fd_sc_hd__or2_4 _6036_ (.A(_0763_),
    .B(_2783_),
    .X(_2785_));
 sky130_fd_sc_hd__nand2_1 _6037_ (.A(net93),
    .B(_2784_),
    .Y(_2786_));
 sky130_fd_sc_hd__a21oi_1 _6038_ (.A1(_1416_),
    .A2(_2785_),
    .B1(net100),
    .Y(_2787_));
 sky130_fd_sc_hd__inv_2 _6039_ (.A(_2787_),
    .Y(_2788_));
 sky130_fd_sc_hd__a21oi_4 _6040_ (.A1(_2782_),
    .A2(_2788_),
    .B1(net123),
    .Y(_2789_));
 sky130_fd_sc_hd__o22a_1 _6041_ (.A1(_1416_),
    .A2(_1673_),
    .B1(_2264_),
    .B2(_2785_),
    .X(_2790_));
 sky130_fd_sc_hd__o21a_1 _6042_ (.A1(net101),
    .A2(_2790_),
    .B1(_2782_),
    .X(_2791_));
 sky130_fd_sc_hd__nor2_1 _6043_ (.A(_0856_),
    .B(_2782_),
    .Y(_2792_));
 sky130_fd_sc_hd__o32a_1 _6044_ (.A1(net124),
    .A2(_2791_),
    .A3(_2792_),
    .B1(net637),
    .B2(_2789_),
    .X(_0366_));
 sky130_fd_sc_hd__o22a_1 _6045_ (.A1(_1416_),
    .A2(_1715_),
    .B1(_2282_),
    .B2(_2785_),
    .X(_2793_));
 sky130_fd_sc_hd__o21a_1 _6046_ (.A1(net101),
    .A2(_2793_),
    .B1(_2782_),
    .X(_2794_));
 sky130_fd_sc_hd__nor2_1 _6047_ (.A(_1014_),
    .B(_2782_),
    .Y(_2795_));
 sky130_fd_sc_hd__o32a_1 _6048_ (.A1(net124),
    .A2(_2794_),
    .A3(_2795_),
    .B1(net680),
    .B2(_2789_),
    .X(_0367_));
 sky130_fd_sc_hd__o22a_1 _6049_ (.A1(_1416_),
    .A2(_1736_),
    .B1(_2293_),
    .B2(_2785_),
    .X(_2796_));
 sky130_fd_sc_hd__o21a_1 _6050_ (.A1(net101),
    .A2(_2796_),
    .B1(_2782_),
    .X(_2797_));
 sky130_fd_sc_hd__nor2_1 _6051_ (.A(_1066_),
    .B(_2782_),
    .Y(_2798_));
 sky130_fd_sc_hd__o32a_1 _6052_ (.A1(net123),
    .A2(_2797_),
    .A3(_2798_),
    .B1(net713),
    .B2(_2789_),
    .X(_0368_));
 sky130_fd_sc_hd__o22a_1 _6053_ (.A1(_1416_),
    .A2(_1754_),
    .B1(_2304_),
    .B2(_2785_),
    .X(_2799_));
 sky130_fd_sc_hd__o21a_1 _6054_ (.A1(net100),
    .A2(_2799_),
    .B1(_2782_),
    .X(_2800_));
 sky130_fd_sc_hd__nor2_1 _6055_ (.A(_1100_),
    .B(_2782_),
    .Y(_2801_));
 sky130_fd_sc_hd__o32a_1 _6056_ (.A1(net123),
    .A2(_2800_),
    .A3(_2801_),
    .B1(net703),
    .B2(_2789_),
    .X(_0369_));
 sky130_fd_sc_hd__o22a_1 _6057_ (.A1(_1416_),
    .A2(_1771_),
    .B1(_2316_),
    .B2(_2785_),
    .X(_2802_));
 sky130_fd_sc_hd__o21a_1 _6058_ (.A1(net100),
    .A2(_2802_),
    .B1(_2782_),
    .X(_2803_));
 sky130_fd_sc_hd__nor2_1 _6059_ (.A(_1150_),
    .B(_2782_),
    .Y(_2804_));
 sky130_fd_sc_hd__o32a_1 _6060_ (.A1(net123),
    .A2(_2803_),
    .A3(_2804_),
    .B1(net662),
    .B2(_2789_),
    .X(_0370_));
 sky130_fd_sc_hd__o22a_1 _6061_ (.A1(_1416_),
    .A2(_1789_),
    .B1(_2328_),
    .B2(_2785_),
    .X(_2805_));
 sky130_fd_sc_hd__o21a_1 _6062_ (.A1(net100),
    .A2(_2805_),
    .B1(_2782_),
    .X(_2806_));
 sky130_fd_sc_hd__nor2_1 _6063_ (.A(_1191_),
    .B(_2782_),
    .Y(_2807_));
 sky130_fd_sc_hd__o32a_1 _6064_ (.A1(net123),
    .A2(_2806_),
    .A3(_2807_),
    .B1(net718),
    .B2(_2789_),
    .X(_0371_));
 sky130_fd_sc_hd__o22a_1 _6065_ (.A1(_1416_),
    .A2(_1807_),
    .B1(_2340_),
    .B2(_2785_),
    .X(_2808_));
 sky130_fd_sc_hd__o21a_1 _6066_ (.A1(net100),
    .A2(_2808_),
    .B1(_2782_),
    .X(_2809_));
 sky130_fd_sc_hd__nor2_1 _6067_ (.A(_1245_),
    .B(_2782_),
    .Y(_2810_));
 sky130_fd_sc_hd__o32a_1 _6068_ (.A1(net123),
    .A2(_2809_),
    .A3(_2810_),
    .B1(net660),
    .B2(_2789_),
    .X(_0372_));
 sky130_fd_sc_hd__a22o_1 _6069_ (.A1(_1415_),
    .A2(_1827_),
    .B1(_2351_),
    .B2(_2784_),
    .X(_2811_));
 sky130_fd_sc_hd__nand2_1 _6070_ (.A(net93),
    .B(_2811_),
    .Y(_2812_));
 sky130_fd_sc_hd__mux2_1 _6071_ (.A0(_1295_),
    .A1(_2812_),
    .S(_2782_),
    .X(_2813_));
 sky130_fd_sc_hd__o22a_1 _6072_ (.A1(net798),
    .A2(_2789_),
    .B1(_2813_),
    .B2(net123),
    .X(_0373_));
 sky130_fd_sc_hd__or2_4 _6073_ (.A(_1995_),
    .B(_2781_),
    .X(_2814_));
 sky130_fd_sc_hd__o2bb2a_1 _6074_ (.A1_N(_2361_),
    .A2_N(_2784_),
    .B1(_1416_),
    .B2(_1847_),
    .X(_2815_));
 sky130_fd_sc_hd__o21a_1 _6075_ (.A1(net100),
    .A2(_2815_),
    .B1(_2814_),
    .X(_2816_));
 sky130_fd_sc_hd__nor2_1 _6076_ (.A(_0856_),
    .B(_2814_),
    .Y(_2817_));
 sky130_fd_sc_hd__a21oi_4 _6077_ (.A1(_2788_),
    .A2(_2814_),
    .B1(net123),
    .Y(_2818_));
 sky130_fd_sc_hd__o32a_1 _6078_ (.A1(net123),
    .A2(_2816_),
    .A3(_2817_),
    .B1(_2818_),
    .B2(net664),
    .X(_0374_));
 sky130_fd_sc_hd__o22a_1 _6079_ (.A1(_1416_),
    .A2(_1866_),
    .B1(_2375_),
    .B2(_2785_),
    .X(_2819_));
 sky130_fd_sc_hd__o21a_1 _6080_ (.A1(net100),
    .A2(_2819_),
    .B1(_2814_),
    .X(_2820_));
 sky130_fd_sc_hd__nor2_1 _6081_ (.A(_1014_),
    .B(_2814_),
    .Y(_2821_));
 sky130_fd_sc_hd__o32a_1 _6082_ (.A1(net123),
    .A2(_2820_),
    .A3(_2821_),
    .B1(net740),
    .B2(_2818_),
    .X(_0375_));
 sky130_fd_sc_hd__o22a_1 _6083_ (.A1(_1416_),
    .A2(_1885_),
    .B1(_2385_),
    .B2(_2785_),
    .X(_2822_));
 sky130_fd_sc_hd__o21a_1 _6084_ (.A1(net100),
    .A2(_2822_),
    .B1(_2814_),
    .X(_2823_));
 sky130_fd_sc_hd__nor2_1 _6085_ (.A(_1066_),
    .B(_2814_),
    .Y(_2824_));
 sky130_fd_sc_hd__o32a_1 _6086_ (.A1(net123),
    .A2(_2823_),
    .A3(_2824_),
    .B1(net583),
    .B2(_2818_),
    .X(_0376_));
 sky130_fd_sc_hd__o22a_1 _6087_ (.A1(_1416_),
    .A2(_1903_),
    .B1(_2393_),
    .B2(_2785_),
    .X(_2825_));
 sky130_fd_sc_hd__o21a_1 _6088_ (.A1(net100),
    .A2(_2825_),
    .B1(_2814_),
    .X(_2826_));
 sky130_fd_sc_hd__nor2_1 _6089_ (.A(_1100_),
    .B(_2814_),
    .Y(_2827_));
 sky130_fd_sc_hd__o32a_1 _6090_ (.A1(net123),
    .A2(_2826_),
    .A3(_2827_),
    .B1(net742),
    .B2(_2818_),
    .X(_0377_));
 sky130_fd_sc_hd__o2bb2a_1 _6091_ (.A1_N(_2403_),
    .A2_N(_2784_),
    .B1(_1416_),
    .B2(_1922_),
    .X(_2828_));
 sky130_fd_sc_hd__o21a_1 _6092_ (.A1(net100),
    .A2(_2828_),
    .B1(_2814_),
    .X(_2829_));
 sky130_fd_sc_hd__nor2_1 _6093_ (.A(_1150_),
    .B(_2814_),
    .Y(_2830_));
 sky130_fd_sc_hd__o32a_1 _6094_ (.A1(net123),
    .A2(_2829_),
    .A3(_2830_),
    .B1(net755),
    .B2(_2818_),
    .X(_0378_));
 sky130_fd_sc_hd__o22a_1 _6095_ (.A1(_1416_),
    .A2(_1943_),
    .B1(_2414_),
    .B2(_2785_),
    .X(_2831_));
 sky130_fd_sc_hd__o21a_1 _6096_ (.A1(net100),
    .A2(_2831_),
    .B1(_2814_),
    .X(_2832_));
 sky130_fd_sc_hd__nor2_1 _6097_ (.A(_1191_),
    .B(_2814_),
    .Y(_2833_));
 sky130_fd_sc_hd__o32a_1 _6098_ (.A1(net123),
    .A2(_2832_),
    .A3(_2833_),
    .B1(net688),
    .B2(_2818_),
    .X(_0379_));
 sky130_fd_sc_hd__o22a_1 _6099_ (.A1(net817),
    .A2(_2784_),
    .B1(_2786_),
    .B2(_2423_),
    .X(_2834_));
 sky130_fd_sc_hd__or2_1 _6100_ (.A(_1415_),
    .B(_2834_),
    .X(_2835_));
 sky130_fd_sc_hd__or3_1 _6101_ (.A(net100),
    .B(_1416_),
    .C(_1960_),
    .X(_2836_));
 sky130_fd_sc_hd__o211a_1 _6102_ (.A1(net817),
    .A2(net93),
    .B1(_2814_),
    .C1(_2836_),
    .X(_2837_));
 sky130_fd_sc_hd__a2bb2o_1 _6103_ (.A1_N(_1245_),
    .A2_N(_2814_),
    .B1(_2835_),
    .B2(_2837_),
    .X(_2838_));
 sky130_fd_sc_hd__mux2_1 _6104_ (.A0(net817),
    .A1(_2838_),
    .S(net112),
    .X(_0380_));
 sky130_fd_sc_hd__o22a_1 _6105_ (.A1(_1416_),
    .A2(_1980_),
    .B1(_2430_),
    .B2(_2785_),
    .X(_2839_));
 sky130_fd_sc_hd__o22a_1 _6106_ (.A1(net814),
    .A2(_2787_),
    .B1(_2839_),
    .B2(net100),
    .X(_2840_));
 sky130_fd_sc_hd__mux2_1 _6107_ (.A0(_1295_),
    .A1(_2840_),
    .S(_2814_),
    .X(_2841_));
 sky130_fd_sc_hd__mux2_1 _6108_ (.A0(net814),
    .A1(_2841_),
    .S(net27),
    .X(_0381_));
 sky130_fd_sc_hd__inv_2 _6109__2 (.A(clknet_leaf_11_wb_clk_i),
    .Y(net219));
 sky130_fd_sc_hd__inv_2 _6110__3 (.A(clknet_leaf_7_wb_clk_i),
    .Y(net220));
 sky130_fd_sc_hd__dfxtp_1 _6111_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(net458),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6112_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(net453),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6113_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(_0042_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6114_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(_0043_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6115_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(_0044_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6116_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(_0045_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6117_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(_0046_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6118_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(net455),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6119_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net226),
    .Q(\z80.tv80s.i_tv80_core.RegAddrA_r[2] ));
 sky130_fd_sc_hd__dfrtp_1 _6120_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(net559),
    .RESET_B(net173),
    .Q(\z80.tv80s.i_tv80_core.R[0] ));
 sky130_fd_sc_hd__dfrtp_1 _6121_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(net616),
    .RESET_B(net173),
    .Q(\z80.tv80s.i_tv80_core.R[1] ));
 sky130_fd_sc_hd__dfrtp_1 _6122_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(net545),
    .RESET_B(net174),
    .Q(\z80.tv80s.i_tv80_core.R[2] ));
 sky130_fd_sc_hd__dfrtp_1 _6123_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(net528),
    .RESET_B(net173),
    .Q(\z80.tv80s.i_tv80_core.R[3] ));
 sky130_fd_sc_hd__dfrtp_1 _6124_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(net614),
    .RESET_B(net173),
    .Q(\z80.tv80s.i_tv80_core.R[4] ));
 sky130_fd_sc_hd__dfrtp_1 _6125_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(net565),
    .RESET_B(net174),
    .Q(\z80.tv80s.i_tv80_core.R[5] ));
 sky130_fd_sc_hd__dfrtp_1 _6126_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(net685),
    .RESET_B(net173),
    .Q(\z80.tv80s.i_tv80_core.R[6] ));
 sky130_fd_sc_hd__dfxtp_1 _6127_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net553),
    .Q(\z80.tv80s.i_tv80_core.RegAddrB_r[2] ));
 sky130_fd_sc_hd__dfxtp_1 _6128_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(net598),
    .Q(\z80.tv80s.i_tv80_core.RegAddrC[2] ));
 sky130_fd_sc_hd__dfxtp_1 _6129_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(_0058_),
    .Q(\z80.tv80s.i_tv80_core.RegAddrC[1] ));
 sky130_fd_sc_hd__dfrtp_1 _6130_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net820),
    .RESET_B(net180),
    .Q(\z80.tv80s.i_tv80_core.mcycles[1] ));
 sky130_fd_sc_hd__dfrtp_1 _6131_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net280),
    .RESET_B(net180),
    .Q(\z80.tv80s.i_tv80_core.mcycles[2] ));
 sky130_fd_sc_hd__dfrtp_1 _6132_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net549),
    .RESET_B(net177),
    .Q(\z80.tv80s.i_tv80_core.mcycles[4] ));
 sky130_fd_sc_hd__dfrtp_1 _6133_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net413),
    .RESET_B(net180),
    .Q(\z80.tv80s.i_tv80_core.mcycles[5] ));
 sky130_fd_sc_hd__dfxtp_1 _6134_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(_0059_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6135_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(net416),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6136_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(_0061_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6137_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(net395),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6138_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(net322),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6139_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(net355),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6140_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(net332),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6141_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(net404),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6142_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(net384),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6143_ (.CLK(clknet_leaf_43_wb_clk_i),
    .D(net312),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6144_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(net316),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6145_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(_0070_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6146_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(net324),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6147_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(net402),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6148_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(net335),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6149_ (.CLK(clknet_leaf_43_wb_clk_i),
    .D(net342),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][7] ));
 sky130_fd_sc_hd__dfrtp_1 _6150_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0075_),
    .RESET_B(net183),
    .Q(\z80.tv80s.i_tv80_core.PreserveC_r ));
 sky130_fd_sc_hd__dfxtp_1 _6151_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(net330),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6152_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(net382),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6153_ (.CLK(clknet_leaf_43_wb_clk_i),
    .D(net314),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6154_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(net294),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6155_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(net398),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6156_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(net326),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6157_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(net337),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6158_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(net360),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][7] ));
 sky130_fd_sc_hd__dfstp_4 _6159_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net796),
    .SET_B(net179),
    .Q(\z80.tv80s.i_tv80_core.ISet[0] ));
 sky130_fd_sc_hd__dfrtp_1 _6160_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net568),
    .RESET_B(net179),
    .Q(\z80.tv80s.i_tv80_core.ISet[1] ));
 sky130_fd_sc_hd__dfrtp_1 _6161_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0002_),
    .RESET_B(net179),
    .Q(\z80.tv80s.i_tv80_core.ISet[2] ));
 sky130_fd_sc_hd__dfrtp_1 _6162_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net479),
    .RESET_B(net179),
    .Q(\z80.tv80s.i_tv80_core.ISet[3] ));
 sky130_fd_sc_hd__dfstp_1 _6163_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0020_),
    .SET_B(net171),
    .Q(net53));
 sky130_fd_sc_hd__dfstp_1 _6164_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0019_),
    .SET_B(net179),
    .Q(\z80.normal_rd_n ));
 sky130_fd_sc_hd__dfstp_1 _6165_ (.CLK(net218),
    .D(_0018_),
    .SET_B(net177),
    .Q(\z80.early_mreq_n ));
 sky130_fd_sc_hd__dfstp_1 _6166_ (.CLK(net219),
    .D(_0017_),
    .SET_B(net177),
    .Q(\z80.early_iorq_n ));
 sky130_fd_sc_hd__dfstp_1 _6167_ (.CLK(net220),
    .D(_0019_),
    .SET_B(net179),
    .Q(\z80.early_rd_n ));
 sky130_fd_sc_hd__dfstp_1 _6168_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0018_),
    .SET_B(net177),
    .Q(\z80.normal_mreq_n ));
 sky130_fd_sc_hd__dfstp_1 _6169_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0017_),
    .SET_B(net177),
    .Q(\z80.normal_iorq_n ));
 sky130_fd_sc_hd__dfxtp_1 _6170_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net286),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6171_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net284),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6172_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0086_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6173_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net339),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6174_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(_0088_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6175_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(_0089_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6176_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net318),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6177_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net481),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6178_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(net489),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6179_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(net357),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6180_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(_0094_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6181_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(_0095_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6182_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(net378),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6183_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(net408),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6184_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(net328),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6185_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(net366),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6186_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net276),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6187_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net420),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6188_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0102_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6189_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net302),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6190_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net432),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6191_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(_0105_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6192_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net274),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6193_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net436),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6194_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(_0108_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6195_ (.CLK(clknet_leaf_43_wb_clk_i),
    .D(net447),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6196_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(net362),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6197_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(net368),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6198_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(_0112_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6199_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(net411),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6200_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(_0114_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6201_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(net388),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6202_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net296),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6203_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net392),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6204_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net351),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6205_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net344),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6206_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(net418),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6207_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net320),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6208_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0122_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6209_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net476),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6210_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net347),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6211_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net380),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6212_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net445),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6213_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0127_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6214_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(_0128_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6215_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net288),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6216_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(net310),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6217_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0131_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6218_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(_0132_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6219_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(net439),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6220_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(_0134_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6221_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(_0135_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6222_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(_0136_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6223_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(_0137_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6224_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(net461),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6225_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(net463),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6226_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net370),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6227_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net513),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6228_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net493),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6229_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net422),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6230_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(_0144_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6231_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(_0145_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6232_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net449),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6233_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0147_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6234_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net278),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6235_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net304),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6236_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net290),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6237_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net372),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6238_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net306),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6239_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(net353),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6240_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net272),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6241_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net282),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][7] ));
 sky130_fd_sc_hd__dfrtp_1 _6242_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net256),
    .RESET_B(net180),
    .Q(\z80.tv80s.i_tv80_core.Pre_XY_F_M[1] ));
 sky130_fd_sc_hd__dfrtp_1 _6243_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net260),
    .RESET_B(net177),
    .Q(\z80.tv80s.i_tv80_core.Pre_XY_F_M[2] ));
 sky130_fd_sc_hd__dfrtp_1 _6244_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net500),
    .RESET_B(net178),
    .Q(\z80.tv80s.i_tv80_core.Pre_XY_F_M[3] ));
 sky130_fd_sc_hd__dfrtp_1 _6245_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net258),
    .RESET_B(net180),
    .Q(\z80.tv80s.i_tv80_core.Pre_XY_F_M[4] ));
 sky130_fd_sc_hd__dfrtp_1 _6246_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net400),
    .RESET_B(net180),
    .Q(\z80.tv80s.i_tv80_core.Pre_XY_F_M[5] ));
 sky130_fd_sc_hd__dfrtp_1 _6247_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net268),
    .RESET_B(net180),
    .Q(\z80.tv80s.i_tv80_core.Pre_XY_F_M[6] ));
 sky130_fd_sc_hd__dfrtp_1 _6248_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net522),
    .RESET_B(net180),
    .Q(\z80.tv80s.i_tv80_core.Pre_XY_F_M[7] ));
 sky130_fd_sc_hd__dfxtp_1 _6249_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net308),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6250_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net300),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6251_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0158_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6252_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0159_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6253_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(_0160_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6254_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(_0161_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6255_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net292),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6256_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net498),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][7] ));
 sky130_fd_sc_hd__dfrtp_1 _6257_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net586),
    .RESET_B(net181),
    .Q(\z80.tv80s.i_tv80_core.IStatus[1] ));
 sky130_fd_sc_hd__dfrtp_1 _6258_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net270),
    .RESET_B(net181),
    .Q(\z80.tv80s.i_tv80_core.IStatus[2] ));
 sky130_fd_sc_hd__dfxtp_1 _6259_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(net441),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6260_ (.CLK(clknet_leaf_43_wb_clk_i),
    .D(_0165_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6261_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_0166_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6262_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(net386),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6263_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(net425),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6264_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(_0169_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6265_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(net349),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6266_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(net374),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][7] ));
 sky130_fd_sc_hd__dfstp_1 _6267_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(net687),
    .SET_B(net182),
    .Q(\z80.tv80s.i_tv80_core.Ap[0] ));
 sky130_fd_sc_hd__dfstp_1 _6268_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(net657),
    .SET_B(net174),
    .Q(\z80.tv80s.i_tv80_core.Ap[1] ));
 sky130_fd_sc_hd__dfstp_1 _6269_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(net683),
    .SET_B(net182),
    .Q(\z80.tv80s.i_tv80_core.Ap[2] ));
 sky130_fd_sc_hd__dfstp_1 _6270_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(net697),
    .SET_B(net182),
    .Q(\z80.tv80s.i_tv80_core.Ap[3] ));
 sky130_fd_sc_hd__dfstp_1 _6271_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(net679),
    .SET_B(net174),
    .Q(\z80.tv80s.i_tv80_core.Ap[4] ));
 sky130_fd_sc_hd__dfstp_1 _6272_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(net675),
    .SET_B(net182),
    .Q(\z80.tv80s.i_tv80_core.Ap[5] ));
 sky130_fd_sc_hd__dfstp_1 _6273_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(net659),
    .SET_B(net182),
    .Q(\z80.tv80s.i_tv80_core.Ap[6] ));
 sky130_fd_sc_hd__dfstp_1 _6274_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(net655),
    .SET_B(net182),
    .Q(\z80.tv80s.i_tv80_core.Ap[7] ));
 sky130_fd_sc_hd__dfstp_1 _6275_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(net735),
    .SET_B(net183),
    .Q(\z80.tv80s.i_tv80_core.Fp[0] ));
 sky130_fd_sc_hd__dfstp_1 _6276_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(net748),
    .SET_B(net183),
    .Q(\z80.tv80s.i_tv80_core.Fp[1] ));
 sky130_fd_sc_hd__dfstp_1 _6277_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(net669),
    .SET_B(net182),
    .Q(\z80.tv80s.i_tv80_core.Fp[2] ));
 sky130_fd_sc_hd__dfstp_1 _6278_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(net731),
    .SET_B(net182),
    .Q(\z80.tv80s.i_tv80_core.Fp[3] ));
 sky130_fd_sc_hd__dfstp_1 _6279_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(net671),
    .SET_B(net183),
    .Q(\z80.tv80s.i_tv80_core.Fp[4] ));
 sky130_fd_sc_hd__dfstp_1 _6280_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(net706),
    .SET_B(net182),
    .Q(\z80.tv80s.i_tv80_core.Fp[5] ));
 sky130_fd_sc_hd__dfstp_1 _6281_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(net702),
    .SET_B(net182),
    .Q(\z80.tv80s.i_tv80_core.Fp[6] ));
 sky130_fd_sc_hd__dfstp_1 _6282_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(net667),
    .SET_B(net182),
    .Q(\z80.tv80s.i_tv80_core.Fp[7] ));
 sky130_fd_sc_hd__dfstp_4 _6283_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0033_),
    .SET_B(net179),
    .Q(net54));
 sky130_fd_sc_hd__dfxtp_4 _6284_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net673),
    .Q(\z80.tv80s.i_tv80_core.BusA[0] ));
 sky130_fd_sc_hd__dfxtp_4 _6285_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(net785),
    .Q(\z80.tv80s.i_tv80_core.BusA[1] ));
 sky130_fd_sc_hd__dfxtp_4 _6286_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net750),
    .Q(\z80.tv80s.i_tv80_core.BusA[2] ));
 sky130_fd_sc_hd__dfxtp_4 _6287_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(net691),
    .Q(\z80.tv80s.i_tv80_core.BusA[3] ));
 sky130_fd_sc_hd__dfxtp_4 _6288_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net708),
    .Q(\z80.tv80s.i_tv80_core.BusA[4] ));
 sky130_fd_sc_hd__dfxtp_4 _6289_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(net727),
    .Q(\z80.tv80s.i_tv80_core.BusA[5] ));
 sky130_fd_sc_hd__dfxtp_4 _6290_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net769),
    .Q(\z80.tv80s.i_tv80_core.BusA[6] ));
 sky130_fd_sc_hd__dfxtp_1 _6291_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net871),
    .Q(\z80.tv80s.i_tv80_core.BusA[7] ));
 sky130_fd_sc_hd__dfrtp_1 _6292_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net622),
    .RESET_B(net185),
    .Q(\z80.tv80s.i_tv80_core.NMI_s ));
 sky130_fd_sc_hd__dfrtp_1 _6293_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0197_),
    .RESET_B(net184),
    .Q(\z80.tv80s.i_tv80_core.IR[0] ));
 sky130_fd_sc_hd__dfrtp_1 _6294_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0198_),
    .RESET_B(net184),
    .Q(\z80.tv80s.i_tv80_core.IR[1] ));
 sky130_fd_sc_hd__dfrtp_1 _6295_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0199_),
    .RESET_B(net184),
    .Q(\z80.tv80s.i_tv80_core.IR[2] ));
 sky130_fd_sc_hd__dfrtp_1 _6296_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0200_),
    .RESET_B(net184),
    .Q(\z80.tv80s.i_tv80_core.IR[3] ));
 sky130_fd_sc_hd__dfrtp_2 _6297_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0201_),
    .RESET_B(net184),
    .Q(\z80.tv80s.i_tv80_core.IR[4] ));
 sky130_fd_sc_hd__dfrtp_1 _6298_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0202_),
    .RESET_B(net184),
    .Q(\z80.tv80s.i_tv80_core.IR[5] ));
 sky130_fd_sc_hd__dfrtp_4 _6299_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0203_),
    .RESET_B(net184),
    .Q(\z80.tv80s.i_tv80_core.IR[6] ));
 sky130_fd_sc_hd__dfrtp_4 _6300_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0204_),
    .RESET_B(net184),
    .Q(\z80.tv80s.i_tv80_core.IR[7] ));
 sky130_fd_sc_hd__dfrtp_1 _6301_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(net531),
    .RESET_B(net183),
    .Q(net48));
 sky130_fd_sc_hd__dfrtp_1 _6302_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net555),
    .RESET_B(net185),
    .Q(net47));
 sky130_fd_sc_hd__dfrtp_1 _6303_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net547),
    .RESET_B(net185),
    .Q(net45));
 sky130_fd_sc_hd__dfrtp_1 _6304_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(net537),
    .RESET_B(net183),
    .Q(net42));
 sky130_fd_sc_hd__dfrtp_1 _6305_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(net541),
    .RESET_B(net183),
    .Q(net41));
 sky130_fd_sc_hd__dfrtp_1 _6306_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(net539),
    .RESET_B(net183),
    .Q(net43));
 sky130_fd_sc_hd__dfrtp_1 _6307_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(net533),
    .RESET_B(net183),
    .Q(net44));
 sky130_fd_sc_hd__dfrtp_1 _6308_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net551),
    .RESET_B(net185),
    .Q(net46));
 sky130_fd_sc_hd__dfstp_4 _6309_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(net853),
    .SET_B(net182),
    .Q(\z80.tv80s.i_tv80_core.ACC[0] ));
 sky130_fd_sc_hd__dfstp_4 _6310_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0214_),
    .SET_B(net174),
    .Q(\z80.tv80s.i_tv80_core.ACC[1] ));
 sky130_fd_sc_hd__dfstp_4 _6311_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0215_),
    .SET_B(net182),
    .Q(\z80.tv80s.i_tv80_core.ACC[2] ));
 sky130_fd_sc_hd__dfstp_4 _6312_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0216_),
    .SET_B(net182),
    .Q(\z80.tv80s.i_tv80_core.ACC[3] ));
 sky130_fd_sc_hd__dfstp_4 _6313_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0217_),
    .SET_B(net174),
    .Q(\z80.tv80s.i_tv80_core.ACC[4] ));
 sky130_fd_sc_hd__dfstp_4 _6314_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0218_),
    .SET_B(net182),
    .Q(\z80.tv80s.i_tv80_core.ACC[5] ));
 sky130_fd_sc_hd__dfstp_4 _6315_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0219_),
    .SET_B(net174),
    .Q(\z80.tv80s.i_tv80_core.ACC[6] ));
 sky130_fd_sc_hd__dfstp_2 _6316_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0220_),
    .SET_B(net174),
    .Q(\z80.tv80s.i_tv80_core.ACC[7] ));
 sky130_fd_sc_hd__dfrtp_1 _6317_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(net570),
    .RESET_B(net173),
    .Q(net58));
 sky130_fd_sc_hd__dfrtp_1 _6318_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(net588),
    .RESET_B(net173),
    .Q(net28));
 sky130_fd_sc_hd__dfrtp_1 _6319_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(net561),
    .RESET_B(net170),
    .Q(net57));
 sky130_fd_sc_hd__dfrtp_1 _6320_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(net576),
    .RESET_B(net170),
    .Q(net56));
 sky130_fd_sc_hd__dfrtp_1 _6321_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(net592),
    .RESET_B(net170),
    .Q(net55));
 sky130_fd_sc_hd__dfrtp_1 _6322_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(net572),
    .RESET_B(net173),
    .Q(net29));
 sky130_fd_sc_hd__dfrtp_1 _6323_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(net602),
    .RESET_B(net173),
    .Q(net30));
 sky130_fd_sc_hd__dfrtp_1 _6324_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(net604),
    .RESET_B(net173),
    .Q(net31));
 sky130_fd_sc_hd__dfrtp_1 _6325_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(net636),
    .RESET_B(net170),
    .Q(net32));
 sky130_fd_sc_hd__dfrtp_1 _6326_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(net557),
    .RESET_B(net173),
    .Q(net33));
 sky130_fd_sc_hd__dfrtp_2 _6327_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(net608),
    .RESET_B(net171),
    .Q(net34));
 sky130_fd_sc_hd__dfrtp_2 _6328_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(net590),
    .RESET_B(net170),
    .Q(net35));
 sky130_fd_sc_hd__dfrtp_2 _6329_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(net632),
    .RESET_B(net170),
    .Q(net36));
 sky130_fd_sc_hd__dfrtp_2 _6330_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(net648),
    .RESET_B(net170),
    .Q(net37));
 sky130_fd_sc_hd__dfrtp_4 _6331_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(net725),
    .RESET_B(net171),
    .Q(net39));
 sky130_fd_sc_hd__dfrtp_2 _6332_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(net630),
    .RESET_B(net170),
    .Q(net40));
 sky130_fd_sc_hd__dfstp_4 _6333_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0237_),
    .SET_B(net183),
    .Q(\z80.tv80s.i_tv80_core.F[0] ));
 sky130_fd_sc_hd__dfstp_4 _6334_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0238_),
    .SET_B(net183),
    .Q(\z80.tv80s.i_tv80_core.F[1] ));
 sky130_fd_sc_hd__dfstp_4 _6335_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0239_),
    .SET_B(net182),
    .Q(\z80.tv80s.i_tv80_core.F[2] ));
 sky130_fd_sc_hd__dfstp_2 _6336_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0240_),
    .SET_B(net183),
    .Q(\z80.tv80s.i_tv80_core.F[3] ));
 sky130_fd_sc_hd__dfstp_2 _6337_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0241_),
    .SET_B(net183),
    .Q(\z80.tv80s.i_tv80_core.F[4] ));
 sky130_fd_sc_hd__dfstp_2 _6338_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0242_),
    .SET_B(net183),
    .Q(\z80.tv80s.i_tv80_core.F[5] ));
 sky130_fd_sc_hd__dfstp_2 _6339_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0243_),
    .SET_B(net185),
    .Q(\z80.tv80s.i_tv80_core.F[6] ));
 sky130_fd_sc_hd__dfstp_2 _6340_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(net834),
    .SET_B(net183),
    .Q(\z80.tv80s.i_tv80_core.F[7] ));
 sky130_fd_sc_hd__dfxtp_1 _6341_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(net430),
    .Q(\z80.tv80s.i_tv80_core.IncDecZ ));
 sky130_fd_sc_hd__dfrtp_1 _6342_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net451),
    .RESET_B(net184),
    .Q(\z80.tv80s.i_tv80_core.Z16_r ));
 sky130_fd_sc_hd__dfrtp_4 _6343_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0247_),
    .RESET_B(net184),
    .Q(\z80.tv80s.i_tv80_core.ALU_Op_r[0] ));
 sky130_fd_sc_hd__dfrtp_4 _6344_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(net826),
    .RESET_B(net184),
    .Q(\z80.tv80s.i_tv80_core.ALU_Op_r[1] ));
 sky130_fd_sc_hd__dfrtp_4 _6345_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0249_),
    .RESET_B(net184),
    .Q(\z80.tv80s.i_tv80_core.ALU_Op_r[2] ));
 sky130_fd_sc_hd__dfrtp_4 _6346_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0250_),
    .RESET_B(net184),
    .Q(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ));
 sky130_fd_sc_hd__dfrtp_4 _6347_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0251_),
    .RESET_B(net184),
    .Q(\z80.tv80s.i_tv80_core.Save_ALU_r ));
 sky130_fd_sc_hd__dfrtp_1 _6348_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net264),
    .RESET_B(net185),
    .Q(\z80.tv80s.i_tv80_core.BTR_r ));
 sky130_fd_sc_hd__dfrtp_1 _6349_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net634),
    .RESET_B(net176),
    .Q(\z80.tv80s.i_tv80_core.Read_To_Reg_r[0] ));
 sky130_fd_sc_hd__dfrtp_1 _6350_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net509),
    .RESET_B(net176),
    .Q(\z80.tv80s.i_tv80_core.Read_To_Reg_r[1] ));
 sky130_fd_sc_hd__dfrtp_1 _6351_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net502),
    .RESET_B(net179),
    .Q(\z80.tv80s.i_tv80_core.Read_To_Reg_r[2] ));
 sky130_fd_sc_hd__dfrtp_1 _6352_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(net465),
    .RESET_B(net179),
    .Q(\z80.tv80s.i_tv80_core.Read_To_Reg_r[3] ));
 sky130_fd_sc_hd__dfrtp_1 _6353_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net721),
    .RESET_B(net179),
    .Q(\z80.tv80s.i_tv80_core.Read_To_Reg_r[4] ));
 sky130_fd_sc_hd__dfrtp_1 _6354_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net626),
    .RESET_B(net184),
    .Q(\z80.tv80s.i_tv80_core.Arith16_r ));
 sky130_fd_sc_hd__dfxtp_2 _6355_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0259_),
    .Q(\z80.tv80s.i_tv80_core.RegAddrB_r[0] ));
 sky130_fd_sc_hd__dfxtp_1 _6356_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(net543),
    .Q(\z80.tv80s.i_tv80_core.RegAddrB_r[1] ));
 sky130_fd_sc_hd__dfrtp_1 _6357_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0261_),
    .RESET_B(net179),
    .Q(\z80.tv80s.i_tv80_core.XY_Ind ));
 sky130_fd_sc_hd__dfrtp_1 _6358_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net468),
    .RESET_B(net179),
    .Q(\z80.tv80s.i_tv80_core.XY_State[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6359_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0263_),
    .RESET_B(net179),
    .Q(\z80.tv80s.i_tv80_core.XY_State[1] ));
 sky130_fd_sc_hd__dfxtp_1 _6360_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0264_),
    .Q(\z80.tv80s.i_tv80_core.RegAddrC[0] ));
 sky130_fd_sc_hd__dfrtp_4 _6361_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(net802),
    .RESET_B(net175),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[0] ));
 sky130_fd_sc_hd__dfrtp_4 _6362_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(net791),
    .RESET_B(net181),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[1] ));
 sky130_fd_sc_hd__dfrtp_4 _6363_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(net804),
    .RESET_B(net175),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[2] ));
 sky130_fd_sc_hd__dfrtp_4 _6364_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(net828),
    .RESET_B(net181),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[3] ));
 sky130_fd_sc_hd__dfrtp_4 _6365_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(net816),
    .RESET_B(net181),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[4] ));
 sky130_fd_sc_hd__dfrtp_4 _6366_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(net822),
    .RESET_B(net181),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[5] ));
 sky130_fd_sc_hd__dfrtp_4 _6367_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(net811),
    .RESET_B(net175),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[6] ));
 sky130_fd_sc_hd__dfrtp_4 _6368_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(net813),
    .RESET_B(net181),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[7] ));
 sky130_fd_sc_hd__dfrtp_1 _6369_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(net594),
    .RESET_B(net172),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[8] ));
 sky130_fd_sc_hd__dfrtp_2 _6370_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(net612),
    .RESET_B(net172),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[9] ));
 sky130_fd_sc_hd__dfrtp_4 _6371_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(net762),
    .RESET_B(net172),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[10] ));
 sky130_fd_sc_hd__dfrtp_4 _6372_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(net777),
    .RESET_B(net172),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[11] ));
 sky130_fd_sc_hd__dfrtp_4 _6373_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(net754),
    .RESET_B(net172),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[12] ));
 sky130_fd_sc_hd__dfrtp_4 _6374_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(net783),
    .RESET_B(net172),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[13] ));
 sky130_fd_sc_hd__dfrtp_2 _6375_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(net752),
    .RESET_B(net172),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[14] ));
 sky130_fd_sc_hd__dfrtp_4 _6376_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(net760),
    .RESET_B(net172),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[15] ));
 sky130_fd_sc_hd__dfrtp_1 _6377_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net474),
    .RESET_B(net176),
    .Q(\z80.tv80s.i_tv80_core.Alternate ));
 sky130_fd_sc_hd__dfxtp_4 _6378_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(net710),
    .Q(\z80.tv80s.i_tv80_core.BusB[0] ));
 sky130_fd_sc_hd__dfxtp_4 _6379_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(net646),
    .Q(\z80.tv80s.i_tv80_core.BusB[1] ));
 sky130_fd_sc_hd__dfxtp_2 _6380_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(net775),
    .Q(\z80.tv80s.i_tv80_core.BusB[2] ));
 sky130_fd_sc_hd__dfxtp_4 _6381_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(net650),
    .Q(\z80.tv80s.i_tv80_core.BusB[3] ));
 sky130_fd_sc_hd__dfxtp_2 _6382_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(net729),
    .Q(\z80.tv80s.i_tv80_core.BusB[4] ));
 sky130_fd_sc_hd__dfxtp_4 _6383_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(net644),
    .Q(\z80.tv80s.i_tv80_core.BusB[5] ));
 sky130_fd_sc_hd__dfxtp_4 _6384_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(net620),
    .Q(\z80.tv80s.i_tv80_core.BusB[6] ));
 sky130_fd_sc_hd__dfxtp_4 _6385_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(net640),
    .Q(\z80.tv80s.i_tv80_core.BusB[7] ));
 sky130_fd_sc_hd__dfxtp_1 _6386_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0290_),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[0] ));
 sky130_fd_sc_hd__dfxtp_1 _6387_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0291_),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[1] ));
 sky130_fd_sc_hd__dfxtp_1 _6388_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net250),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[2] ));
 sky130_fd_sc_hd__dfxtp_1 _6389_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net254),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[3] ));
 sky130_fd_sc_hd__dfxtp_1 _6390_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(net224),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[4] ));
 sky130_fd_sc_hd__dfxtp_1 _6391_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(net248),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[5] ));
 sky130_fd_sc_hd__dfxtp_1 _6392_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net252),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[6] ));
 sky130_fd_sc_hd__dfxtp_1 _6393_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(net234),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[7] ));
 sky130_fd_sc_hd__dfxtp_1 _6394_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(net230),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[8] ));
 sky130_fd_sc_hd__dfxtp_1 _6395_ (.CLK(clknet_leaf_43_wb_clk_i),
    .D(net244),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[9] ));
 sky130_fd_sc_hd__dfxtp_1 _6396_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(net238),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[10] ));
 sky130_fd_sc_hd__dfxtp_1 _6397_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net236),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[11] ));
 sky130_fd_sc_hd__dfxtp_1 _6398_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(net246),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[12] ));
 sky130_fd_sc_hd__dfxtp_1 _6399_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(net242),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[13] ));
 sky130_fd_sc_hd__dfxtp_1 _6400_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(net228),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[14] ));
 sky130_fd_sc_hd__dfxtp_1 _6401_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(net232),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[15] ));
 sky130_fd_sc_hd__dfrtp_1 _6402_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(net582),
    .RESET_B(net170),
    .Q(\z80.tv80s.i_tv80_core.I[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6403_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(net677),
    .RESET_B(net170),
    .Q(\z80.tv80s.i_tv80_core.I[1] ));
 sky130_fd_sc_hd__dfrtp_2 _6404_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(net624),
    .RESET_B(net170),
    .Q(\z80.tv80s.i_tv80_core.I[2] ));
 sky130_fd_sc_hd__dfrtp_2 _6405_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(net628),
    .RESET_B(net170),
    .Q(\z80.tv80s.i_tv80_core.I[3] ));
 sky130_fd_sc_hd__dfrtp_1 _6406_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(net580),
    .RESET_B(net171),
    .Q(\z80.tv80s.i_tv80_core.I[4] ));
 sky130_fd_sc_hd__dfrtp_2 _6407_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(net723),
    .RESET_B(net170),
    .Q(\z80.tv80s.i_tv80_core.I[5] ));
 sky130_fd_sc_hd__dfrtp_2 _6408_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(net733),
    .RESET_B(net171),
    .Q(\z80.tv80s.i_tv80_core.I[6] ));
 sky130_fd_sc_hd__dfrtp_4 _6409_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(net793),
    .RESET_B(net170),
    .Q(\z80.tv80s.i_tv80_core.I[7] ));
 sky130_fd_sc_hd__dfrtp_1 _6410_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(net495),
    .RESET_B(net173),
    .Q(\z80.tv80s.i_tv80_core.R[7] ));
 sky130_fd_sc_hd__dfxtp_1 _6411_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net262),
    .Q(\z80.tv80s.i_tv80_core.RegAddrA_r[0] ));
 sky130_fd_sc_hd__dfxtp_1 _6412_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net240),
    .Q(\z80.tv80s.i_tv80_core.RegAddrA_r[1] ));
 sky130_fd_sc_hd__dfrtp_1 _6413_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(net642),
    .RESET_B(net174),
    .Q(\z80.tv80s.i_tv80_core.PC[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6414_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(net695),
    .RESET_B(net174),
    .Q(\z80.tv80s.i_tv80_core.PC[1] ));
 sky130_fd_sc_hd__dfrtp_2 _6415_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(net618),
    .RESET_B(net174),
    .Q(\z80.tv80s.i_tv80_core.PC[2] ));
 sky130_fd_sc_hd__dfrtp_2 _6416_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(net596),
    .RESET_B(net173),
    .Q(\z80.tv80s.i_tv80_core.PC[3] ));
 sky130_fd_sc_hd__dfrtp_2 _6417_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(net600),
    .RESET_B(net173),
    .Q(\z80.tv80s.i_tv80_core.PC[4] ));
 sky130_fd_sc_hd__dfrtp_2 _6418_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(net578),
    .RESET_B(net173),
    .Q(\z80.tv80s.i_tv80_core.PC[5] ));
 sky130_fd_sc_hd__dfrtp_4 _6419_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(net745),
    .RESET_B(net173),
    .Q(\z80.tv80s.i_tv80_core.PC[6] ));
 sky130_fd_sc_hd__dfrtp_4 _6420_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(net739),
    .RESET_B(net170),
    .Q(\z80.tv80s.i_tv80_core.PC[7] ));
 sky130_fd_sc_hd__dfrtp_4 _6421_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(net809),
    .RESET_B(net171),
    .Q(\z80.tv80s.i_tv80_core.PC[8] ));
 sky130_fd_sc_hd__dfrtp_4 _6422_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(net789),
    .RESET_B(net170),
    .Q(\z80.tv80s.i_tv80_core.PC[9] ));
 sky130_fd_sc_hd__dfrtp_4 _6423_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(net807),
    .RESET_B(net171),
    .Q(\z80.tv80s.i_tv80_core.PC[10] ));
 sky130_fd_sc_hd__dfrtp_4 _6424_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(net800),
    .RESET_B(net171),
    .Q(\z80.tv80s.i_tv80_core.PC[11] ));
 sky130_fd_sc_hd__dfrtp_4 _6425_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(net773),
    .RESET_B(net171),
    .Q(\z80.tv80s.i_tv80_core.PC[12] ));
 sky130_fd_sc_hd__dfrtp_4 _6426_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(net781),
    .RESET_B(net171),
    .Q(\z80.tv80s.i_tv80_core.PC[13] ));
 sky130_fd_sc_hd__dfrtp_4 _6427_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(net767),
    .RESET_B(net172),
    .Q(\z80.tv80s.i_tv80_core.PC[14] ));
 sky130_fd_sc_hd__dfrtp_2 _6428_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(net758),
    .RESET_B(net172),
    .Q(\z80.tv80s.i_tv80_core.PC[15] ));
 sky130_fd_sc_hd__dfstp_1 _6429_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0333_),
    .SET_B(net178),
    .Q(\z80.tv80s.i_tv80_core.i_mcode.MCycle[0] ));
 sky130_fd_sc_hd__dfrtp_4 _6430_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net717),
    .RESET_B(net178),
    .Q(\z80.tv80s.i_tv80_core.i_mcode.MCycle[1] ));
 sky130_fd_sc_hd__dfrtp_4 _6431_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net787),
    .RESET_B(net178),
    .Q(\z80.tv80s.i_tv80_core.i_mcode.MCycle[2] ));
 sky130_fd_sc_hd__dfrtp_4 _6432_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net693),
    .RESET_B(net178),
    .Q(\z80.tv80s.i_tv80_core.i_mcode.MCycle[3] ));
 sky130_fd_sc_hd__dfrtp_1 _6433_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0337_),
    .RESET_B(net178),
    .Q(\z80.tv80s.i_tv80_core.i_mcode.MCycle[4] ));
 sky130_fd_sc_hd__dfrtp_4 _6434_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0338_),
    .RESET_B(net178),
    .Q(\z80.tv80s.i_tv80_core.i_mcode.MCycle[5] ));
 sky130_fd_sc_hd__dfrtp_4 _6435_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net700),
    .RESET_B(net177),
    .Q(\z80.tv80s.i_tv80_core.i_mcode.MCycle[6] ));
 sky130_fd_sc_hd__dfrtp_4 _6436_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net712),
    .RESET_B(net178),
    .Q(\z80.tv80s.i_tv80_core.Halt_FF ));
 sky130_fd_sc_hd__dfrtp_1 _6437_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net653),
    .RESET_B(net178),
    .Q(_0034_));
 sky130_fd_sc_hd__dfrtp_1 _6438_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net610),
    .RESET_B(net178),
    .Q(_0035_));
 sky130_fd_sc_hd__dfrtp_1 _6439_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0031_),
    .RESET_B(net178),
    .Q(_0036_));
 sky130_fd_sc_hd__dfrtp_1 _6440_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0021_),
    .RESET_B(net177),
    .Q(\z80.tv80s.i_tv80_core.Auto_Wait_t1 ));
 sky130_fd_sc_hd__dfrtp_1 _6441_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0028_),
    .RESET_B(net185),
    .Q(\z80.tv80s.i_tv80_core.No_BTR ));
 sky130_fd_sc_hd__dfrtp_4 _6442_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net779),
    .RESET_B(net181),
    .Q(\z80.tv80s.i_tv80_core.IntCycle ));
 sky130_fd_sc_hd__dfrtp_1 _6443_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0022_),
    .RESET_B(net177),
    .Q(\z80.tv80s.i_tv80_core.Auto_Wait_t2 ));
 sky130_fd_sc_hd__dfrtp_1 _6444_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net222),
    .RESET_B(net178),
    .Q(\z80.tv80s.i_tv80_core.BusAck ));
 sky130_fd_sc_hd__dfrtp_1 _6445_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(net14),
    .RESET_B(net184),
    .Q(\z80.tv80s.i_tv80_core.Oldnmi_n ));
 sky130_fd_sc_hd__dfrtp_1 _6446_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0025_),
    .RESET_B(net185),
    .Q(\z80.tv80s.i_tv80_core.INT_s ));
 sky130_fd_sc_hd__dfrtp_2 _6447_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net519),
    .RESET_B(net179),
    .Q(\z80.tv80s.i_tv80_core.NMICycle ));
 sky130_fd_sc_hd__dfrtp_1 _6448_ (.CLK(clknet_2_3__leaf_wb_clk_i),
    .D(_0023_),
    .RESET_B(net185),
    .Q(\z80.tv80s.i_tv80_core.BusReq_s ));
 sky130_fd_sc_hd__dfxtp_1 _6449_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net471),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6450_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net487),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6451_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net515),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6452_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net376),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6453_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(_0347_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6454_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(_0348_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6455_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net390),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6456_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0350_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][7] ));
 sky130_fd_sc_hd__dfstp_2 _6457_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net606),
    .SET_B(net179),
    .Q(net38));
 sky130_fd_sc_hd__dfrtp_4 _6458_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0351_),
    .RESET_B(net181),
    .Q(\z80.tv80s.di_reg[0] ));
 sky130_fd_sc_hd__dfrtp_4 _6459_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0352_),
    .RESET_B(net181),
    .Q(\z80.tv80s.di_reg[1] ));
 sky130_fd_sc_hd__dfrtp_4 _6460_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0353_),
    .RESET_B(net181),
    .Q(\z80.tv80s.di_reg[2] ));
 sky130_fd_sc_hd__dfrtp_4 _6461_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0354_),
    .RESET_B(net181),
    .Q(\z80.tv80s.di_reg[3] ));
 sky130_fd_sc_hd__dfrtp_4 _6462_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0355_),
    .RESET_B(net181),
    .Q(\z80.tv80s.di_reg[4] ));
 sky130_fd_sc_hd__dfrtp_4 _6463_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0356_),
    .RESET_B(net181),
    .Q(\z80.tv80s.di_reg[5] ));
 sky130_fd_sc_hd__dfrtp_4 _6464_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0357_),
    .RESET_B(net181),
    .Q(\z80.tv80s.di_reg[6] ));
 sky130_fd_sc_hd__dfrtp_4 _6465_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0358_),
    .RESET_B(net181),
    .Q(\z80.tv80s.di_reg[7] ));
 sky130_fd_sc_hd__dfstp_1 _6466_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net266),
    .SET_B(net177),
    .Q(\z80.tv80s.i_tv80_core.ts[0] ));
 sky130_fd_sc_hd__dfrtp_1 _6467_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0360_),
    .RESET_B(net177),
    .Q(\z80.tv80s.i_tv80_core.ts[1] ));
 sky130_fd_sc_hd__dfrtp_4 _6468_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net574),
    .RESET_B(net177),
    .Q(\z80.tv80s.i_tv80_core.ts[2] ));
 sky130_fd_sc_hd__dfrtp_4 _6469_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0362_),
    .RESET_B(net177),
    .Q(\z80.tv80s.i_tv80_core.ts[3] ));
 sky130_fd_sc_hd__dfrtp_1 _6470_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net737),
    .RESET_B(net177),
    .Q(\z80.tv80s.i_tv80_core.ts[4] ));
 sky130_fd_sc_hd__dfrtp_1 _6471_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net364),
    .RESET_B(net177),
    .Q(\z80.tv80s.i_tv80_core.ts[5] ));
 sky130_fd_sc_hd__dfrtp_1 _6472_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net298),
    .RESET_B(net177),
    .Q(\z80.tv80s.i_tv80_core.ts[6] ));
 sky130_fd_sc_hd__dfrtp_1 _6473_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net765),
    .RESET_B(net179),
    .Q(\z80.tv80s.i_tv80_core.IntE ));
 sky130_fd_sc_hd__dfrtp_1 _6474_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net843),
    .RESET_B(net180),
    .Q(\z80.tv80s.i_tv80_core.IntE_FF2 ));
 sky130_fd_sc_hd__dfstp_1 _6475_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(net638),
    .SET_B(net175),
    .Q(\z80.tv80s.i_tv80_core.SP[0] ));
 sky130_fd_sc_hd__dfstp_1 _6476_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(net681),
    .SET_B(net176),
    .Q(\z80.tv80s.i_tv80_core.SP[1] ));
 sky130_fd_sc_hd__dfstp_1 _6477_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(net714),
    .SET_B(net176),
    .Q(\z80.tv80s.i_tv80_core.SP[2] ));
 sky130_fd_sc_hd__dfstp_1 _6478_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(net704),
    .SET_B(net176),
    .Q(\z80.tv80s.i_tv80_core.SP[3] ));
 sky130_fd_sc_hd__dfstp_1 _6479_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(net663),
    .SET_B(net176),
    .Q(\z80.tv80s.i_tv80_core.SP[4] ));
 sky130_fd_sc_hd__dfstp_1 _6480_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(net719),
    .SET_B(net175),
    .Q(\z80.tv80s.i_tv80_core.SP[5] ));
 sky130_fd_sc_hd__dfstp_1 _6481_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(net661),
    .SET_B(net176),
    .Q(\z80.tv80s.i_tv80_core.SP[6] ));
 sky130_fd_sc_hd__dfstp_1 _6482_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(_0373_),
    .SET_B(net176),
    .Q(\z80.tv80s.i_tv80_core.SP[7] ));
 sky130_fd_sc_hd__dfstp_1 _6483_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(net665),
    .SET_B(net176),
    .Q(\z80.tv80s.i_tv80_core.SP[8] ));
 sky130_fd_sc_hd__dfstp_1 _6484_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(net741),
    .SET_B(net172),
    .Q(\z80.tv80s.i_tv80_core.SP[9] ));
 sky130_fd_sc_hd__dfstp_1 _6485_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(net584),
    .SET_B(net172),
    .Q(\z80.tv80s.i_tv80_core.SP[10] ));
 sky130_fd_sc_hd__dfstp_1 _6486_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(net743),
    .SET_B(net172),
    .Q(\z80.tv80s.i_tv80_core.SP[11] ));
 sky130_fd_sc_hd__dfstp_2 _6487_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(net756),
    .SET_B(net176),
    .Q(\z80.tv80s.i_tv80_core.SP[12] ));
 sky130_fd_sc_hd__dfstp_1 _6488_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(net689),
    .SET_B(net172),
    .Q(\z80.tv80s.i_tv80_core.SP[13] ));
 sky130_fd_sc_hd__dfstp_2 _6489_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(_0380_),
    .SET_B(net176),
    .Q(\z80.tv80s.i_tv80_core.SP[14] ));
 sky130_fd_sc_hd__dfstp_1 _6490_ (.CLK(clknet_leaf_43_wb_clk_i),
    .D(_0381_),
    .SET_B(net176),
    .Q(\z80.tv80s.i_tv80_core.SP[15] ));
 sky130_fd_sc_hd__buf_1 _6523_ (.A(net26),
    .X(net19));
 sky130_fd_sc_hd__buf_1 _6524_ (.A(net26),
    .X(net20));
 sky130_fd_sc_hd__buf_1 _6525_ (.A(net26),
    .X(net21));
 sky130_fd_sc_hd__buf_1 _6526_ (.A(net26),
    .X(net22));
 sky130_fd_sc_hd__buf_1 _6527_ (.A(net26),
    .X(net23));
 sky130_fd_sc_hd__buf_1 _6528_ (.A(net26),
    .X(net24));
 sky130_fd_sc_hd__buf_1 _6529_ (.A(net26),
    .X(net25));
 sky130_fd_sc_hd__conb_1 ci2406_z80_186 (.LO(net186));
 sky130_fd_sc_hd__conb_1 ci2406_z80_187 (.LO(net187));
 sky130_fd_sc_hd__conb_1 ci2406_z80_188 (.LO(net188));
 sky130_fd_sc_hd__conb_1 ci2406_z80_189 (.LO(net189));
 sky130_fd_sc_hd__conb_1 ci2406_z80_190 (.LO(net190));
 sky130_fd_sc_hd__conb_1 ci2406_z80_191 (.LO(net191));
 sky130_fd_sc_hd__conb_1 ci2406_z80_192 (.LO(net192));
 sky130_fd_sc_hd__conb_1 ci2406_z80_193 (.LO(net193));
 sky130_fd_sc_hd__conb_1 ci2406_z80_194 (.LO(net194));
 sky130_fd_sc_hd__conb_1 ci2406_z80_195 (.LO(net195));
 sky130_fd_sc_hd__conb_1 ci2406_z80_196 (.LO(net196));
 sky130_fd_sc_hd__conb_1 ci2406_z80_197 (.LO(net197));
 sky130_fd_sc_hd__conb_1 ci2406_z80_198 (.LO(net198));
 sky130_fd_sc_hd__conb_1 ci2406_z80_199 (.LO(net199));
 sky130_fd_sc_hd__conb_1 ci2406_z80_200 (.LO(net200));
 sky130_fd_sc_hd__conb_1 ci2406_z80_201 (.LO(net201));
 sky130_fd_sc_hd__conb_1 ci2406_z80_202 (.LO(net202));
 sky130_fd_sc_hd__conb_1 ci2406_z80_203 (.LO(net203));
 sky130_fd_sc_hd__conb_1 ci2406_z80_204 (.LO(net204));
 sky130_fd_sc_hd__conb_1 ci2406_z80_205 (.LO(net205));
 sky130_fd_sc_hd__conb_1 ci2406_z80_206 (.LO(net206));
 sky130_fd_sc_hd__conb_1 ci2406_z80_207 (.LO(net207));
 sky130_fd_sc_hd__conb_1 ci2406_z80_208 (.LO(net208));
 sky130_fd_sc_hd__conb_1 ci2406_z80_209 (.LO(net209));
 sky130_fd_sc_hd__conb_1 ci2406_z80_210 (.LO(net210));
 sky130_fd_sc_hd__conb_1 ci2406_z80_211 (.LO(net211));
 sky130_fd_sc_hd__conb_1 ci2406_z80_212 (.LO(net212));
 sky130_fd_sc_hd__conb_1 ci2406_z80_213 (.LO(net213));
 sky130_fd_sc_hd__conb_1 ci2406_z80_214 (.HI(net214));
 sky130_fd_sc_hd__conb_1 ci2406_z80_215 (.HI(net215));
 sky130_fd_sc_hd__conb_1 ci2406_z80_216 (.HI(net216));
 sky130_fd_sc_hd__conb_1 ci2406_z80_217 (.HI(net217));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_wb_clk_i (.A(wb_clk_i),
    .X(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_13_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_15_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_18_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_21_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_23_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_24_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_25_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_26_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_wb_clk_i (.A(clknet_2_2__leaf_wb_clk_i),
    .X(clknet_leaf_27_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_wb_clk_i (.A(clknet_2_2__leaf_wb_clk_i),
    .X(clknet_leaf_28_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_wb_clk_i (.A(clknet_2_2__leaf_wb_clk_i),
    .X(clknet_leaf_29_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_wb_clk_i (.A(clknet_2_2__leaf_wb_clk_i),
    .X(clknet_leaf_30_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_wb_clk_i (.A(clknet_2_2__leaf_wb_clk_i),
    .X(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_wb_clk_i (.A(clknet_2_2__leaf_wb_clk_i),
    .X(clknet_leaf_32_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_wb_clk_i (.A(clknet_2_2__leaf_wb_clk_i),
    .X(clknet_leaf_33_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_wb_clk_i (.A(clknet_2_2__leaf_wb_clk_i),
    .X(clknet_leaf_34_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_wb_clk_i (.A(clknet_2_2__leaf_wb_clk_i),
    .X(clknet_leaf_35_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_36_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_37_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_38_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_39_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_40_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_41_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_42_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_43_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_44_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_45_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_46_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_47_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_48_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_49_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_50_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_9_wb_clk_i));
 sky130_fd_sc_hd__buf_4 fanout100 (.A(net101),
    .X(net100));
 sky130_fd_sc_hd__buf_6 fanout101 (.A(_0598_),
    .X(net101));
 sky130_fd_sc_hd__buf_4 fanout102 (.A(_0598_),
    .X(net102));
 sky130_fd_sc_hd__buf_6 fanout103 (.A(_0501_),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_4 fanout104 (.A(_0501_),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_8 fanout105 (.A(_0388_),
    .X(net105));
 sky130_fd_sc_hd__buf_6 fanout106 (.A(_0387_),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_4 fanout107 (.A(_0387_),
    .X(net107));
 sky130_fd_sc_hd__buf_4 fanout108 (.A(_2981_),
    .X(net108));
 sky130_fd_sc_hd__buf_4 fanout109 (.A(_2980_),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_8 fanout110 (.A(_2886_),
    .X(net110));
 sky130_fd_sc_hd__buf_4 fanout111 (.A(_2864_),
    .X(net111));
 sky130_fd_sc_hd__buf_6 fanout112 (.A(net27),
    .X(net112));
 sky130_fd_sc_hd__clkbuf_8 fanout113 (.A(net27),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_4 fanout114 (.A(net27),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_8 fanout115 (.A(net116),
    .X(net115));
 sky130_fd_sc_hd__buf_4 fanout116 (.A(net117),
    .X(net116));
 sky130_fd_sc_hd__buf_4 fanout117 (.A(net27),
    .X(net117));
 sky130_fd_sc_hd__clkbuf_8 fanout118 (.A(net119),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_8 fanout119 (.A(_2850_),
    .X(net119));
 sky130_fd_sc_hd__buf_4 fanout120 (.A(_2845_),
    .X(net120));
 sky130_fd_sc_hd__buf_6 fanout121 (.A(net122),
    .X(net121));
 sky130_fd_sc_hd__buf_8 fanout122 (.A(net736),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_8 fanout123 (.A(net124),
    .X(net123));
 sky130_fd_sc_hd__buf_6 fanout124 (.A(net746),
    .X(net124));
 sky130_fd_sc_hd__buf_4 fanout125 (.A(net127),
    .X(net125));
 sky130_fd_sc_hd__buf_2 fanout126 (.A(net127),
    .X(net126));
 sky130_fd_sc_hd__buf_4 fanout127 (.A(net128),
    .X(net127));
 sky130_fd_sc_hd__buf_4 fanout128 (.A(net746),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_8 fanout129 (.A(net651),
    .X(net129));
 sky130_fd_sc_hd__buf_6 fanout130 (.A(net786),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_8 fanout131 (.A(net132),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_8 fanout132 (.A(\z80.tv80s.i_tv80_core.i_mcode.MCycle[1] ),
    .X(net132));
 sky130_fd_sc_hd__buf_4 fanout133 (.A(net134),
    .X(net133));
 sky130_fd_sc_hd__buf_4 fanout134 (.A(net137),
    .X(net134));
 sky130_fd_sc_hd__buf_4 fanout135 (.A(net137),
    .X(net135));
 sky130_fd_sc_hd__buf_6 fanout136 (.A(net137),
    .X(net136));
 sky130_fd_sc_hd__clkbuf_8 fanout137 (.A(net858),
    .X(net137));
 sky130_fd_sc_hd__buf_6 fanout138 (.A(net139),
    .X(net138));
 sky130_fd_sc_hd__buf_8 fanout139 (.A(net864),
    .X(net139));
 sky130_fd_sc_hd__buf_6 fanout140 (.A(net534),
    .X(net140));
 sky130_fd_sc_hd__buf_4 fanout141 (.A(net142),
    .X(net141));
 sky130_fd_sc_hd__clkbuf_8 fanout142 (.A(net872),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_8 fanout143 (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[1] ),
    .X(net143));
 sky130_fd_sc_hd__clkbuf_8 fanout144 (.A(net145),
    .X(net144));
 sky130_fd_sc_hd__buf_4 fanout145 (.A(net146),
    .X(net145));
 sky130_fd_sc_hd__buf_4 fanout146 (.A(net794),
    .X(net146));
 sky130_fd_sc_hd__buf_4 fanout147 (.A(net868),
    .X(net147));
 sky130_fd_sc_hd__buf_4 fanout148 (.A(net149),
    .X(net148));
 sky130_fd_sc_hd__buf_4 fanout149 (.A(\z80.tv80s.i_tv80_core.IR[4] ),
    .X(net149));
 sky130_fd_sc_hd__buf_4 fanout150 (.A(net152),
    .X(net150));
 sky130_fd_sc_hd__buf_2 fanout151 (.A(net152),
    .X(net151));
 sky130_fd_sc_hd__buf_4 fanout152 (.A(net876),
    .X(net152));
 sky130_fd_sc_hd__buf_4 fanout153 (.A(net154),
    .X(net153));
 sky130_fd_sc_hd__buf_4 fanout154 (.A(net867),
    .X(net154));
 sky130_fd_sc_hd__buf_4 fanout155 (.A(net157),
    .X(net155));
 sky130_fd_sc_hd__clkbuf_2 fanout156 (.A(net157),
    .X(net156));
 sky130_fd_sc_hd__clkbuf_4 fanout157 (.A(net866),
    .X(net157));
 sky130_fd_sc_hd__buf_4 fanout158 (.A(net159),
    .X(net158));
 sky130_fd_sc_hd__buf_4 fanout159 (.A(net831),
    .X(net159));
 sky130_fd_sc_hd__buf_4 fanout160 (.A(net161),
    .X(net160));
 sky130_fd_sc_hd__buf_4 fanout161 (.A(net869),
    .X(net161));
 sky130_fd_sc_hd__buf_4 fanout162 (.A(net870),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_8 fanout163 (.A(net824),
    .X(net163));
 sky130_fd_sc_hd__buf_4 fanout164 (.A(net166),
    .X(net164));
 sky130_fd_sc_hd__clkbuf_8 fanout165 (.A(net166),
    .X(net165));
 sky130_fd_sc_hd__clkbuf_8 fanout166 (.A(\z80.tv80s.i_tv80_core.ISet[0] ),
    .X(net166));
 sky130_fd_sc_hd__clkbuf_8 fanout167 (.A(net168),
    .X(net167));
 sky130_fd_sc_hd__buf_6 fanout168 (.A(net861),
    .X(net168));
 sky130_fd_sc_hd__buf_8 fanout169 (.A(\z80.tv80s.i_tv80_core.RegAddrC[2] ),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_8 fanout170 (.A(net171),
    .X(net170));
 sky130_fd_sc_hd__buf_4 fanout171 (.A(net172),
    .X(net171));
 sky130_fd_sc_hd__clkbuf_8 fanout172 (.A(net175),
    .X(net172));
 sky130_fd_sc_hd__clkbuf_8 fanout173 (.A(net175),
    .X(net173));
 sky130_fd_sc_hd__buf_4 fanout174 (.A(net175),
    .X(net174));
 sky130_fd_sc_hd__buf_4 fanout175 (.A(net176),
    .X(net175));
 sky130_fd_sc_hd__buf_4 fanout176 (.A(net18),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_8 fanout177 (.A(net180),
    .X(net177));
 sky130_fd_sc_hd__buf_4 fanout178 (.A(net180),
    .X(net178));
 sky130_fd_sc_hd__clkbuf_8 fanout179 (.A(net180),
    .X(net179));
 sky130_fd_sc_hd__buf_4 fanout180 (.A(net18),
    .X(net180));
 sky130_fd_sc_hd__clkbuf_8 fanout181 (.A(net185),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_8 fanout182 (.A(net183),
    .X(net182));
 sky130_fd_sc_hd__clkbuf_8 fanout183 (.A(net185),
    .X(net183));
 sky130_fd_sc_hd__clkbuf_8 fanout184 (.A(net185),
    .X(net184));
 sky130_fd_sc_hd__clkbuf_8 fanout185 (.A(net18),
    .X(net185));
 sky130_fd_sc_hd__clkbuf_8 fanout59 (.A(_1666_),
    .X(net59));
 sky130_fd_sc_hd__buf_8 fanout60 (.A(_0576_),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_8 fanout61 (.A(_0498_),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_8 fanout63 (.A(_2570_),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_8 fanout64 (.A(_2581_),
    .X(net64));
 sky130_fd_sc_hd__buf_4 fanout65 (.A(net66),
    .X(net65));
 sky130_fd_sc_hd__buf_2 fanout66 (.A(_1683_),
    .X(net66));
 sky130_fd_sc_hd__buf_4 fanout67 (.A(net68),
    .X(net67));
 sky130_fd_sc_hd__buf_4 fanout68 (.A(_1681_),
    .X(net68));
 sky130_fd_sc_hd__buf_4 fanout69 (.A(_0805_),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_8 fanout70 (.A(_0804_),
    .X(net70));
 sky130_fd_sc_hd__buf_4 fanout72 (.A(_2346_),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_8 fanout73 (.A(_0984_),
    .X(net73));
 sky130_fd_sc_hd__buf_6 fanout74 (.A(net75),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_8 fanout75 (.A(_0983_),
    .X(net75));
 sky130_fd_sc_hd__buf_4 fanout76 (.A(_0809_),
    .X(net76));
 sky130_fd_sc_hd__buf_4 fanout77 (.A(_2671_),
    .X(net77));
 sky130_fd_sc_hd__buf_4 fanout78 (.A(_1670_),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_8 fanout79 (.A(_1669_),
    .X(net79));
 sky130_fd_sc_hd__buf_4 fanout80 (.A(_0866_),
    .X(net80));
 sky130_fd_sc_hd__buf_2 fanout81 (.A(_0866_),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_8 fanout82 (.A(_0981_),
    .X(net82));
 sky130_fd_sc_hd__buf_4 fanout83 (.A(_0981_),
    .X(net83));
 sky130_fd_sc_hd__buf_4 fanout84 (.A(_0981_),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_8 fanout85 (.A(_0775_),
    .X(net85));
 sky130_fd_sc_hd__buf_6 fanout86 (.A(_0773_),
    .X(net86));
 sky130_fd_sc_hd__buf_4 fanout87 (.A(net88),
    .X(net87));
 sky130_fd_sc_hd__buf_4 fanout88 (.A(_1418_),
    .X(net88));
 sky130_fd_sc_hd__buf_6 fanout89 (.A(_0772_),
    .X(net89));
 sky130_fd_sc_hd__buf_4 fanout90 (.A(_1417_),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_8 fanout93 (.A(net95),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_8 fanout94 (.A(net95),
    .X(net94));
 sky130_fd_sc_hd__buf_4 fanout95 (.A(_0599_),
    .X(net95));
 sky130_fd_sc_hd__buf_4 fanout96 (.A(_2995_),
    .X(net96));
 sky130_fd_sc_hd__buf_4 fanout97 (.A(_2983_),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_8 fanout98 (.A(net99),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_8 fanout99 (.A(_1685_),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_2 hold1 (.A(\z80.tv80s.i_tv80_core.BusReq_s ),
    .X(net221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(_0298_),
    .X(net230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(_0121_),
    .X(net320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][4] ),
    .X(net321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(_0063_),
    .X(net322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][4] ),
    .X(net323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(_0071_),
    .X(net324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][5] ),
    .X(net325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(_0081_),
    .X(net326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][6] ),
    .X(net327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(_0098_),
    .X(net328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][0] ),
    .X(net329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\z80.tv80s.i_tv80_core.RegBusA_r[15] ),
    .X(net231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(_0076_),
    .X(net330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][6] ),
    .X(net331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(_0065_),
    .X(net332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][6] ),
    .X(net333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][6] ),
    .X(net334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(_0073_),
    .X(net335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][6] ),
    .X(net336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(_0082_),
    .X(net337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][3] ),
    .X(net338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(_0087_),
    .X(net339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(_0305_),
    .X(net232));
 sky130_fd_sc_hd__buf_1 hold120 (.A(net879),
    .X(net340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][7] ),
    .X(net341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(_0074_),
    .X(net342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][3] ),
    .X(net343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(_0119_),
    .X(net344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][2] ),
    .X(net345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][0] ),
    .X(net346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(_0124_),
    .X(net347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][6] ),
    .X(net348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(_0170_),
    .X(net349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\z80.tv80s.i_tv80_core.RegBusA_r[7] ),
    .X(net233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][2] ),
    .X(net350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(_0118_),
    .X(net351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][5] ),
    .X(net352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(_0153_),
    .X(net353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][5] ),
    .X(net354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(_0064_),
    .X(net355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][1] ),
    .X(net356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(_0093_),
    .X(net357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][6] ),
    .X(net358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][7] ),
    .X(net359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(_0297_),
    .X(net234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(_0083_),
    .X(net360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][2] ),
    .X(net361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(_0110_),
    .X(net362));
 sky130_fd_sc_hd__clkbuf_2 hold143 (.A(\z80.tv80s.i_tv80_core.ts[4] ),
    .X(net363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(_0364_),
    .X(net364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][7] ),
    .X(net365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(_0099_),
    .X(net366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][3] ),
    .X(net367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(_0111_),
    .X(net368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][0] ),
    .X(net369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\z80.tv80s.i_tv80_core.RegBusA_r[11] ),
    .X(net235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(_0140_),
    .X(net370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][3] ),
    .X(net371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(_0151_),
    .X(net372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][7] ),
    .X(net373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(_0171_),
    .X(net374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][3] ),
    .X(net375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(_0346_),
    .X(net376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][4] ),
    .X(net377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(_0096_),
    .X(net378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][1] ),
    .X(net379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(_0301_),
    .X(net236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(_0125_),
    .X(net380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][1] ),
    .X(net381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(_0077_),
    .X(net382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][0] ),
    .X(net383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(_0067_),
    .X(net384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][3] ),
    .X(net385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(_0167_),
    .X(net386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][7] ),
    .X(net387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(_0115_),
    .X(net388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][6] ),
    .X(net389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\z80.tv80s.i_tv80_core.RegBusA_r[10] ),
    .X(net237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(_0349_),
    .X(net390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][1] ),
    .X(net391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(_0117_),
    .X(net392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][3] ),
    .X(net393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][3] ),
    .X(net394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(_0062_),
    .X(net395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][5] ),
    .X(net396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][4] ),
    .X(net397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(_0080_),
    .X(net398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(\z80.tv80s.i_tv80_core.Pre_XY_F_M[5] ),
    .X(net399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(_0300_),
    .X(net238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(_0010_),
    .X(net400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][5] ),
    .X(net401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(_0072_),
    .X(net402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][7] ),
    .X(net403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(_0066_),
    .X(net404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(\z80.tv80s.i_tv80_core.Auto_Wait_t2 ),
    .X(net405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(_0736_),
    .X(net406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][5] ),
    .X(net407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(_0097_),
    .X(net408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][2] ),
    .X(net409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\z80.tv80s.i_tv80_core.RegAddrA_r[1] ),
    .X(net239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][5] ),
    .X(net410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold191 (.A(_0113_),
    .X(net411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(\z80.tv80s.i_tv80_core.mcycles[5] ),
    .X(net412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(_0016_),
    .X(net413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][3] ),
    .X(net414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][1] ),
    .X(net415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(_0060_),
    .X(net416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold197 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][4] ),
    .X(net417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold198 (.A(_0120_),
    .X(net418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][1] ),
    .X(net419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(_0341_),
    .X(net222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(_0316_),
    .X(net240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(_0101_),
    .X(net420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][3] ),
    .X(net421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(_0143_),
    .X(net422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][3] ),
    .X(net423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][4] ),
    .X(net424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(_0168_),
    .X(net425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][3] ),
    .X(net426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][2] ),
    .X(net427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][5] ),
    .X(net428));
 sky130_fd_sc_hd__buf_1 hold209 (.A(\z80.tv80s.i_tv80_core.IncDecZ ),
    .X(net429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\z80.tv80s.i_tv80_core.RegBusA_r[13] ),
    .X(net241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold210 (.A(_0245_),
    .X(net430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][4] ),
    .X(net431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(_0104_),
    .X(net432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold213 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][4] ),
    .X(net433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold214 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][2] ),
    .X(net434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][7] ),
    .X(net435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(_0107_),
    .X(net436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold217 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][6] ),
    .X(net437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold218 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][1] ),
    .X(net438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold219 (.A(_0133_),
    .X(net439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(_0303_),
    .X(net242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][0] ),
    .X(net440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold221 (.A(_0164_),
    .X(net441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold222 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][5] ),
    .X(net442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold223 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][5] ),
    .X(net443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][2] ),
    .X(net444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold225 (.A(_0126_),
    .X(net445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold226 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][1] ),
    .X(net446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold227 (.A(_0109_),
    .X(net447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold228 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][6] ),
    .X(net448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold229 (.A(_0146_),
    .X(net449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\z80.tv80s.i_tv80_core.RegBusA_r[9] ),
    .X(net243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold230 (.A(\z80.tv80s.i_tv80_core.Z16_r ),
    .X(net450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold231 (.A(_0246_),
    .X(net451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold232 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][1] ),
    .X(net452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold233 (.A(_0041_),
    .X(net453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold234 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][7] ),
    .X(net454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold235 (.A(_0047_),
    .X(net455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold236 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][3] ),
    .X(net456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold237 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][0] ),
    .X(net457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(_0040_),
    .X(net458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold239 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][1] ),
    .X(net459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(_0299_),
    .X(net244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold240 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][6] ),
    .X(net460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(_0138_),
    .X(net461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold242 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][7] ),
    .X(net462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold243 (.A(_0139_),
    .X(net463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold244 (.A(\z80.tv80s.i_tv80_core.Read_To_Reg_r[3] ),
    .X(net464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold245 (.A(_0256_),
    .X(net465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold246 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][5] ),
    .X(net466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold247 (.A(\z80.tv80s.i_tv80_core.XY_State[0] ),
    .X(net467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold248 (.A(_0262_),
    .X(net468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold249 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][4] ),
    .X(net469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\z80.tv80s.i_tv80_core.RegBusA_r[12] ),
    .X(net245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold250 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][0] ),
    .X(net470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold251 (.A(_0343_),
    .X(net471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold252 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][4] ),
    .X(net472));
 sky130_fd_sc_hd__buf_1 hold253 (.A(\z80.tv80s.i_tv80_core.Alternate ),
    .X(net473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold254 (.A(_0281_),
    .X(net474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold255 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][7] ),
    .X(net475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold256 (.A(_0123_),
    .X(net476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold257 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][2] ),
    .X(net477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold258 (.A(\z80.tv80s.i_tv80_core.ISet[3] ),
    .X(net478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold259 (.A(_0003_),
    .X(net479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(_0302_),
    .X(net246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold260 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][7] ),
    .X(net480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold261 (.A(_0091_),
    .X(net481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold262 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][4] ),
    .X(net482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold263 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][5] ),
    .X(net483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold264 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][2] ),
    .X(net484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold265 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][5] ),
    .X(net485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold266 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][1] ),
    .X(net486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold267 (.A(_0344_),
    .X(net487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold268 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][0] ),
    .X(net488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold269 (.A(_0092_),
    .X(net489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\z80.tv80s.i_tv80_core.RegBusA_r[5] ),
    .X(net247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold270 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][5] ),
    .X(net490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold271 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][4] ),
    .X(net491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold272 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][2] ),
    .X(net492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold273 (.A(_0142_),
    .X(net493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold274 (.A(\z80.tv80s.i_tv80_core.R[7] ),
    .X(net494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold275 (.A(_0314_),
    .X(net495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold276 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][0] ),
    .X(net496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold277 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][7] ),
    .X(net497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold278 (.A(_0163_),
    .X(net498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold279 (.A(\z80.tv80s.i_tv80_core.Pre_XY_F_M[3] ),
    .X(net499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(_0295_),
    .X(net248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold280 (.A(_0008_),
    .X(net500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold281 (.A(\z80.tv80s.i_tv80_core.Read_To_Reg_r[2] ),
    .X(net501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold282 (.A(_0255_),
    .X(net502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold283 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][0] ),
    .X(net503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold284 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][7] ),
    .X(net504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold285 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][3] ),
    .X(net505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold286 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][4] ),
    .X(net506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold287 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][2] ),
    .X(net507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold288 (.A(\z80.tv80s.i_tv80_core.Read_To_Reg_r[1] ),
    .X(net508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold289 (.A(_0254_),
    .X(net509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\z80.tv80s.i_tv80_core.RegBusA_r[2] ),
    .X(net249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold290 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][7] ),
    .X(net510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold291 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][0] ),
    .X(net511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold292 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][1] ),
    .X(net512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold293 (.A(_0141_),
    .X(net513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold294 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][2] ),
    .X(net514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold295 (.A(_0345_),
    .X(net515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold296 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][4] ),
    .X(net516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold297 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][4] ),
    .X(net517));
 sky130_fd_sc_hd__buf_1 hold298 (.A(\z80.tv80s.i_tv80_core.NMI_s ),
    .X(net518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold299 (.A(_0342_),
    .X(net519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\z80.tv80s.i_tv80_core.RegBusA_r[4] ),
    .X(net223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(_0292_),
    .X(net250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold300 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][7] ),
    .X(net520));
 sky130_fd_sc_hd__buf_1 hold301 (.A(net881),
    .X(net521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold302 (.A(_0012_),
    .X(net522));
 sky130_fd_sc_hd__clkbuf_2 hold303 (.A(\z80.tv80s.i_tv80_core.i_mcode.MCycle[4] ),
    .X(net523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold304 (.A(_0588_),
    .X(net524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold305 (.A(_0593_),
    .X(net525));
 sky130_fd_sc_hd__buf_1 hold306 (.A(net878),
    .X(net526));
 sky130_fd_sc_hd__clkbuf_2 hold307 (.A(\z80.tv80s.i_tv80_core.R[3] ),
    .X(net527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold308 (.A(_0052_),
    .X(net528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold309 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][2] ),
    .X(net529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\z80.tv80s.i_tv80_core.RegBusA_r[6] ),
    .X(net251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold310 (.A(net48),
    .X(net530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold311 (.A(_0205_),
    .X(net531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold312 (.A(net44),
    .X(net532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold313 (.A(_0211_),
    .X(net533));
 sky130_fd_sc_hd__buf_1 hold314 (.A(\z80.tv80s.i_tv80_core.XY_Ind ),
    .X(net534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold315 (.A(_2251_),
    .X(net535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold316 (.A(net42),
    .X(net536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold317 (.A(_0208_),
    .X(net537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold318 (.A(net43),
    .X(net538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold319 (.A(_0210_),
    .X(net539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(_0296_),
    .X(net252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold320 (.A(net41),
    .X(net540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold321 (.A(_0209_),
    .X(net541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold322 (.A(\z80.tv80s.i_tv80_core.RegAddrB_r[1] ),
    .X(net542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold323 (.A(_0260_),
    .X(net543));
 sky130_fd_sc_hd__buf_1 hold324 (.A(\z80.tv80s.i_tv80_core.R[2] ),
    .X(net544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold325 (.A(_0051_),
    .X(net545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold326 (.A(net45),
    .X(net546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold327 (.A(_0207_),
    .X(net547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold328 (.A(\z80.tv80s.i_tv80_core.mcycles[4] ),
    .X(net548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold329 (.A(_0015_),
    .X(net549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\z80.tv80s.i_tv80_core.RegBusA_r[3] ),
    .X(net253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold330 (.A(net46),
    .X(net550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold331 (.A(_0212_),
    .X(net551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold332 (.A(\z80.tv80s.i_tv80_core.RegAddrB_r[2] ),
    .X(net552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold333 (.A(_0056_),
    .X(net553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold334 (.A(net47),
    .X(net554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold335 (.A(_0206_),
    .X(net555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold336 (.A(net33),
    .X(net556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold337 (.A(_0230_),
    .X(net557));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold338 (.A(\z80.tv80s.i_tv80_core.R[0] ),
    .X(net558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold339 (.A(_0049_),
    .X(net559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(_0293_),
    .X(net254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold340 (.A(net57),
    .X(net560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold341 (.A(_0223_),
    .X(net561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold342 (.A(\z80.tv80s.i_tv80_core.RegBusA_r[1] ),
    .X(net562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold343 (.A(\z80.tv80s.i_tv80_core.RegBusA_r[0] ),
    .X(net563));
 sky130_fd_sc_hd__clkbuf_2 hold344 (.A(\z80.tv80s.i_tv80_core.R[5] ),
    .X(net564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold345 (.A(_0054_),
    .X(net565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold346 (.A(\z80.tv80s.i_tv80_core.XY_State[1] ),
    .X(net566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold347 (.A(\z80.tv80s.i_tv80_core.ISet[1] ),
    .X(net567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold348 (.A(_0001_),
    .X(net568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold349 (.A(net58),
    .X(net569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\z80.tv80s.i_tv80_core.Pre_XY_F_M[1] ),
    .X(net255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold350 (.A(_0221_),
    .X(net570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold351 (.A(net29),
    .X(net571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold352 (.A(_0226_),
    .X(net572));
 sky130_fd_sc_hd__clkbuf_2 hold353 (.A(net880),
    .X(net573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold354 (.A(_0361_),
    .X(net574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold355 (.A(net56),
    .X(net575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold356 (.A(_0224_),
    .X(net576));
 sky130_fd_sc_hd__buf_1 hold357 (.A(\z80.tv80s.i_tv80_core.PC[5] ),
    .X(net577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold358 (.A(_0322_),
    .X(net578));
 sky130_fd_sc_hd__buf_1 hold359 (.A(\z80.tv80s.i_tv80_core.I[4] ),
    .X(net579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(_0006_),
    .X(net256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold360 (.A(_0310_),
    .X(net580));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold361 (.A(\z80.tv80s.i_tv80_core.I[0] ),
    .X(net581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold362 (.A(_0306_),
    .X(net582));
 sky130_fd_sc_hd__buf_1 hold363 (.A(\z80.tv80s.i_tv80_core.SP[10] ),
    .X(net583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold364 (.A(_0376_),
    .X(net584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold365 (.A(\z80.tv80s.i_tv80_core.IStatus[1] ),
    .X(net585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold366 (.A(_0004_),
    .X(net586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold367 (.A(net28),
    .X(net587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold368 (.A(_0222_),
    .X(net588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold369 (.A(net35),
    .X(net589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\z80.tv80s.i_tv80_core.Pre_XY_F_M[4] ),
    .X(net257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold370 (.A(_0232_),
    .X(net590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold371 (.A(net55),
    .X(net591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold372 (.A(_0225_),
    .X(net592));
 sky130_fd_sc_hd__buf_1 hold373 (.A(\z80.tv80s.i_tv80_core.TmpAddr[8] ),
    .X(net593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold374 (.A(_0273_),
    .X(net594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold375 (.A(\z80.tv80s.i_tv80_core.PC[3] ),
    .X(net595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold376 (.A(_0320_),
    .X(net596));
 sky130_fd_sc_hd__buf_2 hold377 (.A(\z80.tv80s.i_tv80_core.RegAddrC[2] ),
    .X(net597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold378 (.A(_0057_),
    .X(net598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold379 (.A(\z80.tv80s.i_tv80_core.PC[4] ),
    .X(net599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(_0009_),
    .X(net258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold380 (.A(_0321_),
    .X(net600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold381 (.A(net30),
    .X(net601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold382 (.A(_0227_),
    .X(net602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold383 (.A(net31),
    .X(net603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold384 (.A(_0228_),
    .X(net604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold385 (.A(\z80.tv80s.i_tv80_core.ts[0] ),
    .X(net605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold386 (.A(_0032_),
    .X(net606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold387 (.A(net34),
    .X(net607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold388 (.A(_0231_),
    .X(net608));
 sky130_fd_sc_hd__buf_2 hold389 (.A(\z80.tv80s.i_tv80_core.i_mcode.MCycle[5] ),
    .X(net609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\z80.tv80s.i_tv80_core.Pre_XY_F_M[2] ),
    .X(net259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold390 (.A(_0030_),
    .X(net610));
 sky130_fd_sc_hd__buf_1 hold391 (.A(\z80.tv80s.i_tv80_core.TmpAddr[9] ),
    .X(net611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold392 (.A(_0274_),
    .X(net612));
 sky130_fd_sc_hd__buf_1 hold393 (.A(\z80.tv80s.i_tv80_core.R[4] ),
    .X(net613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold394 (.A(_0053_),
    .X(net614));
 sky130_fd_sc_hd__buf_1 hold395 (.A(\z80.tv80s.i_tv80_core.R[1] ),
    .X(net615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold396 (.A(_0050_),
    .X(net616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold397 (.A(\z80.tv80s.i_tv80_core.PC[2] ),
    .X(net617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold398 (.A(_0319_),
    .X(net618));
 sky130_fd_sc_hd__buf_1 hold399 (.A(\z80.tv80s.i_tv80_core.BusB[6] ),
    .X(net619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(_0294_),
    .X(net224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(_0007_),
    .X(net260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold400 (.A(_0288_),
    .X(net620));
 sky130_fd_sc_hd__clkbuf_2 hold401 (.A(\z80.tv80s.i_tv80_core.NMICycle ),
    .X(net621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold402 (.A(_0196_),
    .X(net622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold403 (.A(\z80.tv80s.i_tv80_core.I[2] ),
    .X(net623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold404 (.A(_0308_),
    .X(net624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold405 (.A(\z80.tv80s.i_tv80_core.Arith16_r ),
    .X(net625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold406 (.A(_0258_),
    .X(net626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold407 (.A(\z80.tv80s.i_tv80_core.I[3] ),
    .X(net627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold408 (.A(_0309_),
    .X(net628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold409 (.A(net40),
    .X(net629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\z80.tv80s.i_tv80_core.RegAddrA_r[0] ),
    .X(net261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold410 (.A(_0236_),
    .X(net630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold411 (.A(net36),
    .X(net631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold412 (.A(_0233_),
    .X(net632));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold413 (.A(\z80.tv80s.i_tv80_core.Read_To_Reg_r[0] ),
    .X(net633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold414 (.A(_0253_),
    .X(net634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold415 (.A(net32),
    .X(net635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold416 (.A(_0229_),
    .X(net636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold417 (.A(\z80.tv80s.i_tv80_core.SP[0] ),
    .X(net637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold418 (.A(_0366_),
    .X(net638));
 sky130_fd_sc_hd__buf_1 hold419 (.A(\z80.tv80s.i_tv80_core.BusB[7] ),
    .X(net639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(_0315_),
    .X(net262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold420 (.A(_0289_),
    .X(net640));
 sky130_fd_sc_hd__buf_1 hold421 (.A(\z80.tv80s.i_tv80_core.PC[0] ),
    .X(net641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold422 (.A(_0317_),
    .X(net642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold423 (.A(\z80.tv80s.i_tv80_core.BusB[5] ),
    .X(net643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold424 (.A(_0287_),
    .X(net644));
 sky130_fd_sc_hd__buf_1 hold425 (.A(\z80.tv80s.i_tv80_core.BusB[1] ),
    .X(net645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold426 (.A(_0283_),
    .X(net646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold427 (.A(net37),
    .X(net647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold428 (.A(_0234_),
    .X(net648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold429 (.A(\z80.tv80s.i_tv80_core.BusB[3] ),
    .X(net649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\z80.tv80s.i_tv80_core.BTR_r ),
    .X(net263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold430 (.A(_0285_),
    .X(net650));
 sky130_fd_sc_hd__clkbuf_2 hold431 (.A(\z80.tv80s.i_tv80_core.i_mcode.MCycle[6] ),
    .X(net651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold432 (.A(_0591_),
    .X(net652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold433 (.A(_0029_),
    .X(net653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold434 (.A(\z80.tv80s.i_tv80_core.Ap[7] ),
    .X(net654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold435 (.A(_0179_),
    .X(net655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold436 (.A(\z80.tv80s.i_tv80_core.Ap[1] ),
    .X(net656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold437 (.A(_0173_),
    .X(net657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold438 (.A(\z80.tv80s.i_tv80_core.Ap[6] ),
    .X(net658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold439 (.A(_0178_),
    .X(net659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(_0252_),
    .X(net264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold440 (.A(\z80.tv80s.i_tv80_core.SP[6] ),
    .X(net660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold441 (.A(_0372_),
    .X(net661));
 sky130_fd_sc_hd__buf_1 hold442 (.A(\z80.tv80s.i_tv80_core.SP[4] ),
    .X(net662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold443 (.A(_0370_),
    .X(net663));
 sky130_fd_sc_hd__buf_1 hold444 (.A(\z80.tv80s.i_tv80_core.SP[8] ),
    .X(net664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold445 (.A(_0374_),
    .X(net665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold446 (.A(\z80.tv80s.i_tv80_core.Fp[7] ),
    .X(net666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold447 (.A(_0187_),
    .X(net667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold448 (.A(\z80.tv80s.i_tv80_core.Fp[2] ),
    .X(net668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold449 (.A(_0182_),
    .X(net669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\z80.tv80s.i_tv80_core.ts[6] ),
    .X(net265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold450 (.A(\z80.tv80s.i_tv80_core.Fp[4] ),
    .X(net670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold451 (.A(_0184_),
    .X(net671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold452 (.A(\z80.tv80s.i_tv80_core.BusA[0] ),
    .X(net672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold453 (.A(_0188_),
    .X(net673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold454 (.A(\z80.tv80s.i_tv80_core.Ap[5] ),
    .X(net674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold455 (.A(_0177_),
    .X(net675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold456 (.A(\z80.tv80s.i_tv80_core.I[1] ),
    .X(net676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold457 (.A(_0307_),
    .X(net677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold458 (.A(\z80.tv80s.i_tv80_core.Ap[4] ),
    .X(net678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold459 (.A(_0176_),
    .X(net679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(_0359_),
    .X(net266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold460 (.A(\z80.tv80s.i_tv80_core.SP[1] ),
    .X(net680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold461 (.A(_0367_),
    .X(net681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold462 (.A(\z80.tv80s.i_tv80_core.Ap[2] ),
    .X(net682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold463 (.A(_0174_),
    .X(net683));
 sky130_fd_sc_hd__buf_1 hold464 (.A(\z80.tv80s.i_tv80_core.R[6] ),
    .X(net684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold465 (.A(_0055_),
    .X(net685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold466 (.A(\z80.tv80s.i_tv80_core.Ap[0] ),
    .X(net686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold467 (.A(_0172_),
    .X(net687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold468 (.A(\z80.tv80s.i_tv80_core.SP[13] ),
    .X(net688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold469 (.A(_0379_),
    .X(net689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\z80.tv80s.i_tv80_core.Pre_XY_F_M[6] ),
    .X(net267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold470 (.A(\z80.tv80s.i_tv80_core.BusA[3] ),
    .X(net690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold471 (.A(_0191_),
    .X(net691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold472 (.A(\z80.tv80s.i_tv80_core.i_mcode.MCycle[3] ),
    .X(net692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold473 (.A(_0336_),
    .X(net693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold474 (.A(\z80.tv80s.i_tv80_core.PC[1] ),
    .X(net694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold475 (.A(_0318_),
    .X(net695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold476 (.A(\z80.tv80s.i_tv80_core.Ap[3] ),
    .X(net696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold477 (.A(_0175_),
    .X(net697));
 sky130_fd_sc_hd__clkbuf_2 hold478 (.A(_0036_),
    .X(net698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold479 (.A(_2774_),
    .X(net699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(_0011_),
    .X(net268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold480 (.A(_0339_),
    .X(net700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold481 (.A(\z80.tv80s.i_tv80_core.Fp[6] ),
    .X(net701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold482 (.A(_0186_),
    .X(net702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold483 (.A(\z80.tv80s.i_tv80_core.SP[3] ),
    .X(net703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold484 (.A(_0369_),
    .X(net704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold485 (.A(\z80.tv80s.i_tv80_core.Fp[5] ),
    .X(net705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold486 (.A(_0185_),
    .X(net706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold487 (.A(\z80.tv80s.i_tv80_core.BusA[4] ),
    .X(net707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold488 (.A(_0192_),
    .X(net708));
 sky130_fd_sc_hd__clkbuf_2 hold489 (.A(\z80.tv80s.i_tv80_core.BusB[0] ),
    .X(net709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\z80.tv80s.i_tv80_core.IStatus[2] ),
    .X(net269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold490 (.A(_0282_),
    .X(net710));
 sky130_fd_sc_hd__buf_1 hold491 (.A(\z80.tv80s.i_tv80_core.Halt_FF ),
    .X(net711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold492 (.A(_0024_),
    .X(net712));
 sky130_fd_sc_hd__buf_1 hold493 (.A(\z80.tv80s.i_tv80_core.SP[2] ),
    .X(net713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold494 (.A(_0368_),
    .X(net714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold495 (.A(\z80.tv80s.i_tv80_core.No_BTR ),
    .X(net715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold496 (.A(_0719_),
    .X(net716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold497 (.A(_0334_),
    .X(net717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold498 (.A(\z80.tv80s.i_tv80_core.SP[5] ),
    .X(net718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold499 (.A(_0371_),
    .X(net719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\z80.tv80s.i_tv80_core.RegAddrA_r[2] ),
    .X(net225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(_0005_),
    .X(net270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold500 (.A(\z80.tv80s.i_tv80_core.Read_To_Reg_r[4] ),
    .X(net720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold501 (.A(_0257_),
    .X(net721));
 sky130_fd_sc_hd__buf_1 hold502 (.A(\z80.tv80s.i_tv80_core.I[5] ),
    .X(net722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold503 (.A(_0311_),
    .X(net723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold504 (.A(net39),
    .X(net724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold505 (.A(_0235_),
    .X(net725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold506 (.A(\z80.tv80s.i_tv80_core.BusA[5] ),
    .X(net726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold507 (.A(_0193_),
    .X(net727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold508 (.A(\z80.tv80s.i_tv80_core.BusB[4] ),
    .X(net728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold509 (.A(_0286_),
    .X(net729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][6] ),
    .X(net271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold510 (.A(\z80.tv80s.i_tv80_core.Fp[3] ),
    .X(net730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold511 (.A(_0183_),
    .X(net731));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold512 (.A(\z80.tv80s.i_tv80_core.I[6] ),
    .X(net732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold513 (.A(_0312_),
    .X(net733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold514 (.A(\z80.tv80s.i_tv80_core.Fp[0] ),
    .X(net734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold515 (.A(_0180_),
    .X(net735));
 sky130_fd_sc_hd__clkbuf_2 hold516 (.A(\z80.tv80s.i_tv80_core.ts[3] ),
    .X(net736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold517 (.A(_0363_),
    .X(net737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold518 (.A(\z80.tv80s.i_tv80_core.PC[7] ),
    .X(net738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold519 (.A(_0324_),
    .X(net739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(_0154_),
    .X(net272));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold520 (.A(\z80.tv80s.i_tv80_core.SP[9] ),
    .X(net740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold521 (.A(_0375_),
    .X(net741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold522 (.A(\z80.tv80s.i_tv80_core.SP[11] ),
    .X(net742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold523 (.A(_0377_),
    .X(net743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold524 (.A(\z80.tv80s.i_tv80_core.PC[6] ),
    .X(net744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold525 (.A(_0323_),
    .X(net745));
 sky130_fd_sc_hd__buf_2 hold526 (.A(\z80.tv80s.i_tv80_core.BusAck ),
    .X(net746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold527 (.A(\z80.tv80s.i_tv80_core.Fp[1] ),
    .X(net747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold528 (.A(_0181_),
    .X(net748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold529 (.A(\z80.tv80s.i_tv80_core.BusA[2] ),
    .X(net749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][6] ),
    .X(net273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold530 (.A(_0190_),
    .X(net750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold531 (.A(\z80.tv80s.i_tv80_core.TmpAddr[14] ),
    .X(net751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold532 (.A(_0279_),
    .X(net752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold533 (.A(\z80.tv80s.i_tv80_core.TmpAddr[12] ),
    .X(net753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold534 (.A(_0277_),
    .X(net754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold535 (.A(\z80.tv80s.i_tv80_core.SP[12] ),
    .X(net755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold536 (.A(_0378_),
    .X(net756));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold537 (.A(\z80.tv80s.i_tv80_core.PC[15] ),
    .X(net757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold538 (.A(_0332_),
    .X(net758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold539 (.A(\z80.tv80s.i_tv80_core.TmpAddr[15] ),
    .X(net759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(_0106_),
    .X(net274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold540 (.A(_0280_),
    .X(net760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold541 (.A(\z80.tv80s.i_tv80_core.TmpAddr[10] ),
    .X(net761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold542 (.A(_0275_),
    .X(net762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold543 (.A(\z80.tv80s.i_tv80_core.IntE ),
    .X(net763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold544 (.A(_0731_),
    .X(net764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold545 (.A(_0026_),
    .X(net765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold546 (.A(\z80.tv80s.i_tv80_core.PC[14] ),
    .X(net766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold547 (.A(_0331_),
    .X(net767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold548 (.A(\z80.tv80s.i_tv80_core.BusA[6] ),
    .X(net768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold549 (.A(_0194_),
    .X(net769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][0] ),
    .X(net275));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold550 (.A(_0035_),
    .X(net770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold551 (.A(_2761_),
    .X(net771));
 sky130_fd_sc_hd__buf_1 hold552 (.A(\z80.tv80s.i_tv80_core.PC[12] ),
    .X(net772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold553 (.A(_0329_),
    .X(net773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold554 (.A(\z80.tv80s.i_tv80_core.BusB[2] ),
    .X(net774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold555 (.A(_0284_),
    .X(net775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold556 (.A(\z80.tv80s.i_tv80_core.TmpAddr[11] ),
    .X(net776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold557 (.A(_0276_),
    .X(net777));
 sky130_fd_sc_hd__clkbuf_2 hold558 (.A(\z80.tv80s.i_tv80_core.IntCycle ),
    .X(net778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold559 (.A(_0340_),
    .X(net779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(_0100_),
    .X(net276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold560 (.A(\z80.tv80s.i_tv80_core.PC[13] ),
    .X(net780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold561 (.A(_0330_),
    .X(net781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold562 (.A(\z80.tv80s.i_tv80_core.TmpAddr[13] ),
    .X(net782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold563 (.A(_0278_),
    .X(net783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold564 (.A(\z80.tv80s.i_tv80_core.BusA[1] ),
    .X(net784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold565 (.A(_0189_),
    .X(net785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold566 (.A(\z80.tv80s.i_tv80_core.i_mcode.MCycle[2] ),
    .X(net786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold567 (.A(_0335_),
    .X(net787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold568 (.A(\z80.tv80s.i_tv80_core.PC[9] ),
    .X(net788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold569 (.A(_0326_),
    .X(net789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][0] ),
    .X(net277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold570 (.A(\z80.tv80s.i_tv80_core.TmpAddr[1] ),
    .X(net790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold571 (.A(_0266_),
    .X(net791));
 sky130_fd_sc_hd__clkbuf_2 hold572 (.A(\z80.tv80s.i_tv80_core.I[7] ),
    .X(net792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold573 (.A(_0313_),
    .X(net793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold574 (.A(\z80.tv80s.i_tv80_core.IR[5] ),
    .X(net794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold575 (.A(_2935_),
    .X(net795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold576 (.A(_0000_),
    .X(net796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold577 (.A(_0034_),
    .X(net797));
 sky130_fd_sc_hd__buf_1 hold578 (.A(\z80.tv80s.i_tv80_core.SP[7] ),
    .X(net798));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold579 (.A(\z80.tv80s.i_tv80_core.PC[11] ),
    .X(net799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(_0148_),
    .X(net278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold580 (.A(_0328_),
    .X(net800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold581 (.A(\z80.tv80s.i_tv80_core.TmpAddr[0] ),
    .X(net801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold582 (.A(_0265_),
    .X(net802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold583 (.A(\z80.tv80s.i_tv80_core.TmpAddr[2] ),
    .X(net803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold584 (.A(_0267_),
    .X(net804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold585 (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ),
    .X(net805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold586 (.A(\z80.tv80s.i_tv80_core.PC[10] ),
    .X(net806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold587 (.A(_0327_),
    .X(net807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold588 (.A(\z80.tv80s.i_tv80_core.PC[8] ),
    .X(net808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold589 (.A(_0325_),
    .X(net809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(\z80.tv80s.i_tv80_core.mcycles[2] ),
    .X(net279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold590 (.A(\z80.tv80s.i_tv80_core.TmpAddr[6] ),
    .X(net810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold591 (.A(_0271_),
    .X(net811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold592 (.A(\z80.tv80s.i_tv80_core.TmpAddr[7] ),
    .X(net812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold593 (.A(_0272_),
    .X(net813));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold594 (.A(\z80.tv80s.i_tv80_core.SP[15] ),
    .X(net814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold595 (.A(\z80.tv80s.i_tv80_core.TmpAddr[4] ),
    .X(net815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold596 (.A(_0269_),
    .X(net816));
 sky130_fd_sc_hd__buf_1 hold597 (.A(\z80.tv80s.i_tv80_core.SP[14] ),
    .X(net817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold598 (.A(\z80.tv80s.i_tv80_core.F[5] ),
    .X(net818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold599 (.A(\z80.tv80s.i_tv80_core.mcycles[1] ),
    .X(net819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(_0048_),
    .X(net226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(_0014_),
    .X(net280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold600 (.A(_0013_),
    .X(net820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold601 (.A(\z80.tv80s.i_tv80_core.TmpAddr[5] ),
    .X(net821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold602 (.A(_0270_),
    .X(net822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold603 (.A(\z80.tv80s.i_tv80_core.F[3] ),
    .X(net823));
 sky130_fd_sc_hd__clkbuf_2 hold604 (.A(\z80.tv80s.i_tv80_core.ISet[2] ),
    .X(net824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold605 (.A(_2220_),
    .X(net825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold606 (.A(_0248_),
    .X(net826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold607 (.A(\z80.tv80s.i_tv80_core.TmpAddr[3] ),
    .X(net827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold608 (.A(_0268_),
    .X(net828));
 sky130_fd_sc_hd__buf_2 hold609 (.A(\z80.tv80s.i_tv80_core.ts[2] ),
    .X(net829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][7] ),
    .X(net281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold610 (.A(\z80.tv80s.i_tv80_core.F[4] ),
    .X(net830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold611 (.A(\z80.tv80s.i_tv80_core.IR[1] ),
    .X(net831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold612 (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[2] ),
    .X(net832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold613 (.A(\z80.tv80s.i_tv80_core.F[7] ),
    .X(net833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold614 (.A(_0244_),
    .X(net834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold615 (.A(\z80.tv80s.i_tv80_core.IR[6] ),
    .X(net835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold616 (.A(\z80.tv80s.di_reg[0] ),
    .X(net836));
 sky130_fd_sc_hd__buf_1 hold617 (.A(\z80.tv80s.i_tv80_core.Save_ALU_r ),
    .X(net837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold618 (.A(\z80.tv80s.di_reg[1] ),
    .X(net838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold619 (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[0] ),
    .X(net839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(_0155_),
    .X(net282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold620 (.A(\z80.tv80s.di_reg[5] ),
    .X(net840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold621 (.A(\z80.tv80s.di_reg[4] ),
    .X(net841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold622 (.A(\z80.tv80s.i_tv80_core.IntE_FF2 ),
    .X(net842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold623 (.A(_0027_),
    .X(net843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold624 (.A(\z80.tv80s.di_reg[3] ),
    .X(net844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold625 (.A(\z80.tv80s.i_tv80_core.IR[7] ),
    .X(net845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold626 (.A(\z80.tv80s.di_reg[2] ),
    .X(net846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold627 (.A(\z80.tv80s.di_reg[6] ),
    .X(net847));
 sky130_fd_sc_hd__buf_1 hold628 (.A(\z80.tv80s.di_reg[7] ),
    .X(net848));
 sky130_fd_sc_hd__buf_1 hold629 (.A(\z80.tv80s.i_tv80_core.ACC[7] ),
    .X(net849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][1] ),
    .X(net283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold630 (.A(\z80.tv80s.i_tv80_core.ACC[1] ),
    .X(net850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold631 (.A(\z80.tv80s.i_tv80_core.ACC[4] ),
    .X(net851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold632 (.A(\z80.tv80s.i_tv80_core.ACC[0] ),
    .X(net852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold633 (.A(_0213_),
    .X(net853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold634 (.A(\z80.tv80s.i_tv80_core.F[6] ),
    .X(net854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold635 (.A(\z80.tv80s.i_tv80_core.ACC[2] ),
    .X(net855));
 sky130_fd_sc_hd__buf_1 hold636 (.A(\z80.tv80s.i_tv80_core.F[2] ),
    .X(net856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold637 (.A(\z80.tv80s.i_tv80_core.ACC[6] ),
    .X(net857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold638 (.A(\z80.tv80s.i_tv80_core.i_mcode.MCycle[0] ),
    .X(net858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold639 (.A(\z80.tv80s.i_tv80_core.ACC[5] ),
    .X(net859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(_0085_),
    .X(net284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold640 (.A(\z80.tv80s.i_tv80_core.ts[2] ),
    .X(net860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold641 (.A(\z80.tv80s.i_tv80_core.RegAddrC[1] ),
    .X(net861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold642 (.A(\z80.tv80s.i_tv80_core.ACC[3] ),
    .X(net862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold643 (.A(\z80.tv80s.i_tv80_core.F[0] ),
    .X(net863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold644 (.A(\z80.tv80s.i_tv80_core.RegAddrC[0] ),
    .X(net864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold645 (.A(\z80.tv80s.i_tv80_core.F[1] ),
    .X(net865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold646 (.A(\z80.tv80s.i_tv80_core.IR[2] ),
    .X(net866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold647 (.A(\z80.tv80s.i_tv80_core.IR[3] ),
    .X(net867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold648 (.A(\z80.tv80s.i_tv80_core.IR[4] ),
    .X(net868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold649 (.A(\z80.tv80s.i_tv80_core.IR[0] ),
    .X(net869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][0] ),
    .X(net285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold650 (.A(\z80.tv80s.i_tv80_core.BusA[7] ),
    .X(net870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold651 (.A(_0195_),
    .X(net871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold652 (.A(\z80.tv80s.i_tv80_core.RegAddrB_r[0] ),
    .X(net872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold653 (.A(\z80.tv80s.i_tv80_core.Read_To_Reg_r[0] ),
    .X(net873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold654 (.A(\z80.tv80s.i_tv80_core.ts[4] ),
    .X(net874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold655 (.A(\z80.tv80s.i_tv80_core.i_mcode.MCycle[0] ),
    .X(net875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold656 (.A(\z80.tv80s.i_tv80_core.IR[3] ),
    .X(net876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold657 (.A(\z80.tv80s.i_tv80_core.Save_ALU_r ),
    .X(net877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold658 (.A(\z80.tv80s.i_tv80_core.PreserveC_r ),
    .X(net878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold659 (.A(\z80.tv80s.i_tv80_core.Auto_Wait_t1 ),
    .X(net879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(_0084_),
    .X(net286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold660 (.A(\z80.tv80s.i_tv80_core.ts[1] ),
    .X(net880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold661 (.A(\z80.tv80s.i_tv80_core.Pre_XY_F_M[7] ),
    .X(net881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][5] ),
    .X(net287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(_0129_),
    .X(net288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][2] ),
    .X(net289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\z80.tv80s.i_tv80_core.RegBusA_r[14] ),
    .X(net227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(_0150_),
    .X(net290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][6] ),
    .X(net291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(_0162_),
    .X(net292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][3] ),
    .X(net293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(_0079_),
    .X(net294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][0] ),
    .X(net295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(_0116_),
    .X(net296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(\z80.tv80s.i_tv80_core.ts[5] ),
    .X(net297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(_0365_),
    .X(net298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][1] ),
    .X(net299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(_0304_),
    .X(net228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(_0157_),
    .X(net300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][3] ),
    .X(net301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(_0103_),
    .X(net302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][1] ),
    .X(net303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(_0149_),
    .X(net304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][4] ),
    .X(net305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(_0152_),
    .X(net306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][0] ),
    .X(net307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(_0156_),
    .X(net308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][6] ),
    .X(net309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\z80.tv80s.i_tv80_core.RegBusA_r[8] ),
    .X(net229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(_0130_),
    .X(net310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][1] ),
    .X(net311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(_0068_),
    .X(net312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][2] ),
    .X(net313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(_0078_),
    .X(net314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][2] ),
    .X(net315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(_0069_),
    .X(net316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][6] ),
    .X(net317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(_0090_),
    .X(net318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][5] ),
    .X(net319));
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(custom_settings[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(io_in[26]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_2 input11 (.A(io_in[27]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_2 input12 (.A(io_in[28]),
    .X(net12));
 sky130_fd_sc_hd__buf_2 input13 (.A(io_in[29]),
    .X(net13));
 sky130_fd_sc_hd__buf_1 input14 (.A(io_in[30]),
    .X(net14));
 sky130_fd_sc_hd__buf_1 input15 (.A(io_in[31]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(io_in[35]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_4 input17 (.A(io_in[4]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_4 input18 (.A(rst_n),
    .X(net18));
 sky130_fd_sc_hd__buf_1 input2 (.A(custom_settings[1]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(custom_settings[2]),
    .X(net3));
 sky130_fd_sc_hd__buf_1 input4 (.A(custom_settings[3]),
    .X(net4));
 sky130_fd_sc_hd__buf_1 input5 (.A(custom_settings[4]),
    .X(net5));
 sky130_fd_sc_hd__dlymetal6s2s_1 input6 (.A(io_in[22]),
    .X(net6));
 sky130_fd_sc_hd__buf_1 input7 (.A(io_in[23]),
    .X(net7));
 sky130_fd_sc_hd__dlymetal6s2s_1 input8 (.A(io_in[24]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_2 input9 (.A(io_in[25]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_4 max_cap62 (.A(_1688_),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_4 max_cap71 (.A(_0798_),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_2 max_cap91 (.A(net92),
    .X(net91));
 sky130_fd_sc_hd__buf_12 output19 (.A(net19),
    .X(io_oeb[22]));
 sky130_fd_sc_hd__buf_12 output20 (.A(net20),
    .X(io_oeb[23]));
 sky130_fd_sc_hd__buf_12 output21 (.A(net21),
    .X(io_oeb[24]));
 sky130_fd_sc_hd__buf_12 output22 (.A(net22),
    .X(io_oeb[25]));
 sky130_fd_sc_hd__buf_12 output23 (.A(net23),
    .X(io_oeb[26]));
 sky130_fd_sc_hd__buf_12 output24 (.A(net24),
    .X(io_oeb[27]));
 sky130_fd_sc_hd__buf_12 output25 (.A(net25),
    .X(io_oeb[28]));
 sky130_fd_sc_hd__buf_12 output26 (.A(net26),
    .X(io_oeb[29]));
 sky130_fd_sc_hd__buf_12 output27 (.A(net117),
    .X(io_out[0]));
 sky130_fd_sc_hd__buf_12 output28 (.A(net28),
    .X(io_out[10]));
 sky130_fd_sc_hd__buf_12 output29 (.A(net29),
    .X(io_out[11]));
 sky130_fd_sc_hd__buf_12 output30 (.A(net30),
    .X(io_out[12]));
 sky130_fd_sc_hd__buf_12 output31 (.A(net31),
    .X(io_out[13]));
 sky130_fd_sc_hd__buf_12 output32 (.A(net32),
    .X(io_out[14]));
 sky130_fd_sc_hd__buf_12 output33 (.A(net33),
    .X(io_out[15]));
 sky130_fd_sc_hd__buf_12 output34 (.A(net34),
    .X(io_out[16]));
 sky130_fd_sc_hd__buf_12 output35 (.A(net35),
    .X(io_out[17]));
 sky130_fd_sc_hd__buf_12 output36 (.A(net36),
    .X(io_out[18]));
 sky130_fd_sc_hd__buf_12 output37 (.A(net37),
    .X(io_out[19]));
 sky130_fd_sc_hd__buf_12 output38 (.A(net38),
    .X(io_out[1]));
 sky130_fd_sc_hd__buf_12 output39 (.A(net39),
    .X(io_out[20]));
 sky130_fd_sc_hd__buf_12 output40 (.A(net40),
    .X(io_out[21]));
 sky130_fd_sc_hd__buf_12 output41 (.A(net41),
    .X(io_out[22]));
 sky130_fd_sc_hd__buf_12 output42 (.A(net42),
    .X(io_out[23]));
 sky130_fd_sc_hd__buf_12 output43 (.A(net43),
    .X(io_out[24]));
 sky130_fd_sc_hd__buf_12 output44 (.A(net44),
    .X(io_out[25]));
 sky130_fd_sc_hd__buf_12 output45 (.A(net45),
    .X(io_out[26]));
 sky130_fd_sc_hd__buf_12 output46 (.A(net46),
    .X(io_out[27]));
 sky130_fd_sc_hd__buf_12 output47 (.A(net47),
    .X(io_out[28]));
 sky130_fd_sc_hd__buf_12 output48 (.A(net48),
    .X(io_out[29]));
 sky130_fd_sc_hd__buf_12 output49 (.A(net49),
    .X(io_out[2]));
 sky130_fd_sc_hd__buf_12 output50 (.A(net50),
    .X(io_out[32]));
 sky130_fd_sc_hd__buf_12 output51 (.A(net51),
    .X(io_out[33]));
 sky130_fd_sc_hd__buf_12 output52 (.A(net52),
    .X(io_out[34]));
 sky130_fd_sc_hd__buf_12 output53 (.A(net53),
    .X(io_out[3]));
 sky130_fd_sc_hd__buf_12 output54 (.A(net54),
    .X(io_out[5]));
 sky130_fd_sc_hd__buf_12 output55 (.A(net55),
    .X(io_out[6]));
 sky130_fd_sc_hd__buf_12 output56 (.A(net56),
    .X(io_out[7]));
 sky130_fd_sc_hd__buf_12 output57 (.A(net57),
    .X(io_out[8]));
 sky130_fd_sc_hd__buf_12 output58 (.A(net58),
    .X(io_out[9]));
 sky130_fd_sc_hd__buf_2 wire92 (.A(_1500_),
    .X(net92));
 assign io_oeb[0] = net186;
 assign io_oeb[10] = net195;
 assign io_oeb[11] = net196;
 assign io_oeb[12] = net197;
 assign io_oeb[13] = net198;
 assign io_oeb[14] = net199;
 assign io_oeb[15] = net200;
 assign io_oeb[16] = net201;
 assign io_oeb[17] = net202;
 assign io_oeb[18] = net203;
 assign io_oeb[19] = net204;
 assign io_oeb[1] = net187;
 assign io_oeb[20] = net205;
 assign io_oeb[21] = net206;
 assign io_oeb[2] = net188;
 assign io_oeb[30] = net215;
 assign io_oeb[31] = net216;
 assign io_oeb[32] = net207;
 assign io_oeb[33] = net208;
 assign io_oeb[34] = net209;
 assign io_oeb[35] = net217;
 assign io_oeb[3] = net189;
 assign io_oeb[4] = net214;
 assign io_oeb[5] = net190;
 assign io_oeb[6] = net191;
 assign io_oeb[7] = net192;
 assign io_oeb[8] = net193;
 assign io_oeb[9] = net194;
 assign io_out[30] = net211;
 assign io_out[31] = net212;
 assign io_out[35] = net213;
 assign io_out[4] = net210;
endmodule

